 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "11000001",3 => "11100100",4 => "01110101",5 => "01010011",6 => "00110011",7 => "11110110",8 => "01010001",9 => "01000111",10 => "01100011",11 => "00110000",12 => "11100111",13 => "10010011",14 => "10011111",15 => "11001101",16 => "10001101",17 => "00001000",18 => "10011110",19 => "11111011",20 => "00111011",21 => "10101000",22 => "00000111",23 => "11011010",24 => "11111011",25 => "01000110",26 => "10010110",27 => "10001000",28 => "01110011",29 => "10000110",30 => "00000000",31 => "00000100",32 => "00111010",33 => "01101010",34 => "11101100",35 => "01110001",36 => "00000101",37 => "01111110",38 => "10010111",39 => "11111110",40 => "00011001",41 => "11011011",42 => "00101010",43 => "00111001",44 => "10110111",45 => "01011001",46 => "11100111",47 => "00010101",48 => "01001110",49 => "11010010",50 => "10101100",51 => "00010010",52 => "11001001",53 => "01001100",54 => "11011010",55 => "11110010",56 => "00111001",57 => "01010000",58 => "10010000",59 => "01111110",60 => "00111100",61 => "00001010",62 => "11011100",63 => "01010001",64 => "01011101",65 => "00101011",66 => "10010101",67 => "01000011",68 => "00010101",69 => "11001001",70 => "00000110",71 => "01000000",72 => "10000101",73 => "10001100",74 => "11100001",75 => "01110101",76 => "00101111",77 => "00110110",78 => "10001011",79 => "11010000",80 => "10010011",81 => "01100011",82 => "10000111",83 => "00101100",84 => "00110011",85 => "11010110",86 => "11101110",87 => "10010111",88 => "01011001",89 => "11110011",90 => "01110101",91 => "11101101",92 => "01111011",93 => "01001000",94 => "11110111",95 => "10110011",96 => "01100101",97 => "00011101",98 => "11011010",99 => "10001100",100 => "01110100",101 => "01100110",102 => "11111101",103 => "00010000",104 => "00110110",105 => "01100111",106 => "00110110",107 => "00110001",108 => "00011100",109 => "10010001",110 => "01011001",111 => "01100110",112 => "00001011",113 => "11011100",114 => "01110000",115 => "00111100",116 => "10110100",117 => "00101011",118 => "10000011",119 => "01010010",120 => "11000011",121 => "10110000",122 => "10111001",123 => "01100001",124 => "01101001",125 => "01100011",126 => "01111110",127 => "10100111",128 => "11110101",129 => "11100111",130 => "11001000",131 => "11110110",132 => "10110111",133 => "01110000",134 => "10001011",135 => "00001010",136 => "10001110",137 => "00001100",138 => "11000011",139 => "00011100",140 => "01010100",141 => "11011000",142 => "00100111",143 => "00100110",144 => "10100100",145 => "10001011",146 => "01101110",147 => "00111110",148 => "00111111",149 => "11101100",150 => "10010000",151 => "10000100",152 => "10111010",153 => "10001000",154 => "01101010",155 => "01110000",156 => "11111101",157 => "11110100",158 => "10111101",159 => "11111100",160 => "01110101",161 => "00100011",162 => "00111001",163 => "00110011",164 => "01000010",165 => "00111001",166 => "10101110",167 => "10101100",168 => "00100010",169 => "11000001",170 => "00001110",171 => "01110011",172 => "00011100",173 => "10000101",174 => "11111011",175 => "10100100",176 => "01100100",177 => "11000010",178 => "11101010",179 => "00001100",180 => "01101011",181 => "11111110",182 => "10101110",183 => "01000000",184 => "00011101",185 => "00001010",186 => "11011000",187 => "01101110",188 => "10001110",189 => "11001100",190 => "10111100",191 => "01101110",192 => "11110001",193 => "01110001",194 => "01101100",195 => "11111110",196 => "01110000",197 => "10101000",198 => "10001100",199 => "01111111",200 => "01001000",201 => "01111101",202 => "11001111",203 => "00000100",204 => "01100101",205 => "01110011",206 => "11110101",207 => "11101101",208 => "10001111",209 => "11101110",210 => "11110011",211 => "10011110",212 => "11100011",213 => "11100111",214 => "11111100",215 => "01110000",216 => "00111010",217 => "11100101",218 => "11001011",219 => "01000110",220 => "11001100",221 => "00001010",222 => "10111011",223 => "01010000",224 => "10111100",225 => "00110101",226 => "00111000",227 => "11101011",228 => "10101100",229 => "00111010",230 => "00010001",231 => "01101101",232 => "01110001",233 => "01100101",234 => "10010011",235 => "00011000",236 => "00011011",237 => "00111111",238 => "00110111",239 => "10111011",240 => "01011101",241 => "11011011",242 => "11110001",243 => "00000010",244 => "01100100",245 => "10101101",246 => "11100111",247 => "00000001",248 => "11110000",249 => "10110011",250 => "01011001",251 => "01111011",252 => "11000010",253 => "10100010",254 => "00100000",255 => "00111011",256 => "00111000",257 => "00001111",258 => "01011101",259 => "10101000",260 => "01011110",261 => "01100001",262 => "01001100",263 => "00101110",264 => "11100100",265 => "11101110",266 => "01110100",267 => "10000011",268 => "01111111",269 => "01110010",270 => "01110000",271 => "10000111",272 => "01101001",273 => "01101100",274 => "01000101",275 => "10000111",276 => "11000110",277 => "10111110",278 => "11100110",279 => "00011001",280 => "10100010",281 => "10111010",282 => "11001110",283 => "10111001",284 => "01100001",285 => "01010101",286 => "01010011",287 => "00001101",288 => "00101001",289 => "11011000",290 => "01101111",291 => "10000110",292 => "00010010",293 => "01011100",294 => "11111110",295 => "00100010",296 => "10001010",297 => "00001011",298 => "01100001",299 => "11110001",300 => "11101101",301 => "11001000",302 => "00110000",303 => "11001011",304 => "00011011",305 => "01010101",306 => "00110001",307 => "00000101",308 => "11111101",309 => "01001001",310 => "01110110",311 => "00110010",312 => "11000101",313 => "01010110",314 => "00001110",315 => "11010101",316 => "10111001",317 => "01111010",318 => "11001011",319 => "11100010",320 => "01001000",321 => "10100101",322 => "01011111",323 => "10010011",324 => "11110010",325 => "01000100",326 => "11000001",327 => "01101101",328 => "01101111",329 => "11011110",330 => "11011010",331 => "00010100",332 => "10000010",333 => "01000101",334 => "10100010",335 => "10101011",336 => "01110100",337 => "00001111",338 => "10100000",339 => "10011001",340 => "11111101",341 => "11001110",342 => "11101101",343 => "11111110",344 => "11011101",345 => "10110010",346 => "11111001",347 => "10000000",348 => "00001111",349 => "11101100",350 => "00111110",351 => "10110010",352 => "01110011",353 => "01001100",354 => "10001110",355 => "01111011",356 => "01010110",357 => "11111110",358 => "10100000",359 => "10100001",360 => "11000010",361 => "01010100",362 => "11100100",363 => "01001011",364 => "01100000",365 => "00110010",366 => "11111000",367 => "11111010",368 => "10110010",369 => "01000110",370 => "11011100",371 => "11110010",372 => "01110100",373 => "10100110",374 => "10000001",375 => "11011001",376 => "01101111",377 => "00011101",378 => "10000001",379 => "01001110",380 => "11010110",381 => "10110101",382 => "01101000",383 => "11011110",384 => "00111100",385 => "01101100",386 => "01011100",387 => "01110011",388 => "10010100",389 => "00000010",390 => "10110110",391 => "10100011",392 => "11000000",393 => "01011111",394 => "10101001",395 => "10010111",396 => "11010011",397 => "10011100",398 => "10010011",399 => "01001010",400 => "01010101",401 => "00101000",402 => "10111010",403 => "11110011",404 => "10011010",405 => "10000001",406 => "01011111",407 => "01011110",408 => "11100010",409 => "10111000",410 => "00001001",411 => "01010101",412 => "00101000",413 => "00101101",414 => "01101001",415 => "11001101",416 => "00011101",417 => "00000100",418 => "00000101",419 => "11111111",420 => "11000101",421 => "11111001",422 => "00100001",423 => "00100000",424 => "00001000",425 => "00100100",426 => "00110011",427 => "11001001",428 => "11111010",429 => "01001100",430 => "00100001",431 => "10011110",432 => "01011010",433 => "00000111",434 => "01001000",435 => "01001101",436 => "01100111",437 => "10110100",438 => "01011011",439 => "01111111",440 => "00101101",441 => "01110001",442 => "01010001",443 => "01111010",444 => "00010111",445 => "00101111",446 => "00100000",447 => "11100101",448 => "00100100",449 => "01111011",450 => "01100101",451 => "01101101",452 => "10101111",453 => "10001001",454 => "01010001",455 => "11101001",456 => "01010010",457 => "00100101",458 => "11010100",459 => "11011111",460 => "00011100",461 => "10101001",462 => "00011011",463 => "11100101",464 => "00100011",465 => "10001000",466 => "00101001",467 => "00010101",468 => "10100100",469 => "10001110",470 => "00000100",471 => "10100000",472 => "00110110",473 => "00111000",474 => "00110100",475 => "01100011",476 => "00111001",477 => "00001010",478 => "11001100",479 => "11000000",480 => "10101110",481 => "00001111",482 => "00001001",483 => "00101110",484 => "00100101",485 => "01011111",486 => "01100010",487 => "00111010",488 => "01111101",489 => "10010000",490 => "00001111",491 => "01001011",492 => "01001100",493 => "10101010",494 => "11101011",495 => "11010011",496 => "10111110",497 => "00010011",498 => "11110000",499 => "10101000",500 => "11011110",501 => "11110010",502 => "01010101",503 => "11001101",504 => "00111010",505 => "01001010",506 => "01010100",507 => "00111110",508 => "00110111",509 => "10011001",510 => "11011000",511 => "11111100",512 => "11010001",513 => "00010011",514 => "01001001",515 => "01100101",516 => "01100111",517 => "01100000",518 => "11101100",519 => "01000010",520 => "11101011",521 => "11011111",522 => "10011001",523 => "01101011",524 => "11010100",525 => "00111111",526 => "10001001",527 => "01110000",528 => "01111011",529 => "10110110",530 => "00110011",531 => "10010011",532 => "01000110",533 => "01111101",534 => "00001101",535 => "01101111",536 => "00001010",537 => "01000110",538 => "00101000",539 => "01110100",540 => "00100111",541 => "00100111",542 => "01100110",543 => "00100011",544 => "10000011",545 => "10100011",546 => "00101101",547 => "00100000",548 => "01000011",549 => "11101111",550 => "01000000",551 => "01101110",552 => "00011011",553 => "01011000",554 => "01111100",555 => "11011000",556 => "11000101",557 => "00000011",558 => "00100011",559 => "11110000",560 => "11011111",561 => "10101111",562 => "11011100",563 => "00110110",564 => "00101100",565 => "00000100",566 => "11001110",567 => "10010101",568 => "11011101",569 => "11101100",570 => "11111001",571 => "01110111",572 => "00001111",573 => "00011010",574 => "11001111",575 => "11000101",576 => "00110110",577 => "11100000",578 => "01000001",579 => "01111110",580 => "10101101",581 => "10001000",582 => "00101101",583 => "10101000",584 => "11110111",585 => "10110100",586 => "11101010",587 => "00011010",588 => "10000100",589 => "10100000",590 => "00100111",591 => "01100111",592 => "11001010",593 => "01001110",594 => "01100100",595 => "00000110",596 => "10101010",597 => "10110010",598 => "01100011",599 => "01011001",600 => "11101111",601 => "10110100",602 => "00100011",603 => "00000101",604 => "11010100",605 => "11011000",606 => "00011010",607 => "11100001",608 => "00011110",609 => "10101110",610 => "10010100",611 => "11111001",612 => "11000100",613 => "10111010",614 => "11101011",615 => "11101110",616 => "10110110",617 => "11001100",618 => "11101011",619 => "11001101",620 => "00100111",621 => "10000000",622 => "10100100",623 => "10110100",624 => "10110111",625 => "10011100",626 => "10001111",627 => "11101111",628 => "00001000",629 => "00100000",630 => "00111111",631 => "11110000",632 => "11011010",633 => "11011100",634 => "01011100",635 => "00101011",636 => "00100011",637 => "01000110",638 => "11001100",639 => "10000000",640 => "00010000",641 => "10101101",642 => "00000110",643 => "10000001",644 => "01011011",645 => "11010110",646 => "11001101",647 => "10010011",648 => "11010111",649 => "01111011",650 => "11001101",651 => "10101001",652 => "11010111",653 => "01110100",654 => "01110111",655 => "00000100",656 => "11111100",657 => "00001101",658 => "10001111",659 => "10011011",660 => "11000110",661 => "01110100",662 => "00110010",663 => "11000100",664 => "11111101",665 => "00100000",666 => "11000110",667 => "11111001",668 => "00110101",669 => "01011101",670 => "10111101",671 => "10100111",672 => "00010100",673 => "00110111",674 => "11100001",675 => "00001010",676 => "11010101",677 => "11110010",678 => "00110001",679 => "11110001",680 => "11001111",681 => "11100111",682 => "01010101",683 => "00111010",684 => "10100101",685 => "11111111",686 => "00000100",687 => "11111011",688 => "10010100",689 => "10100011",690 => "11010110",691 => "00100101",692 => "10000011",693 => "11010110",694 => "00010000",695 => "10111011",696 => "11011001",697 => "00011001",698 => "01001000",699 => "10111011",700 => "01001111",701 => "01101010",702 => "10011001",703 => "00101110",704 => "00111011",705 => "11011000",706 => "10111000",707 => "10111010",708 => "10110110",709 => "10111100",710 => "10110110",711 => "11001000",712 => "00110111",713 => "10110001",714 => "01100111",715 => "10011110",716 => "11101011",717 => "11010100",718 => "00010000",719 => "11101010",720 => "01111011",721 => "11000000",722 => "11010001",723 => "00011101",724 => "00100101",725 => "01010100",726 => "01011010",727 => "10100110",728 => "10001001",729 => "10111011",730 => "11111000",731 => "10011010",732 => "00111110",733 => "00110111",734 => "11100101",735 => "00110110",736 => "01001101",737 => "11000000",738 => "01000101",739 => "11001110",740 => "10101001",741 => "10110111",742 => "11000010",743 => "11101101",744 => "00001000",745 => "10101111",746 => "00111111",747 => "00001110",748 => "01101001",749 => "01010110",750 => "00110110",751 => "11100011",752 => "00111100",753 => "01101010",754 => "00001011",755 => "01011111",756 => "10001110",757 => "00010100",758 => "11100111",759 => "10010011",760 => "00000000",761 => "00010011",762 => "01111110",763 => "11001000",764 => "11111110",765 => "00001110",766 => "10101101",767 => "01001011",768 => "11010000",769 => "00001101",770 => "01101100",771 => "10001001",772 => "01000000",773 => "00000101",774 => "01110000",775 => "11100101",776 => "01111000",777 => "10111011",778 => "01101110",779 => "11101110",780 => "10100000",781 => "11001010",782 => "10001110",783 => "11001000",784 => "11001000",785 => "01011000",786 => "01010100",787 => "00101100",788 => "10100110",789 => "10000101",790 => "11110110",791 => "00111100",792 => "01100001",793 => "00010000",794 => "11110001",795 => "11010100",796 => "00000011",797 => "01111011",798 => "10110100",799 => "00101011",800 => "10110011",801 => "00001100",802 => "01100011",803 => "10001011",804 => "10111111",805 => "01010001",806 => "00111010",807 => "11011001",808 => "00101100",809 => "11000010",810 => "01000111",811 => "10000110",812 => "00001001",813 => "11011110",814 => "10010101",815 => "00110110",816 => "00010110",817 => "00010011",818 => "10000011",819 => "00001011",820 => "10000001",821 => "10110000",822 => "01110010",823 => "00001111",824 => "11010001",825 => "01011010",826 => "11011111",827 => "01101110",828 => "10110100",829 => "00001010",830 => "00101110",831 => "10000111",832 => "10001001",833 => "11011110",834 => "00010011",835 => "00110010",836 => "00011011",837 => "10000100",838 => "00110001",839 => "11011110",840 => "00101111",841 => "01011000",842 => "10111100",843 => "11100101",844 => "10001110",845 => "00110110",846 => "10110101",847 => "00001110",848 => "00111000",849 => "01111011",850 => "11100101",851 => "01101111",852 => "10000000",853 => "01111110",854 => "00010011",855 => "00010000",856 => "11100110",857 => "00001011",858 => "11000100",859 => "01000110",860 => "00011000",861 => "10011010",862 => "11001111",863 => "10100011",864 => "01011000",865 => "01111001",866 => "11111010",867 => "10000110",868 => "01110101",869 => "01100101",870 => "11101111",871 => "01000111",872 => "10001101",873 => "11100001",874 => "01000010",875 => "11101000",876 => "10110011",877 => "11101100",878 => "01101100",879 => "01000011",880 => "11100010",881 => "00110110",882 => "01010000",883 => "00110101",884 => "00011010",885 => "11011000",886 => "10010111",887 => "10100001",888 => "10001000",889 => "11001110",890 => "01111110",891 => "11000101",892 => "11010110",893 => "11001010",894 => "01001011",895 => "00010100",896 => "01101000",897 => "10001010",898 => "11100111",899 => "00010110",900 => "00011110",901 => "10101111",902 => "00100111",903 => "00100010",904 => "11110010",905 => "01100100",906 => "00011001",907 => "11011110",908 => "10010010",909 => "01111000",910 => "10000100",911 => "01010100",912 => "00111010",913 => "01000001",914 => "00010000",915 => "00010101",916 => "00001100",917 => "10101111",918 => "00011001",919 => "01000101",920 => "00011101",921 => "01011010",922 => "11111100",923 => "01110000",924 => "01101100",925 => "00000101",926 => "00111001",927 => "11111110",928 => "01101010",929 => "00100100",930 => "01111100",931 => "00100100",932 => "10101101",933 => "00110100",934 => "01001101",935 => "10101011",936 => "10011001",937 => "01100011",938 => "00111011",939 => "01000110",940 => "11011011",941 => "01010100",942 => "11100011",943 => "11101100",944 => "11100010",945 => "11011000",946 => "11110111",947 => "11010100",948 => "10100010",949 => "00101110",950 => "10111010",951 => "10111010",952 => "11111001",953 => "11110100",954 => "01101001",955 => "11000111",956 => "11101001",957 => "00000000",958 => "10101011",959 => "01111101",960 => "11010011",961 => "00110111",962 => "10110101",963 => "00001100",964 => "00001110",965 => "10001110",966 => "00101111",967 => "11101100",968 => "00010111",969 => "10000011",970 => "01101110",971 => "00110101",972 => "10100000",973 => "00010000",974 => "01111011",975 => "10100011",976 => "10011010",977 => "01100000",978 => "01111110",979 => "01011100",980 => "01111001",981 => "01101001",982 => "11000100",983 => "10000101",984 => "11100100",985 => "10001111",986 => "11001101",987 => "11001111",988 => "01011000",989 => "00001000",990 => "11110100",991 => "01101101",992 => "11010111",993 => "00110111",994 => "11001110",995 => "00110110",996 => "11010000",997 => "11111100",998 => "00101011",999 => "10000000",1000 => "10010011",1001 => "01001101",1002 => "11011111",1003 => "11010011",1004 => "01110100",1005 => "00111000",1006 => "11110101",1007 => "00111011",1008 => "01100100",1009 => "11100110",1010 => "00101011",1011 => "11111101",1012 => "10011101",1013 => "11111111",1014 => "00110101",1015 => "11110001",1016 => "01100100",1017 => "01011000",1018 => "00011110",1019 => "01000010",1020 => "00000010",1021 => "10100101",1022 => "11110000",1023 => "00010100",1024 => "10110001",1025 => "11010111",1026 => "01010110",1027 => "00011100",1028 => "10111011",1029 => "10010000",1030 => "11011001",1031 => "11110100",1032 => "01010000",1033 => "10000010",1034 => "00101111",1035 => "10110000",1036 => "01100010",1037 => "10010110",1038 => "01011000",1039 => "10011011",1040 => "01001011",1041 => "00100001",1042 => "00100010",1043 => "00011111",1044 => "11100111",1045 => "10111110",1046 => "11111110",1047 => "10111000",1048 => "01101011",1049 => "10100000",1050 => "00111000",1051 => "01111110",1052 => "11110001",1053 => "01110100",1054 => "00101101",1055 => "00011001",1056 => "01000110",1057 => "01110110",1058 => "10111000",1059 => "01010000",1060 => "11101000",1061 => "00111110",1062 => "11110101",1063 => "01101111",1064 => "10101110",1065 => "01110111",1066 => "00011000",1067 => "10101011",1068 => "11000011",1069 => "01100110",1070 => "01011101",1071 => "11110010",1072 => "11101100",1073 => "11101110",1074 => "00100110",1075 => "10000000",1076 => "00111000",1077 => "10101010",1078 => "01111100",1079 => "00110000",1080 => "10101100",1081 => "01111001",1082 => "00100111",1083 => "10101111",1084 => "00000100",1085 => "11010111",1086 => "11001001",1087 => "01001100",1088 => "11111010",1089 => "00010111",1090 => "10110100",1091 => "01000011",1092 => "11110000",1093 => "00000100",1094 => "11001111",1095 => "00110010",1096 => "11100111",1097 => "01100101",1098 => "00100010",1099 => "00010001",1100 => "01001011",1101 => "01000111",1102 => "10001001",1103 => "00111101",1104 => "11001111",1105 => "00101000",1106 => "11101100",1107 => "00101101",1108 => "10001101",1109 => "11000111",1110 => "10001011",1111 => "00101110",1112 => "00100000",1113 => "10110000",1114 => "11011010",1115 => "10001101",1116 => "01111000",1117 => "10011011",1118 => "01010011",1119 => "00101101",1120 => "11010000",1121 => "00111111",1122 => "10001000",1123 => "00100001",1124 => "00111001",1125 => "00010100",1126 => "10010010",1127 => "11001100",1128 => "00001101",1129 => "00101111",1130 => "10110100",1131 => "11111000",1132 => "01110001",1133 => "01011101",1134 => "00000011",1135 => "11100101",1136 => "10011101",1137 => "00011100",1138 => "00001010",1139 => "00101011",1140 => "11001101",1141 => "10011010",1142 => "11101011",1143 => "10100010",1144 => "10000111",1145 => "10000001",1146 => "10011111",1147 => "00001001",1148 => "00000110",1149 => "11101100",1150 => "00100111",1151 => "00101001",1152 => "11011111",1153 => "00001100",1154 => "10001110",1155 => "01110100",1156 => "01001010",1157 => "01001000",1158 => "11100001",1159 => "10101110",1160 => "10000011",1161 => "00101111",1162 => "01010101",1163 => "10101110",1164 => "11111101",1165 => "01000000",1166 => "01101001",1167 => "01000011",1168 => "10010000",1169 => "11101010",1170 => "10111011",1171 => "10111000",1172 => "10100011",1173 => "01100000",1174 => "10000100",1175 => "00011011",1176 => "01011100",1177 => "10100010",1178 => "01010011",1179 => "01011001",1180 => "01100111",1181 => "10111111",1182 => "11111001",1183 => "10010000",1184 => "11100111",1185 => "10000011",1186 => "00100111",1187 => "11010100",1188 => "01111010",1189 => "10011110",1190 => "01110001",1191 => "00010000",1192 => "11010110",1193 => "00101110",1194 => "11111100",1195 => "11011001",1196 => "11101111",1197 => "01001001",1198 => "00111011",1199 => "10100111",1200 => "00100100",1201 => "00011101",1202 => "01111100",1203 => "00001100",1204 => "00111100",1205 => "11000011",1206 => "00011010",1207 => "00011101",1208 => "00011011",1209 => "10011100",1210 => "01100110",1211 => "10101110",1212 => "11000011",1213 => "10011101",1214 => "00000110",1215 => "10110001",1216 => "01110010",1217 => "01000011",1218 => "01111001",1219 => "10010000",1220 => "10011100",1221 => "10101000",1222 => "00101110",1223 => "10101110",1224 => "00100010",1225 => "00011100",1226 => "01100011",1227 => "11000101",1228 => "00001101",1229 => "11111110",1230 => "10111011",1231 => "11000111",1232 => "01011011",1233 => "11001110",1234 => "00100111",1235 => "11111100",1236 => "11001111",1237 => "00001111",1238 => "10101100",1239 => "11110001",1240 => "11011110",1241 => "01111111",1242 => "01111101",1243 => "01101101",1244 => "01111101",1245 => "10111100",1246 => "00111010",1247 => "11101110",1248 => "10110010",1249 => "10110111",1250 => "00101100",1251 => "01111101",1252 => "10001001",1253 => "10111010",1254 => "00110101",1255 => "10010011",1256 => "01110101",1257 => "10111110",1258 => "10000011",1259 => "10100011",1260 => "11100011",1261 => "10001111",1262 => "11010001",1263 => "11011010",1264 => "00100010",1265 => "11111101",1266 => "10101010",1267 => "11101001",1268 => "00101110",1269 => "01101100",1270 => "01101110",1271 => "11100111",1272 => "00001111",1273 => "11011001",1274 => "11010100",1275 => "11110111",1276 => "01100100",1277 => "00001010",1278 => "00010100",1279 => "01111001",1280 => "10010110",1281 => "01001000",1282 => "11110101",1283 => "01100010",1284 => "01010101",1285 => "00011111",1286 => "01000010",1287 => "01100001",1288 => "01011011",1289 => "01001111",1290 => "01010100",1291 => "00111110",1292 => "10000010",1293 => "01011010",1294 => "10010010",1295 => "01101000",1296 => "10000101",1297 => "11011001",1298 => "11001111",1299 => "00011010",1300 => "00000111",1301 => "01001011",1302 => "00011001",1303 => "10100010",1304 => "11010100",1305 => "11100100",1306 => "00111111",1307 => "11011100",1308 => "11100000",1309 => "01011011",1310 => "10010000",1311 => "01011110",1312 => "00100101",1313 => "01110101",1314 => "00111000",1315 => "00111110",1316 => "01001010",1317 => "00111111",1318 => "00011010",1319 => "01011000",1320 => "01100111",1321 => "11010001",1322 => "10011000",1323 => "00101000",1324 => "10001111",1325 => "01100000",1326 => "11101100",1327 => "01001000",1328 => "00011010",1329 => "01110100",1330 => "11111100",1331 => "01011010",1332 => "00001101",1333 => "00010001",1334 => "10100001",1335 => "11010111",1336 => "01011000",1337 => "00111110",1338 => "00010111",1339 => "10001011",1340 => "00011101",1341 => "00000111",1342 => "10001100",1343 => "10110011",1344 => "10110100",1345 => "01111101",1346 => "11011010",1347 => "10100111",1348 => "01100000",1349 => "01100000",1350 => "11000110",1351 => "01100001",1352 => "11111001",1353 => "10000101",1354 => "01110000",1355 => "00110110",1356 => "00001010",1357 => "01101100",1358 => "11010100",1359 => "10101100",1360 => "01011111",1361 => "00101011",1362 => "00010111",1363 => "01100100",1364 => "01111010",1365 => "10001100",1366 => "10010001",1367 => "11111100",1368 => "10111000",1369 => "01100111",1370 => "00101011",1371 => "10011011",1372 => "11011110",1373 => "11101011",1374 => "00010010",1375 => "11111000",1376 => "11011110",1377 => "11010010",1378 => "10011001",1379 => "01110001",1380 => "10010111",1381 => "01110001",1382 => "01101110",1383 => "01001001",1384 => "00100001",1385 => "10101101",1386 => "00010111",1387 => "00000011",1388 => "01100110",1389 => "01110101",1390 => "00110110",1391 => "01110110",1392 => "11000111",1393 => "00000001",1394 => "10100101",1395 => "00010010",1396 => "11011100",1397 => "11010111",1398 => "01111110",1399 => "01000000",1400 => "11011001",1401 => "00001101",1402 => "11101010",1403 => "01110001",1404 => "00110110",1405 => "00011101",1406 => "01101000",1407 => "01000001",1408 => "11100011",1409 => "11000010",1410 => "10101111",1411 => "10111010",1412 => "00000011",1413 => "00001111",1414 => "11011100",1415 => "11101000",1416 => "10101001",1417 => "11110100",1418 => "00010110",1419 => "11101000",1420 => "00011100",1421 => "01011010",1422 => "00110000",1423 => "00110111",1424 => "10000000",1425 => "01001110",1426 => "10111101",1427 => "00111111",1428 => "11000011",1429 => "01010111",1430 => "10000001",1431 => "11110111",1432 => "01010101",1433 => "01100101",1434 => "00001001",1435 => "11101011",1436 => "01001001",1437 => "00111101",1438 => "11001101",1439 => "10000001",1440 => "00001100",1441 => "10111101",1442 => "01101000",1443 => "10100011",1444 => "01011001",1445 => "11101000",1446 => "00010100",1447 => "01111011",1448 => "11010011",1449 => "11000100",1450 => "10101110",1451 => "11001100",1452 => "10110011",1453 => "10001100",1454 => "00011101",1455 => "11000110",1456 => "10111000",1457 => "11010100",1458 => "10010100",1459 => "00001111",1460 => "00000111",1461 => "10011111",1462 => "00001101",1463 => "00000110",1464 => "11110100",1465 => "01001111",1466 => "11011110",1467 => "01000000",1468 => "11100001",1469 => "01000000",1470 => "01100100",1471 => "10110110",1472 => "10001100",1473 => "01110011",1474 => "00100011",1475 => "10010010",1476 => "11111001",1477 => "10101011",1478 => "10101011",1479 => "00100001",1480 => "10000111",1481 => "01110100",1482 => "10100001",1483 => "11111111",1484 => "10111001",1485 => "10101001",1486 => "00011001",1487 => "01110100",1488 => "10111000",1489 => "11101101",1490 => "00011011",1491 => "10000101",1492 => "11000011",1493 => "11001101",1494 => "11011111",1495 => "10101110",1496 => "01011100",1497 => "01101000",1498 => "11111010",1499 => "10100100",1500 => "00001000",1501 => "00111011",1502 => "10111011",1503 => "11101100",1504 => "11010101",1505 => "11010010",1506 => "01100001",1507 => "10110100",1508 => "01010010",1509 => "01110100",1510 => "01000001",1511 => "10010000",1512 => "00111110",1513 => "10111101",1514 => "10001100",1515 => "01010011",1516 => "10101000",1517 => "01010111",1518 => "11101001",1519 => "10111000",1520 => "11100100",1521 => "10100100",1522 => "01010101",1523 => "11101101",1524 => "10001001",1525 => "10100100",1526 => "00101000",1527 => "11110001",1528 => "10101101",1529 => "01001010",1530 => "11001011",1531 => "00011011",1532 => "10001100",1533 => "11010111",1534 => "01101111",1535 => "00010100",1536 => "11110111",1537 => "10011100",1538 => "01110101",1539 => "00010111",1540 => "10110110",1541 => "01111011",1542 => "01000011",1543 => "11010000",1544 => "11111010",1545 => "00111100",1546 => "01010110",1547 => "01111011",1548 => "11101001",1549 => "10010011",1550 => "11000010",1551 => "10001100",1552 => "01101101",1553 => "11100111",1554 => "10000110",1555 => "11001110",1556 => "01111000",1557 => "00010110",1558 => "11011001",1559 => "10010100",1560 => "00010000",1561 => "10010001",1562 => "10010100",1563 => "01011100",1564 => "10111110",1565 => "01011000",1566 => "00100000",1567 => "11001000",1568 => "11111100",1569 => "11011000",1570 => "00100100",1571 => "10001111",1572 => "10100100",1573 => "00000000",1574 => "11011101",1575 => "01001110",1576 => "11010011",1577 => "01011011",1578 => "00011000",1579 => "01101011",1580 => "00110111",1581 => "00111100",1582 => "10110100",1583 => "11000011",1584 => "11010000",1585 => "01011100",1586 => "10111100",1587 => "10000101",1588 => "11100100",1589 => "10010001",1590 => "11111000",1591 => "10101011",1592 => "00101101",1593 => "10011001",1594 => "10101011",1595 => "00010010",1596 => "01100100",1597 => "01100101",1598 => "10000101",1599 => "00010101",1600 => "11011111",1601 => "00101100",1602 => "00111101",1603 => "00001100",1604 => "10010101",1605 => "00111010",1606 => "11111011",1607 => "01100000",1608 => "00111100",1609 => "11101010",1610 => "01110111",1611 => "00010000",1612 => "11000000",1613 => "00011011",1614 => "10110011",1615 => "10100111",1616 => "00100000",1617 => "00000010",1618 => "11111110",1619 => "00000001",1620 => "01110011",1621 => "10101111",1622 => "10000000",1623 => "00010010",1624 => "01100101",1625 => "10010111",1626 => "01010000",1627 => "10001110",1628 => "00011011",1629 => "01000011",1630 => "00010011",1631 => "00101010",1632 => "10001000",1633 => "00001101",1634 => "10001101",1635 => "10111001",1636 => "10101000",1637 => "10101001",1638 => "11001000",1639 => "11011000",1640 => "01010010",1641 => "11111010",1642 => "00000101",1643 => "01011001",1644 => "00011000",1645 => "11010111",1646 => "11001101",1647 => "10100100",1648 => "01111100",1649 => "00000101",1650 => "10010010",1651 => "10000000",1652 => "00011011",1653 => "11101111",1654 => "10001000",1655 => "11110000",1656 => "01100100",1657 => "11010011",1658 => "01000001",1659 => "01010101",1660 => "00110001",1661 => "10011010",1662 => "01010101",1663 => "11110010",1664 => "00011101",1665 => "11101011",1666 => "00000100",1667 => "00110011",1668 => "01010001",1669 => "00111010",1670 => "00100111",1671 => "11011001",1672 => "00111001",1673 => "10101100",1674 => "01110101",1675 => "10001110",1676 => "00100100",1677 => "11101011",1678 => "11111000",1679 => "00111000",1680 => "11101011",1681 => "01001000",1682 => "11010010",1683 => "00110000",1684 => "11000011",1685 => "00111010",1686 => "10010110",1687 => "01001101",1688 => "01111101",1689 => "01101111",1690 => "10001101",1691 => "10000100",1692 => "00010010",1693 => "10100000",1694 => "00111101",1695 => "00010011",1696 => "11010011",1697 => "01101001",1698 => "11000111",1699 => "11111101",1700 => "01110010",1701 => "11000111",1702 => "11111110",1703 => "10001010",1704 => "10101001",1705 => "00011001",1706 => "00001000",1707 => "11111001",1708 => "01101100",1709 => "10001000",1710 => "00111001",1711 => "01010011",1712 => "11100101",1713 => "00011011",1714 => "10000110",1715 => "11010101",1716 => "01101111",1717 => "10110001",1718 => "10101011",1719 => "00100111",1720 => "01110001",1721 => "11000010",1722 => "11111110",1723 => "01001001",1724 => "01101011",1725 => "11101100",1726 => "00110000",1727 => "11011000",1728 => "00011000",1729 => "00110010",1730 => "00111101",1731 => "00010100",1732 => "10110101",1733 => "00000101",1734 => "10001101",1735 => "00110101",1736 => "00101111",1737 => "10101011",1738 => "01001110",1739 => "01000001",1740 => "11010011",1741 => "00100010",1742 => "10110010",1743 => "01011111",1744 => "10011010",1745 => "00110010",1746 => "10000001",1747 => "00001101",1748 => "10001011",1749 => "10010001",1750 => "00001000",1751 => "01100110",1752 => "01000011",1753 => "00101101",1754 => "00100111",1755 => "10001010",1756 => "11111111",1757 => "11010001",1758 => "10011010",1759 => "11111110",1760 => "10100000",1761 => "10010101",1762 => "00101011",1763 => "00101100",1764 => "11100100",1765 => "10101101",1766 => "11100000",1767 => "00000000",1768 => "11000100",1769 => "00100011",1770 => "11110010",1771 => "11101000",1772 => "00010010",1773 => "11001001",1774 => "11011101",1775 => "11101110",1776 => "01110101",1777 => "10100011",1778 => "10010101",1779 => "10001110",1780 => "11000111",1781 => "10111001",1782 => "10110100",1783 => "11111101",1784 => "11111110",1785 => "01110100",1786 => "11110101",1787 => "00100101",1788 => "10010101",1789 => "01001001",1790 => "11110110",1791 => "10000000",1792 => "10110110",1793 => "01101011",1794 => "11101010",1795 => "01001111",1796 => "01001011",1797 => "10110100",1798 => "01011101",1799 => "10100100",1800 => "00011001",1801 => "10000001",1802 => "11001111",1803 => "01000000",1804 => "11101111",1805 => "11000011",1806 => "10111000",1807 => "00010101",1808 => "00000001",1809 => "00101011",1810 => "10010011",1811 => "10011100",1812 => "10011011",1813 => "11010111",1814 => "10001010",1815 => "00001000",1816 => "11001011",1817 => "10010010",1818 => "00111110",1819 => "01001110",1820 => "00101110",1821 => "10110101",1822 => "00111000",1823 => "11101100",1824 => "00111110",1825 => "11011110",1826 => "01111110",1827 => "01001000",1828 => "01011101",1829 => "11101110",1830 => "00000100",1831 => "10000001",1832 => "00100111",1833 => "11010100",1834 => "10000111",1835 => "11011011",1836 => "10000010",1837 => "01010101",1838 => "01111101",1839 => "10011001",1840 => "00000011",1841 => "10001110",1842 => "11111000",1843 => "10101111",1844 => "10000011",1845 => "11001011",1846 => "01111000",1847 => "01100100",1848 => "10110010",1849 => "00110010",1850 => "01110111",1851 => "01111100",1852 => "00000010",1853 => "01111011",1854 => "10001100",1855 => "11010101",1856 => "00100010",1857 => "11101110",1858 => "01101011",1859 => "00011001",1860 => "11011000",1861 => "11110110",1862 => "01100100",1863 => "10001110",1864 => "10011011",1865 => "10101010",1866 => "11010111",1867 => "00010110",1868 => "10000111",1869 => "10110101",1870 => "01100000",1871 => "01011110",1872 => "10100110",1873 => "01000111",1874 => "00011011",1875 => "10000101",1876 => "00001111",1877 => "10101110",1878 => "10110111",1879 => "11101011",1880 => "01101000",1881 => "10100110",1882 => "01001011",1883 => "10011101",1884 => "10001110",1885 => "01111111",1886 => "10011101",1887 => "00100001",1888 => "11010001",1889 => "00110111",1890 => "11111000",1891 => "01110100",1892 => "11000100",1893 => "10000100",1894 => "01111111",1895 => "11100110",1896 => "00110101",1897 => "10011110",1898 => "00000110",1899 => "00110010",1900 => "10110001",1901 => "01111100",1902 => "00011011",1903 => "00000110",1904 => "10101101",1905 => "00100000",1906 => "11000011",1907 => "01111111",1908 => "11100010",1909 => "10111010",1910 => "00011010",1911 => "10000110",1912 => "11100010",1913 => "01000101",1914 => "10011110",1915 => "01010011",1916 => "01110111",1917 => "01001111",1918 => "01101011",1919 => "00000111",1920 => "10001011",1921 => "00001110",1922 => "00000001",1923 => "11101111",1924 => "11101000",1925 => "10010010",1926 => "00101011",1927 => "01010010",1928 => "11000000",1929 => "01101100",1930 => "10001001",1931 => "10111100",1932 => "00101010",1933 => "00011000",1934 => "01000101",1935 => "10100010",1936 => "11101000",1937 => "11011110",1938 => "01010111",1939 => "10011000",1940 => "10000011",1941 => "00101010",1942 => "00101010",1943 => "00000100",1944 => "10110101",1945 => "10001100",1946 => "11011111",1947 => "00101001",1948 => "10011110",1949 => "01001010",1950 => "00101110",1951 => "10110110",1952 => "00101101",1953 => "01110110",1954 => "01111001",1955 => "01111001",1956 => "00011111",1957 => "01010100",1958 => "10001100",1959 => "11100010",1960 => "11011010",1961 => "00001001",1962 => "11011100",1963 => "11000111",1964 => "11010010",1965 => "10110001",1966 => "10000010",1967 => "01110101",1968 => "10001100",1969 => "01010000",1970 => "11110111",1971 => "01101011",1972 => "00000100",1973 => "01001000",1974 => "10000101",1975 => "01001000",1976 => "11101001",1977 => "00000010",1978 => "11001100",1979 => "01111110",1980 => "00110100",1981 => "01110010",1982 => "01101110",1983 => "00010011",1984 => "00010010",1985 => "10011100",1986 => "10010110",1987 => "10000110",1988 => "11111011",1989 => "11100111",1990 => "10001000",1991 => "00010010",1992 => "11001011",1993 => "10001110",1994 => "11011111",1995 => "11001011",1996 => "01011110",1997 => "10111101",1998 => "11111010",1999 => "00011011",2000 => "11111010",2001 => "10010111",2002 => "00100000",2003 => "11111110",2004 => "10000001",2005 => "00001101",2006 => "00101000",2007 => "01111100",2008 => "10011101",2009 => "11100000",2010 => "10100100",2011 => "11111101",2012 => "01001101",2013 => "10100111",2014 => "10111010",2015 => "11101010",2016 => "11100001",2017 => "00100011",2018 => "01001100",2019 => "10111000",2020 => "10110011",2021 => "10010000",2022 => "00111001",2023 => "11100111",2024 => "01100001",2025 => "00110100",2026 => "11011110",2027 => "01010011",2028 => "11101111",2029 => "01111001",2030 => "01101001",2031 => "10000001",2032 => "11000010",2033 => "01010101",2034 => "01010110",2035 => "00101010",2036 => "01010111",2037 => "01110001",2038 => "11000001",2039 => "11111111",2040 => "11001110",2041 => "11100010",2042 => "10000111",2043 => "00011111",2044 => "11101001",2045 => "01011110",2046 => "01010111",2047 => "01101001",2048 => "00101111",2049 => "01001001",2050 => "11011111",2051 => "11101110",2052 => "11110000",2053 => "10011000",2054 => "00000001",2055 => "01011100",2056 => "00000011",2057 => "11110101",2058 => "10111011",2059 => "10101001",2060 => "10110011",2061 => "00001010",2062 => "10001010",2063 => "00001001",2064 => "11111010",2065 => "00011100",2066 => "10101111",2067 => "11001110",2068 => "11111001",2069 => "01010101",2070 => "11101110",2071 => "10000101",2072 => "10011010",2073 => "00100000",2074 => "11011000",2075 => "11011000",2076 => "00100010",2077 => "11011000",2078 => "00010101",2079 => "01010111",2080 => "10001111",2081 => "00110010",2082 => "00110011",2083 => "00011111",2084 => "01111000",2085 => "01010111",2086 => "01111011",2087 => "00110001",2088 => "00101001",2089 => "10100101",2090 => "01011100",2091 => "00101010",2092 => "01010000",2093 => "11101011",2094 => "11010111",2095 => "10011001",2096 => "10101101",2097 => "00100010",2098 => "00110000",2099 => "01111111",2100 => "00000101",2101 => "00110111",2102 => "01100101",2103 => "11000001",2104 => "01101111",2105 => "11000011",2106 => "01111100",2107 => "10110010",2108 => "01000101",2109 => "10001000",2110 => "10011101",2111 => "01001011",2112 => "10101000",2113 => "01011011",2114 => "01010100",2115 => "01100000",2116 => "00110000",2117 => "11001001",2118 => "11100111",2119 => "10110000",2120 => "11010001",2121 => "11100111",2122 => "00000011",2123 => "01111100",2124 => "00000010",2125 => "01000011",2126 => "10011110",2127 => "00000101",2128 => "00010001",2129 => "01010100",2130 => "00100001",2131 => "00110001",2132 => "00011111",2133 => "00001100",2134 => "11101100",2135 => "10001111",2136 => "11001111",2137 => "10101100",2138 => "00010101",2139 => "11010001",2140 => "10101110",2141 => "00001000",2142 => "11111100",2143 => "01110110",2144 => "00001101",2145 => "10011101",2146 => "01100101",2147 => "10111011",2148 => "10101110",2149 => "11111110",2150 => "10111110",2151 => "10101100",2152 => "01011100",2153 => "00100111",2154 => "10001111",2155 => "01100111",2156 => "00010010",2157 => "00110100",2158 => "00111000",2159 => "01100011",2160 => "00100011",2161 => "11010111",2162 => "01011101",2163 => "00101011",2164 => "00110000",2165 => "00111100",2166 => "11001100",2167 => "11101101",2168 => "11000010",2169 => "00111100",2170 => "10110011",2171 => "00010100",2172 => "10100101",2173 => "01101011",2174 => "00110110",2175 => "00110111",2176 => "01101010",2177 => "11000110",2178 => "01010100",2179 => "10111001",2180 => "11100110",2181 => "00111101",2182 => "11011001",2183 => "11000010",2184 => "11000011",2185 => "01100000",2186 => "11011001",2187 => "10000101",2188 => "11001010",2189 => "10001000",2190 => "01101000",2191 => "01101101",2192 => "01110001",2193 => "00100110",2194 => "11001000",2195 => "01111010",2196 => "11000110",2197 => "10010100",2198 => "01101100",2199 => "11011101",2200 => "11001001",2201 => "01001101",2202 => "11100000",2203 => "10011010",2204 => "01011110",2205 => "11111100",2206 => "10110011",2207 => "01000101",2208 => "00100010",2209 => "00110001",2210 => "10110100",2211 => "01110011",2212 => "10101101",2213 => "10001110",2214 => "11000000",2215 => "10001001",2216 => "11000110",2217 => "00100001",2218 => "00011011",2219 => "01011110",2220 => "01110101",2221 => "00110001",2222 => "00001100",2223 => "10001011",2224 => "00010101",2225 => "10011010",2226 => "00101101",2227 => "01001111",2228 => "10010110",2229 => "00111101",2230 => "10001101",2231 => "10111101",2232 => "11101011",2233 => "10111111",2234 => "10010011",2235 => "11011011",2236 => "10111011",2237 => "10001000",2238 => "00110110",2239 => "10000010",2240 => "01100001",2241 => "01100000",2242 => "11000111",2243 => "01000100",2244 => "01101001",2245 => "01101010",2246 => "01000001",2247 => "11100100",2248 => "10001100",2249 => "01100111",2250 => "10101000",2251 => "01000111",2252 => "01011000",2253 => "10000110",2254 => "10011110",2255 => "01010001",2256 => "01000110",2257 => "11101100",2258 => "10110010",2259 => "11101011",2260 => "00001100",2261 => "10100101",2262 => "11110110",2263 => "11101000",2264 => "11000111",2265 => "00100111",2266 => "11010110",2267 => "00000011",2268 => "11111100",2269 => "10001101",2270 => "11000010",2271 => "10010001",2272 => "10010010",2273 => "01110110",2274 => "11111111",2275 => "01101100",2276 => "01011001",2277 => "11101010",2278 => "01011001",2279 => "11001011",2280 => "10001010",2281 => "11001010",2282 => "11111001",2283 => "01100001",2284 => "01011101",2285 => "00110000",2286 => "01001001",2287 => "00010111",2288 => "01011110",2289 => "01110000",2290 => "01111010",2291 => "10010010",2292 => "11100101",2293 => "01110000",2294 => "01000111",2295 => "11000101",2296 => "10101101",2297 => "10100100",2298 => "10011000",2299 => "00000111",2300 => "00010000",2301 => "00100100",2302 => "11100011",2303 => "10101010",2304 => "01100010",2305 => "10011110",2306 => "00001000",2307 => "00111001",2308 => "10110001",2309 => "10010011",2310 => "11001011",2311 => "10010101",2312 => "11111110",2313 => "10110101",2314 => "01000100",2315 => "10100011",2316 => "01000111",2317 => "01110000",2318 => "00011100",2319 => "11110110",2320 => "10110100",2321 => "10010001",2322 => "10011110",2323 => "01001000",2324 => "01101100",2325 => "11001101",2326 => "11100000",2327 => "10101001",2328 => "00010110",2329 => "11110001",2330 => "11111010",2331 => "10100010",2332 => "11110100",2333 => "01001001",2334 => "00101110",2335 => "00111000",2336 => "01110000",2337 => "00111101",2338 => "11011001",2339 => "11110111",2340 => "00110000",2341 => "00111111",2342 => "01011110",2343 => "11110010",2344 => "00010010",2345 => "11111010",2346 => "11100101",2347 => "11100111",2348 => "11001010",2349 => "01000101",2350 => "10111100",2351 => "01111000",2352 => "00001011",2353 => "01011100",2354 => "11111100",2355 => "01110101",2356 => "10111100",2357 => "10011100",2358 => "01010001",2359 => "10101100",2360 => "00100110",2361 => "11101111",2362 => "00100000",2363 => "00111001",2364 => "11010111",2365 => "10110000",2366 => "11001010",2367 => "00010101",2368 => "10011000",2369 => "00100110",2370 => "11000110",2371 => "10111001",2372 => "00100010",2373 => "01101001",2374 => "11001100",2375 => "11000001",2376 => "01111111",2377 => "01010110",2378 => "10011100",2379 => "11001101",2380 => "11110100",2381 => "11101111",2382 => "01001110",2383 => "10010010",2384 => "00010001",2385 => "00010101",2386 => "11000001",2387 => "10000001",2388 => "01011010",2389 => "10000110",2390 => "10111100",2391 => "00110010",2392 => "00010100",2393 => "00010010",2394 => "01001100",2395 => "01111011",2396 => "11101100",2397 => "01010111",2398 => "11001110",2399 => "10000110",2400 => "10011000",2401 => "11111000",2402 => "10110100",2403 => "00001111",2404 => "00101001",2405 => "10011110",2406 => "01011001",2407 => "11111110",2408 => "10110101",2409 => "00011010",2410 => "10010110",2411 => "00100010",2412 => "01011100",2413 => "10111010",2414 => "11001010",2415 => "10010111",2416 => "11000101",2417 => "01100101",2418 => "01110010",2419 => "01011011",2420 => "10100010",2421 => "11001111",2422 => "00111111",2423 => "01100101",2424 => "11111100",2425 => "01010111",2426 => "00001010",2427 => "10110000",2428 => "01000110",2429 => "00111010",2430 => "00111100",2431 => "11100010",2432 => "00100000",2433 => "11111000",2434 => "11111110",2435 => "01000100",2436 => "10101100",2437 => "01011000",2438 => "01010100",2439 => "11111011",2440 => "01011110",2441 => "10111100",2442 => "11010111",2443 => "01011110",2444 => "11110001",2445 => "00010100",2446 => "11000100",2447 => "11000010",2448 => "10001010",2449 => "11011100",2450 => "10100011",2451 => "00000011",2452 => "11101101",2453 => "00101011",2454 => "10010100",2455 => "11001111",2456 => "00100000",2457 => "01110111",2458 => "01101101",2459 => "11110101",2460 => "11101001",2461 => "00111001",2462 => "11001110",2463 => "10111000",2464 => "00111110",2465 => "01100111",2466 => "10011011",2467 => "01010010",2468 => "01110010",2469 => "11100001",2470 => "01100100",2471 => "10100110",2472 => "01001010",2473 => "10111001",2474 => "11111000",2475 => "00100110",2476 => "00101000",2477 => "11110000",2478 => "11101111",2479 => "11011000",2480 => "11010001",2481 => "11110100",2482 => "11110000",2483 => "10001110",2484 => "11000011",2485 => "00000101",2486 => "00000110",2487 => "10111110",2488 => "10001111",2489 => "00010001",2490 => "11100011",2491 => "10110110",2492 => "10001010",2493 => "01110001",2494 => "11010101",2495 => "10011000",2496 => "10000001",2497 => "11000011",2498 => "01101011",2499 => "01010010",2500 => "10101011",2501 => "00100100",2502 => "10101001",2503 => "01010001",2504 => "11100111",2505 => "11001101",2506 => "10001111",2507 => "10011100",2508 => "10011110",2509 => "01001101",2510 => "01110001",2511 => "01100100",2512 => "11111001",2513 => "11101111",2514 => "01101000",2515 => "10001000",2516 => "11000001",2517 => "11001010",2518 => "11100100",2519 => "11001101",2520 => "01010100",2521 => "00101100",2522 => "10000111",2523 => "11010100",2524 => "10101100",2525 => "11111010",2526 => "00011001",2527 => "01010010",2528 => "11111011",2529 => "00100011",2530 => "00100111",2531 => "01001110",2532 => "10010111",2533 => "00000011",2534 => "00011100",2535 => "11010110",2536 => "11110011",2537 => "00111101",2538 => "00100010",2539 => "00101000",2540 => "10111111",2541 => "11010111",2542 => "01010100",2543 => "00011101",2544 => "00111000",2545 => "01101011",2546 => "01001101",2547 => "00100001",2548 => "10100010",2549 => "01111000",2550 => "11110010",2551 => "00101011",2552 => "01110010",2553 => "11011101",2554 => "00010101",2555 => "11111001",2556 => "10100101",2557 => "10101010",2558 => "11100101",2559 => "11001110",2560 => "10010001",2561 => "11001011",2562 => "11110110",2563 => "01101001",2564 => "10110000",2565 => "00011010",2566 => "11100011",2567 => "11000100",2568 => "11000100",2569 => "11111010",2570 => "11110101",2571 => "01111111",2572 => "01101101",2573 => "11110111",2574 => "00010011",2575 => "11000010",2576 => "11001111",2577 => "00111101",2578 => "01110111",2579 => "11000011",2580 => "10111001",2581 => "10001100",2582 => "11000110",2583 => "10011101",2584 => "10001101",2585 => "11110001",2586 => "11010011",2587 => "10100010",2588 => "00110110",2589 => "00000100",2590 => "11001110",2591 => "00000101",2592 => "00000110",2593 => "01110110",2594 => "00001000",2595 => "00001101",2596 => "10101111",2597 => "00011111",2598 => "10000011",2599 => "11011011",2600 => "01010101",2601 => "00011111",2602 => "00011111",2603 => "01100001",2604 => "11001101",2605 => "00001010",2606 => "01100110",2607 => "11001001",2608 => "10110010",2609 => "11001001",2610 => "00010010",2611 => "11000100",2612 => "00011111",2613 => "01101111",2614 => "01000010",2615 => "00111010",2616 => "11111000",2617 => "00010000",2618 => "01100010",2619 => "00101110",2620 => "00011100",2621 => "00000100",2622 => "10000110",2623 => "10111001",2624 => "10101001",2625 => "10001100",2626 => "11000111",2627 => "00001100",2628 => "11011011",2629 => "01010101",2630 => "00111011",2631 => "00011011",2632 => "01001101",2633 => "11110110",2634 => "10001011",2635 => "11011110",2636 => "11110011",2637 => "01101010",2638 => "01000000",2639 => "10110001",2640 => "10110100",2641 => "11110110",2642 => "01110110",2643 => "00111001",2644 => "00000100",2645 => "11101010",2646 => "11100100",2647 => "01001011",2648 => "00011001",2649 => "10110000",2650 => "00001100",2651 => "10110011",2652 => "00101111",2653 => "00110010",2654 => "11001101",2655 => "01111000",2656 => "10110101",2657 => "11110000",2658 => "00010100",2659 => "10110011",2660 => "00110111",2661 => "00100001",2662 => "00111010",2663 => "11000100",2664 => "10110000",2665 => "01110000",2666 => "00011000",2667 => "11010111",2668 => "10100101",2669 => "10000001",2670 => "01101011",2671 => "00110110",2672 => "01010111",2673 => "11100000",2674 => "10111100",2675 => "01011111",2676 => "11001001",2677 => "11011101",2678 => "01100000",2679 => "10110110",2680 => "01011001",2681 => "11111000",2682 => "01000001",2683 => "01101111",2684 => "11011101",2685 => "10100010",2686 => "01111010",2687 => "01110100",2688 => "00000000",2689 => "00100011",2690 => "11001001",2691 => "01111101",2692 => "00010001",2693 => "10000110",2694 => "01000001",2695 => "01011110",2696 => "00110010",2697 => "10010010",2698 => "10101100",2699 => "00000101",2700 => "00110000",2701 => "01101010",2702 => "10100100",2703 => "11111001",2704 => "11101001",2705 => "00010010",2706 => "00001111",2707 => "01000110",2708 => "10011110",2709 => "11011111",2710 => "00111111",2711 => "00010010",2712 => "00110010",2713 => "11001111",2714 => "01101100",2715 => "01001101",2716 => "10010001",2717 => "10101001",2718 => "00100110",2719 => "01001010",2720 => "01100001",2721 => "00101010",2722 => "00111010",2723 => "11000111",2724 => "11111001",2725 => "01000111",2726 => "00111101",2727 => "01101011",2728 => "10100010",2729 => "10111001",2730 => "01101101",2731 => "10100111",2732 => "11101011",2733 => "11101101",2734 => "00000110",2735 => "01011011",2736 => "01111110",2737 => "11001000",2738 => "10011111",2739 => "00101110",2740 => "10010010",2741 => "01011010",2742 => "11010000",2743 => "11100000",2744 => "01010100",2745 => "11000000",2746 => "11011100",2747 => "00101111",2748 => "00110110",2749 => "01000110",2750 => "01000111",2751 => "01011100",2752 => "01101011",2753 => "10101010",2754 => "00010011",2755 => "10101111",2756 => "10110001",2757 => "11001110",2758 => "10000001",2759 => "11001110",2760 => "11011101",2761 => "10010011",2762 => "11011010",2763 => "01000101",2764 => "10001010",2765 => "01010001",2766 => "10101001",2767 => "01110010",2768 => "11010101",2769 => "10001101",2770 => "10000100",2771 => "10101111",2772 => "01110011",2773 => "01000011",2774 => "10111110",2775 => "10101010",2776 => "00110110",2777 => "00010100",2778 => "01110110",2779 => "01111001",2780 => "10111010",2781 => "00010111",2782 => "11000000",2783 => "10001111",2784 => "11111010",2785 => "00101011",2786 => "10101100",2787 => "01001110",2788 => "00100010",2789 => "01000011",2790 => "11001110",2791 => "10010011",2792 => "01110010",2793 => "10111001",2794 => "10111100",2795 => "10111110",2796 => "00101000",2797 => "01100001",2798 => "01110101",2799 => "00100101",2800 => "00011101",2801 => "10001101",2802 => "00010101",2803 => "00100000",2804 => "00001001",2805 => "01001110",2806 => "11111110",2807 => "10111000",2808 => "00101100",2809 => "00011110",2810 => "10001010",2811 => "10011010",2812 => "01011011",2813 => "10000111",2814 => "10011101",2815 => "00010111",2816 => "11001011",2817 => "10000000",2818 => "10101001",2819 => "00110000",2820 => "00111100",2821 => "10000010",2822 => "11001010",2823 => "01111010",2824 => "11000110",2825 => "00010110",2826 => "00100101",2827 => "11100000",2828 => "01110001",2829 => "01000101",2830 => "01000111",2831 => "11000010",2832 => "11110011",2833 => "00000010",2834 => "11000111",2835 => "01011111",2836 => "00010001",2837 => "11010000",2838 => "10000111",2839 => "11010000",2840 => "11110111",2841 => "11000110",2842 => "00100110",2843 => "10110001",2844 => "11001110",2845 => "11010011",2846 => "00001110",2847 => "10011010",2848 => "00111011",2849 => "01010101",2850 => "10101001",2851 => "01100110",2852 => "01001011",2853 => "00110111",2854 => "11011001",2855 => "01110101",2856 => "00110000",2857 => "11111111",2858 => "01001100",2859 => "10101010",2860 => "10111101",2861 => "01111110",2862 => "10010111",2863 => "00111101",2864 => "00110110",2865 => "00000011",2866 => "10011111",2867 => "10001010",2868 => "10011110",2869 => "00110110",2870 => "01100101",2871 => "11000101",2872 => "11010000",2873 => "10101011",2874 => "10101100",2875 => "00000001",2876 => "11110010",2877 => "11011010",2878 => "11101111",2879 => "11111001",2880 => "00010111",2881 => "01100001",2882 => "00011101",2883 => "10110010",2884 => "11000100",2885 => "11111101",2886 => "01011110",2887 => "10111001",2888 => "01101001",2889 => "00111000",2890 => "01011001",2891 => "00011010",2892 => "11101101",2893 => "11000100",2894 => "10000000",2895 => "11111011",2896 => "10011010",2897 => "11010101",2898 => "01101000",2899 => "10011010",2900 => "10111100",2901 => "10110111",2902 => "11111000",2903 => "11111110",2904 => "11000000",2905 => "10111101",2906 => "11111010",2907 => "10110110",2908 => "10100010",2909 => "11001000",2910 => "01100100",2911 => "10000001",2912 => "00011111",2913 => "00011010",2914 => "11000110",2915 => "01101111",2916 => "00101010",2917 => "11111000",2918 => "11000001",2919 => "01111110",2920 => "10001000",2921 => "11101000",2922 => "01010001",2923 => "01101010",2924 => "10110111",2925 => "00101101",2926 => "01111001",2927 => "10110111",2928 => "10011010",2929 => "11011111",2930 => "11100110",2931 => "01111000",2932 => "00110001",2933 => "10111100",2934 => "11010001",2935 => "00000000",2936 => "11000010",2937 => "10110111",2938 => "11001111",2939 => "11011010",2940 => "01100110",2941 => "01110011",2942 => "00100111",2943 => "01000010",2944 => "01010001",2945 => "11000000",2946 => "10101100",2947 => "01100110",2948 => "11000010",2949 => "10011101",2950 => "00000100",2951 => "10111101",2952 => "00111001",2953 => "11100000",2954 => "01101011",2955 => "00100101",2956 => "01111011",2957 => "00010111",2958 => "11000000",2959 => "11100111",2960 => "01101000",2961 => "01111110",2962 => "01010111",2963 => "01111110",2964 => "11101111",2965 => "00010111",2966 => "00100100",2967 => "11111010",2968 => "11001111",2969 => "10000110",2970 => "10111111",2971 => "10100110",2972 => "11010001",2973 => "00100001",2974 => "00000000",2975 => "00010110",2976 => "01111110",2977 => "11110011",2978 => "11000010",2979 => "11101101",2980 => "01101001",2981 => "10110010",2982 => "11101001",2983 => "10111110",2984 => "00101000",2985 => "11001111",2986 => "11011100",2987 => "11010001",2988 => "10000101",2989 => "00000000",2990 => "11100010",2991 => "11111001",2992 => "10011001",2993 => "11000110",2994 => "10111000",2995 => "10111010",2996 => "11111100",2997 => "11110100",2998 => "00011010",2999 => "10000110",3000 => "00101010",3001 => "10001010",3002 => "10100011",3003 => "00111110",3004 => "00011101",3005 => "00110011",3006 => "11110010",3007 => "01000111",3008 => "10000000",3009 => "00100001",3010 => "10011100",3011 => "01110110",3012 => "11110000",3013 => "01111110",3014 => "01111000",3015 => "10101111",3016 => "11100000",3017 => "01000110",3018 => "11011001",3019 => "11111000",3020 => "00000010",3021 => "10100101",3022 => "11111100",3023 => "01011101",3024 => "11010000",3025 => "10100000",3026 => "10111000",3027 => "01001000",3028 => "11100011",3029 => "00011101",3030 => "11110001",3031 => "10110111",3032 => "00000100",3033 => "10111101",3034 => "00010101",3035 => "11111100",3036 => "01010010",3037 => "01110001",3038 => "11110101",3039 => "10111110",3040 => "11000011",3041 => "01010101",3042 => "10000011",3043 => "11110101",3044 => "01100010",3045 => "11111100",3046 => "11011001",3047 => "10111011",3048 => "11111110",3049 => "00100010",3050 => "11001000",3051 => "11110001",3052 => "10000010",3053 => "00001100",3054 => "00011011",3055 => "01010011",3056 => "01000101",3057 => "11010111",3058 => "00101111",3059 => "00111111",3060 => "00111010",3061 => "01001010",3062 => "11100100",3063 => "00000101",3064 => "10111000",3065 => "10010111",3066 => "11011001",3067 => "10100000",3068 => "00111011",3069 => "11001001",3070 => "11101100",3071 => "01010001",3072 => "10110011",3073 => "11011100",3074 => "11000111",3075 => "10011100",3076 => "10110111",3077 => "00011001",3078 => "00001100",3079 => "00011010",3080 => "00001101",3081 => "11010100",3082 => "01111101",3083 => "01110010",3084 => "10000010",3085 => "10101111",3086 => "11100001",3087 => "01110001",3088 => "00000110",3089 => "11001111",3090 => "00001100",3091 => "11111101",3092 => "11011111",3093 => "11101101",3094 => "00001100",3095 => "00101100",3096 => "01111001",3097 => "10001000",3098 => "11100010",3099 => "11001001",3100 => "11011101",3101 => "11000111",3102 => "01000000",3103 => "10110001",3104 => "01011100",3105 => "00100000",3106 => "01111001",3107 => "11101011",3108 => "00100000",3109 => "01110110",3110 => "10111101",3111 => "00000111",3112 => "10010011",3113 => "00111100",3114 => "01001101",3115 => "11100100",3116 => "01000110",3117 => "10000110",3118 => "11001001",3119 => "01100010",3120 => "00100010",3121 => "10101011",3122 => "10000010",3123 => "01111110",3124 => "01101011",3125 => "10110001",3126 => "00010010",3127 => "11001001",3128 => "10111100",3129 => "11001101",3130 => "11100100",3131 => "10010011",3132 => "10011001",3133 => "01000111",3134 => "01010001",3135 => "10110000",3136 => "10100010",3137 => "00000011",3138 => "10111000",3139 => "01100101",3140 => "10001001",3141 => "10111111",3142 => "00011101",3143 => "10101111",3144 => "00011000",3145 => "00010010",3146 => "00010000",3147 => "00111001",3148 => "00010010",3149 => "01001111",3150 => "01001100",3151 => "10111110",3152 => "00110110",3153 => "00010010",3154 => "11000100",3155 => "10100100",3156 => "00001100",3157 => "10101111",3158 => "11001001",3159 => "01011000",3160 => "00101101",3161 => "10000001",3162 => "11111111",3163 => "00011001",3164 => "01010100",3165 => "00011010",3166 => "10010101",3167 => "10000000",3168 => "01010101",3169 => "11101011",3170 => "10010001",3171 => "10000110",3172 => "10000011",3173 => "00001000",3174 => "10011001",3175 => "01110101",3176 => "01011111",3177 => "01010100",3178 => "11110001",3179 => "00100010",3180 => "11011010",3181 => "11010100",3182 => "10100111",3183 => "00111010",3184 => "01101111",3185 => "01001111",3186 => "11010101",3187 => "01100101",3188 => "10010011",3189 => "11111000",3190 => "00101111",3191 => "01110100",3192 => "01011001",3193 => "01101001",3194 => "00111010",3195 => "11101111",3196 => "01010110",3197 => "01101101",3198 => "00001000",3199 => "01111010",3200 => "11001010",3201 => "11011111",3202 => "10000110",3203 => "10101100",3204 => "10110011",3205 => "01101111",3206 => "00000000",3207 => "01100100",3208 => "11010011",3209 => "00010011",3210 => "10101000",3211 => "01000101",3212 => "10111110",3213 => "01110011",3214 => "11001100",3215 => "11110111",3216 => "01110010",3217 => "11100000",3218 => "00100100",3219 => "11101000",3220 => "11110111",3221 => "00110000",3222 => "00101000",3223 => "00101110",3224 => "00011000",3225 => "00101111",3226 => "11001110",3227 => "00010100",3228 => "11111001",3229 => "11000110",3230 => "10100000",3231 => "01011100",3232 => "10011000",3233 => "00011000",3234 => "01101000",3235 => "11110010",3236 => "00000001",3237 => "00110111",3238 => "11110110",3239 => "00000011",3240 => "00100101",3241 => "00011011",3242 => "01001000",3243 => "00001000",3244 => "00110101",3245 => "11111110",3246 => "01001110",3247 => "11000000",3248 => "00100000",3249 => "01000111",3250 => "00101010",3251 => "10111011",3252 => "10110011",3253 => "00011010",3254 => "10110100",3255 => "01111001",3256 => "10111000",3257 => "00011111",3258 => "00010101",3259 => "10111110",3260 => "11101010",3261 => "11000101",3262 => "11111100",3263 => "00101101",3264 => "00100100",3265 => "01110010",3266 => "11100000",3267 => "00000011",3268 => "00110101",3269 => "00110001",3270 => "00100111",3271 => "11100011",3272 => "11110111",3273 => "10110111",3274 => "11111001",3275 => "01000100",3276 => "10100010",3277 => "10010100",3278 => "00000010",3279 => "01101000",3280 => "00111010",3281 => "11000011",3282 => "11011110",3283 => "00011000",3284 => "00011001",3285 => "01001010",3286 => "10011000",3287 => "01110011",3288 => "11111010",3289 => "10000111",3290 => "11101001",3291 => "10100111",3292 => "10011010",3293 => "10010110",3294 => "10001011",3295 => "01010001",3296 => "11001010",3297 => "11101111",3298 => "00111001",3299 => "10111110",3300 => "01000010",3301 => "00101010",3302 => "10100010",3303 => "11001011",3304 => "10101101",3305 => "01010100",3306 => "11011011",3307 => "11100010",3308 => "00010011",3309 => "00000010",3310 => "11101111",3311 => "10000001",3312 => "10100101",3313 => "01010110",3314 => "10000111",3315 => "01111101",3316 => "10011010",3317 => "00001101",3318 => "00110111",3319 => "11101001",3320 => "10100000",3321 => "01001100",3322 => "01100110",3323 => "10001110",3324 => "01101111",3325 => "11010000",3326 => "00101010",3327 => "11000000",3328 => "00010100",3329 => "11111111",3330 => "01001011",3331 => "01001011",3332 => "10100110",3333 => "11100011",3334 => "10110100",3335 => "11001111",3336 => "11000100",3337 => "11000111",3338 => "00000111",3339 => "01001111",3340 => "01001011",3341 => "01101111",3342 => "01010000",3343 => "01101110",3344 => "10000000",3345 => "00001000",3346 => "01111111",3347 => "00010000",3348 => "10000111",3349 => "10110000",3350 => "01101100",3351 => "00010111",3352 => "01111000",3353 => "11001100",3354 => "11000001",3355 => "10101100",3356 => "11100111",3357 => "00110011",3358 => "00111011",3359 => "00100011",3360 => "11001010",3361 => "10111110",3362 => "00001001",3363 => "01001111",3364 => "11010001",3365 => "00111100",3366 => "00110100",3367 => "11100111",3368 => "00000101",3369 => "01000011",3370 => "10001101",3371 => "00111001",3372 => "00100100",3373 => "01000111",3374 => "00110000",3375 => "11011011",3376 => "01001011",3377 => "10001111",3378 => "01000010",3379 => "10000011",3380 => "01101000",3381 => "00101111",3382 => "00001010",3383 => "11001000",3384 => "00001010",3385 => "11111011",3386 => "00011101",3387 => "00100001",3388 => "10001011",3389 => "11101100",3390 => "11100100",3391 => "00100111",3392 => "01111101",3393 => "01001001",3394 => "10011101",3395 => "01000110",3396 => "00101101",3397 => "11010100",3398 => "11101110",3399 => "01010111",3400 => "00110111",3401 => "11000111",3402 => "10100111",3403 => "10000001",3404 => "01101110",3405 => "00110101",3406 => "11001011",3407 => "11000000",3408 => "01111011",3409 => "01110100",3410 => "11011111",3411 => "11010101",3412 => "10010111",3413 => "00001010",3414 => "00110111",3415 => "01110110",3416 => "10010010",3417 => "00101100",3418 => "00100000",3419 => "10011111",3420 => "01111011",3421 => "01010111",3422 => "01011000",3423 => "01000111",3424 => "11101101",3425 => "10111011",3426 => "00000110",3427 => "01110000",3428 => "01111011",3429 => "00010001",3430 => "10101111",3431 => "01011010",3432 => "11100000",3433 => "00101110",3434 => "00100110",3435 => "00110011",3436 => "10000111",3437 => "10101011",3438 => "11111011",3439 => "00110001",3440 => "00111010",3441 => "11111010",3442 => "10111000",3443 => "11000101",3444 => "11110111",3445 => "01100010",3446 => "00011100",3447 => "01111110",3448 => "10001100",3449 => "11010111",3450 => "00111001",3451 => "11110001",3452 => "11000011",3453 => "10101101",3454 => "00011001",3455 => "11101001",3456 => "10001001",3457 => "00000101",3458 => "10111111",3459 => "10010101",3460 => "11001101",3461 => "11111111",3462 => "10100101",3463 => "01101111",3464 => "10100101",3465 => "01101010",3466 => "01011001",3467 => "00001100",3468 => "10010101",3469 => "10101101",3470 => "00010111",3471 => "11100001",3472 => "10000101",3473 => "10011100",3474 => "00100100",3475 => "00101110",3476 => "00100001",3477 => "11000011",3478 => "01011110",3479 => "01110100",3480 => "11101100",3481 => "01001110",3482 => "11010010",3483 => "01101001",3484 => "01010000",3485 => "10010010",3486 => "01000101",3487 => "10111111",3488 => "01001000",3489 => "11010101",3490 => "10100000",3491 => "11010110",3492 => "11010001",3493 => "01010010",3494 => "00101101",3495 => "01111111",3496 => "11100101",3497 => "00000111",3498 => "10100110",3499 => "00001001",3500 => "11111110",3501 => "01111010",3502 => "10101110",3503 => "00010101",3504 => "11001101",3505 => "01100001",3506 => "01000011",3507 => "10010001",3508 => "10111101",3509 => "01011101",3510 => "10100110",3511 => "00000101",3512 => "01000101",3513 => "00110110",3514 => "01101100",3515 => "01110101",3516 => "01110101",3517 => "00100110",3518 => "10011000",3519 => "01001110",3520 => "11101010",3521 => "10000001",3522 => "00001111",3523 => "00010001",3524 => "10101101",3525 => "00000001",3526 => "11100101",3527 => "11111010",3528 => "10100000",3529 => "11110000",3530 => "00111110",3531 => "00010010",3532 => "10111000",3533 => "11000000",3534 => "01100010",3535 => "01000011",3536 => "00000101",3537 => "00111000",3538 => "00111001",3539 => "11110101",3540 => "10111000",3541 => "11100011",3542 => "01100011",3543 => "11001110",3544 => "01001101",3545 => "01111000",3546 => "01111110",3547 => "01010011",3548 => "11000011",3549 => "01100111",3550 => "10101010",3551 => "01100110",3552 => "11001101",3553 => "00000000",3554 => "00101110",3555 => "01001101",3556 => "00000111",3557 => "00101011",3558 => "10001001",3559 => "10100001",3560 => "11100101",3561 => "01101101",3562 => "10010011",3563 => "00000111",3564 => "01101011",3565 => "01000110",3566 => "10111111",3567 => "11010000",3568 => "00100001",3569 => "00110001",3570 => "11011110",3571 => "10110000",3572 => "10010110",3573 => "11000010",3574 => "01110010",3575 => "10001111",3576 => "11011110",3577 => "10011101",3578 => "10010011",3579 => "01010101",3580 => "10000000",3581 => "00011101",3582 => "00110101",3583 => "11001001",3584 => "11110000",3585 => "00111001",3586 => "11110110",3587 => "10111000",3588 => "00010100",3589 => "11011010",3590 => "10000100",3591 => "01010111",3592 => "10001100",3593 => "01101011",3594 => "11111011",3595 => "00000110",3596 => "00100001",3597 => "11000001",3598 => "00010110",3599 => "11100010",3600 => "01000101",3601 => "00100001",3602 => "10000100",3603 => "11001101",3604 => "00110101",3605 => "00110100",3606 => "11001101",3607 => "10011110",3608 => "00000100",3609 => "11001111",3610 => "11000111",3611 => "00110000",3612 => "01100110",3613 => "00111100",3614 => "01101110",3615 => "11100001",3616 => "01011010",3617 => "00001110",3618 => "11100110",3619 => "01011101",3620 => "01101011",3621 => "10010000",3622 => "00000110",3623 => "01000101",3624 => "01110110",3625 => "10010111",3626 => "00001010",3627 => "10011010",3628 => "01101110",3629 => "01111110",3630 => "10001011",3631 => "00111000",3632 => "10011110",3633 => "00000101",3634 => "10010110",3635 => "11011101",3636 => "01000100",3637 => "01000000",3638 => "10110001",3639 => "11100111",3640 => "11110011",3641 => "01000111",3642 => "00101110",3643 => "11001011",3644 => "01011110",3645 => "11000111",3646 => "11001110",3647 => "00110100",3648 => "01100101",3649 => "01101100",3650 => "11010110",3651 => "11000000",3652 => "01100011",3653 => "10000010",3654 => "01001010",3655 => "00100001",3656 => "00111110",3657 => "11111001",3658 => "11111001",3659 => "11111110",3660 => "01100001",3661 => "11111010",3662 => "10101010",3663 => "11001110",3664 => "10110110",3665 => "01011100",3666 => "00100010",3667 => "01101001",3668 => "10110010",3669 => "01101110",3670 => "01000111",3671 => "11101010",3672 => "10100110",3673 => "10111001",3674 => "01010101",3675 => "11110100",3676 => "00101101",3677 => "00010010",3678 => "11000101",3679 => "11101001",3680 => "11010100",3681 => "10111000",3682 => "11000101",3683 => "01010101",3684 => "11010101",3685 => "10110101",3686 => "11000111",3687 => "00010000",3688 => "11111111",3689 => "01101101",3690 => "11010011",3691 => "01111001",3692 => "01010001",3693 => "01111101",3694 => "10111001",3695 => "10111101",3696 => "01100001",3697 => "10110111",3698 => "10110111",3699 => "10100001",3700 => "00000011",3701 => "11010100",3702 => "00100011",3703 => "11110010",3704 => "10010001",3705 => "00011100",3706 => "11010110",3707 => "10100010",3708 => "10101100",3709 => "11001010",3710 => "00011100",3711 => "01101111",3712 => "01001100",3713 => "10110000",3714 => "10101001",3715 => "00001010",3716 => "11000100",3717 => "11010101",3718 => "10001001",3719 => "11111010",3720 => "01111111",3721 => "11010110",3722 => "01010010",3723 => "01001001",3724 => "10000011",3725 => "11010101",3726 => "01001010",3727 => "10001011",3728 => "10100001",3729 => "00111100",3730 => "00101001",3731 => "10100001",3732 => "01000110",3733 => "01011011",3734 => "01111111",3735 => "11001011",3736 => "10100011",3737 => "10110010",3738 => "10101001",3739 => "01000011",3740 => "11010010",3741 => "10010011",3742 => "10010101",3743 => "01000010",3744 => "01101100",3745 => "11000110",3746 => "00000010",3747 => "11010001",3748 => "00001110",3749 => "01011010",3750 => "01100001",3751 => "01100111",3752 => "01011011",3753 => "01000110",3754 => "00010101",3755 => "01111101",3756 => "00101010",3757 => "01001000",3758 => "00111011",3759 => "11111011",3760 => "00100111",3761 => "11001100",3762 => "11000101",3763 => "00101100",3764 => "01101110",3765 => "01001100",3766 => "01010000",3767 => "01011101",3768 => "01100111",3769 => "00100101",3770 => "10101010",3771 => "00101110",3772 => "01101001",3773 => "11001010",3774 => "00110100",3775 => "00100110",3776 => "01011010",3777 => "11000000",3778 => "00010100",3779 => "11000010",3780 => "01011010",3781 => "01001101",3782 => "11101110",3783 => "01110011",3784 => "00100000",3785 => "11101100",3786 => "11011011",3787 => "10111011",3788 => "10110000",3789 => "00111100",3790 => "01101100",3791 => "01011011",3792 => "01101111",3793 => "00011101",3794 => "00111111",3795 => "01101011",3796 => "11110111",3797 => "00110000",3798 => "11011001",3799 => "11011100",3800 => "01010100",3801 => "10111001",3802 => "10100000",3803 => "00000100",3804 => "11010100",3805 => "01010010",3806 => "00101110",3807 => "01111100",3808 => "11010000",3809 => "10010011",3810 => "01111101",3811 => "00100110",3812 => "01110111",3813 => "11110100",3814 => "00111100",3815 => "01000101",3816 => "01011010",3817 => "01011000",3818 => "10101001",3819 => "11110100",3820 => "01100001",3821 => "10001011",3822 => "11101100",3823 => "01101010",3824 => "11111010",3825 => "00110100",3826 => "10010000",3827 => "00001101",3828 => "10100100",3829 => "01111100",3830 => "11011010",3831 => "00011100",3832 => "01101010",3833 => "11010000",3834 => "01001111",3835 => "10100011",3836 => "10010001",3837 => "11000110",3838 => "00001001",3839 => "00000101",3840 => "10011011",3841 => "00110110",3842 => "00111001",3843 => "11001000",3844 => "01110010",3845 => "10001000",3846 => "00101110",3847 => "00111011",3848 => "11011110",3849 => "10100100",3850 => "00001011",3851 => "01011010",3852 => "11100100",3853 => "11001000",3854 => "00100101",3855 => "11110010",3856 => "00010010",3857 => "10110001",3858 => "10010101",3859 => "11101110",3860 => "10101001",3861 => "11111111",3862 => "00010110",3863 => "00111000",3864 => "11110001",3865 => "11000010",3866 => "11000101",3867 => "10011010",3868 => "00000011",3869 => "10101100",3870 => "00001100",3871 => "11011011",3872 => "10100000",3873 => "01110101",3874 => "10001100",3875 => "10010111",3876 => "11111101",3877 => "01111110",3878 => "10000101",3879 => "11011100",3880 => "10001011",3881 => "01010101",3882 => "01001011",3883 => "11011111",3884 => "11111011",3885 => "10011000",3886 => "10110000",3887 => "00011001",3888 => "01110101",3889 => "11110000",3890 => "11010110",3891 => "00100101",3892 => "00001101",3893 => "00100101",3894 => "11111000",3895 => "00110110",3896 => "10101100",3897 => "10111111",3898 => "11000100",3899 => "00100001",3900 => "00000110",3901 => "00111010",3902 => "00010001",3903 => "10110100",3904 => "01110100",3905 => "00100100",3906 => "01010110",3907 => "01011001",3908 => "11111100",3909 => "01100101",3910 => "01100100",3911 => "10010010",3912 => "11101001",3913 => "10011010",3914 => "00010100",3915 => "00001001",3916 => "10100000",3917 => "10010010",3918 => "11101010",3919 => "00001100",3920 => "10111100",3921 => "10000110",3922 => "11010000",3923 => "01010101",3924 => "10010100",3925 => "10010111",3926 => "10000110",3927 => "10001110",3928 => "11010101",3929 => "10000001",3930 => "11100000",3931 => "11111110",3932 => "00010111",3933 => "10101111",3934 => "00100011",3935 => "00110111",3936 => "01011100",3937 => "10100100",3938 => "11101101",3939 => "00111111",3940 => "00100010",3941 => "11100011",3942 => "00101011",3943 => "00110011",3944 => "11010101",3945 => "10001011",3946 => "01111010",3947 => "00000111",3948 => "11110100",3949 => "10000110",3950 => "00000111",3951 => "11110101",3952 => "11011000",3953 => "01000010",3954 => "10000001",3955 => "10111010",3956 => "00110100",3957 => "10100110",3958 => "01101001",3959 => "00011111",3960 => "01000110",3961 => "00011000",3962 => "01111011",3963 => "11110011",3964 => "10000001",3965 => "10010000",3966 => "00100110",3967 => "10101101",3968 => "01000110",3969 => "10010010",3970 => "11010001",3971 => "00101110",3972 => "11100010",3973 => "10101000",3974 => "00001100",3975 => "01110010",3976 => "01000101",3977 => "10010101",3978 => "00111110",3979 => "10111000",3980 => "11101000",3981 => "00100011",3982 => "00111111",3983 => "10111000",3984 => "00011010",3985 => "10000011",3986 => "00111000",3987 => "10101101",3988 => "00100100",3989 => "11110000",3990 => "01110011",3991 => "11000011",3992 => "00001011",3993 => "11011111",3994 => "01110000",3995 => "00001000",3996 => "00101110",3997 => "10000001",3998 => "01111010",3999 => "01011000",4000 => "10110000",4001 => "01100101",4002 => "11100101",4003 => "10111000",4004 => "10000001",4005 => "01011010",4006 => "11000101",4007 => "01010011",4008 => "11000001",4009 => "11100111",4010 => "00111001",4011 => "00100111",4012 => "11111010",4013 => "00001110",4014 => "10111010",4015 => "01011001",4016 => "10111011",4017 => "11001110",4018 => "00010010",4019 => "01011110",4020 => "00010101",4021 => "00110010",4022 => "11100101",4023 => "01001000",4024 => "01010001",4025 => "11110001",4026 => "10111110",4027 => "11111001",4028 => "10011010",4029 => "00101101",4030 => "10111011",4031 => "00110001",4032 => "01010010",4033 => "11110001",4034 => "11010011",4035 => "10101101",4036 => "11100111",4037 => "10101111",4038 => "01101111",4039 => "11100000",4040 => "10100010",4041 => "11011010",4042 => "00010010",4043 => "10110010",4044 => "10010000",4045 => "00110100",4046 => "01011101",4047 => "11011011",4048 => "00000100",4049 => "00011111",4050 => "00100110",4051 => "11111100",4052 => "00000010",4053 => "00100000",4054 => "00000000",4055 => "00111010",4056 => "01010100",4057 => "01010111",4058 => "11011100",4059 => "10000011",4060 => "00001000",4061 => "00100011",4062 => "01110110",4063 => "00011000",4064 => "10000101",4065 => "11111101",4066 => "11100110",4067 => "01100111",4068 => "11011010",4069 => "00001011",4070 => "01110111",4071 => "00001010",4072 => "01100001",4073 => "01010111",4074 => "11011110",4075 => "11110001",4076 => "00101100",4077 => "01000011",4078 => "11001100",4079 => "01110100",4080 => "01000011",4081 => "00001111",4082 => "10011110",4083 => "11110110",4084 => "01000001",4085 => "10001101",4086 => "11000000",4087 => "01111011",4088 => "10000111",4089 => "00111000",4090 => "00111110",4091 => "10010111",4092 => "01101111",4093 => "10001110",4094 => "00110001",4095 => "11001011",4096 => "01000011",4097 => "10101000",4098 => "10110011",4099 => "01100000",4100 => "11011010",4101 => "00010110",4102 => "10111011",4103 => "01010100",4104 => "11110101",4105 => "10111010",4106 => "00100000",4107 => "01000111",4108 => "10010110",4109 => "00100100",4110 => "11110111",4111 => "01111101",4112 => "00011110",4113 => "10101111",4114 => "10001100",4115 => "00101011",4116 => "11101001",4117 => "00110101",4118 => "11110001",4119 => "11101110",4120 => "11000111",4121 => "11011101",4122 => "00010010",4123 => "10100011",4124 => "00010001",4125 => "11000110",4126 => "10110011",4127 => "11110010",4128 => "01111111",4129 => "10011010",4130 => "11101100",4131 => "11101000",4132 => "00011010",4133 => "01100111",4134 => "01100000",4135 => "10110101",4136 => "00011011",4137 => "00001101",4138 => "10010100",4139 => "10110100",4140 => "11101001",4141 => "11110011",4142 => "01110101",4143 => "00001111",4144 => "00001110",4145 => "00101001",4146 => "00011001",4147 => "01101110",4148 => "10101111",4149 => "11011000",4150 => "00111101",4151 => "11001100",4152 => "10101100",4153 => "01000011",4154 => "00011110",4155 => "10100010",4156 => "00111111",4157 => "00111011",4158 => "11010001",4159 => "00100111",4160 => "01011011",4161 => "00111010",4162 => "00011110",4163 => "01001101",4164 => "00011000",4165 => "11011101",4166 => "10001101",4167 => "01100111",4168 => "00110111",4169 => "01100110",4170 => "01011101",4171 => "11010000",4172 => "10011010",4173 => "00011111",4174 => "00111111",4175 => "10111101",4176 => "11110010",4177 => "00010000",4178 => "01110010",4179 => "11011010",4180 => "01110011",4181 => "01101101",4182 => "10011110",4183 => "11110101",4184 => "10011000",4185 => "10111110",4186 => "01110000",4187 => "01010010",4188 => "01010110",4189 => "01101101",4190 => "01010000",4191 => "00100111",4192 => "11110010",4193 => "00101111",4194 => "01111011",4195 => "10110111",4196 => "10110110",4197 => "01010101",4198 => "11111110",4199 => "10000011",4200 => "11100110",4201 => "11011000",4202 => "10101100",4203 => "00101010",4204 => "11110101",4205 => "10110000",4206 => "01111101",4207 => "01011001",4208 => "10110010",4209 => "00101010",4210 => "11110101",4211 => "00101000",4212 => "11000011",4213 => "00111101",4214 => "01110111",4215 => "01011001",4216 => "01111100",4217 => "01010110",4218 => "11001010",4219 => "11010111",4220 => "00000000",4221 => "01001011",4222 => "11011101",4223 => "00101011",4224 => "11000100",4225 => "01010001",4226 => "00111001",4227 => "10110111",4228 => "01110001",4229 => "00001101",4230 => "00101110",4231 => "00100000",4232 => "00000111",4233 => "00110011",4234 => "00100010",4235 => "01101000",4236 => "00110111",4237 => "01001011",4238 => "11001000",4239 => "01110000",4240 => "01101110",4241 => "11001111",4242 => "10100000",4243 => "11110101",4244 => "01110110",4245 => "00100001",4246 => "11000100",4247 => "10011000",4248 => "10001100",4249 => "10101110",4250 => "10011110",4251 => "01010101",4252 => "11111010",4253 => "00010101",4254 => "11011111",4255 => "01000100",4256 => "01010101",4257 => "10010001",4258 => "00100101",4259 => "00110011",4260 => "00010001",4261 => "01101111",4262 => "01000001",4263 => "10001010",4264 => "11001010",4265 => "00011100",4266 => "11010000",4267 => "00110010",4268 => "00011011",4269 => "10010000",4270 => "01000011",4271 => "00000000",4272 => "11101000",4273 => "01101011",4274 => "01111111",4275 => "01111011",4276 => "00100011",4277 => "11000100",4278 => "00101011",4279 => "00111111",4280 => "10000001",4281 => "10011011",4282 => "10011100",4283 => "00011110",4284 => "10000000",4285 => "00111011",4286 => "11100110",4287 => "11101110",4288 => "00011001",4289 => "11100110",4290 => "01011110",4291 => "01011100",4292 => "01110111",4293 => "01100100",4294 => "10011100",4295 => "00011100",4296 => "11101111",4297 => "11010110",4298 => "10000111",4299 => "10011110",4300 => "01000110",4301 => "11011010",4302 => "01010100",4303 => "00110101",4304 => "10010000",4305 => "10111100",4306 => "00001110",4307 => "01010110",4308 => "11010000",4309 => "01010001",4310 => "00001011",4311 => "00000001",4312 => "11001010",4313 => "11000100",4314 => "10100101",4315 => "00010101",4316 => "00010011",4317 => "10001011",4318 => "10110100",4319 => "01010000",4320 => "01110001",4321 => "10000101",4322 => "10111111",4323 => "01111010",4324 => "01111010",4325 => "10101110",4326 => "11111110",4327 => "11010000",4328 => "10001100",4329 => "00101011",4330 => "00000011",4331 => "01001000",4332 => "01111000",4333 => "10000101",4334 => "11100110",4335 => "11110011",4336 => "10011001",4337 => "11000001",4338 => "11010011",4339 => "00110010",4340 => "01100001",4341 => "01111110",4342 => "00110011",4343 => "10100111",4344 => "10000000",4345 => "10000011",4346 => "00000101",4347 => "01110110",4348 => "00111110",4349 => "10011100",4350 => "11100101",4351 => "01000101",4352 => "11010110",4353 => "11000111",4354 => "01011100",4355 => "00100001",4356 => "11111001",4357 => "10111011",4358 => "10001111",4359 => "10000001",4360 => "11111001",4361 => "00011001",4362 => "11001110",4363 => "10001111",4364 => "01000010",4365 => "11111001",4366 => "11010101",4367 => "11111100",4368 => "10101010",4369 => "11110000",4370 => "11000101",4371 => "00100111",4372 => "10000100",4373 => "01100001",4374 => "11001000",4375 => "00010000",4376 => "10111001",4377 => "00001111",4378 => "11010101",4379 => "11000010",4380 => "11100010",4381 => "10111100",4382 => "00110011",4383 => "00101110",4384 => "00111001",4385 => "10011100",4386 => "00110101",4387 => "10000110",4388 => "00000010",4389 => "01101111",4390 => "11111101",4391 => "11001111",4392 => "00000010",4393 => "10000011",4394 => "01011100",4395 => "10101000",4396 => "00100100",4397 => "10001101",4398 => "00111011",4399 => "01011000",4400 => "00100110",4401 => "01001110",4402 => "01000111",4403 => "00110010",4404 => "00101111",4405 => "10111100",4406 => "01110100",4407 => "11111111",4408 => "11000101",4409 => "11011110",4410 => "00011011",4411 => "11000110",4412 => "00111100",4413 => "00000101",4414 => "11000011",4415 => "11101001",4416 => "01000010",4417 => "00001111",4418 => "00001010",4419 => "00010101",4420 => "01110001",4421 => "01010001",4422 => "00110010",4423 => "11010000",4424 => "11100100",4425 => "01010000",4426 => "10111000",4427 => "01000011",4428 => "10011101",4429 => "11011010",4430 => "11000000",4431 => "10101001",4432 => "11101001",4433 => "11110111",4434 => "01100101",4435 => "01011000",4436 => "11010001",4437 => "00000111",4438 => "00100011",4439 => "10100011",4440 => "10100010",4441 => "11011100",4442 => "11100010",4443 => "00011100",4444 => "00011011",4445 => "00001100",4446 => "01010001",4447 => "00001010",4448 => "00001101",4449 => "10100001",4450 => "10111000",4451 => "00100010",4452 => "11011110",4453 => "00100110",4454 => "01101111",4455 => "10011010",4456 => "01000111",4457 => "00010110",4458 => "10111001",4459 => "00011111",4460 => "00111111",4461 => "10010101",4462 => "10100101",4463 => "00001001",4464 => "01101011",4465 => "00001000",4466 => "10001110",4467 => "10001010",4468 => "10110101",4469 => "01110001",4470 => "10010101",4471 => "00111100",4472 => "11000010",4473 => "11101111",4474 => "11011110",4475 => "01000011",4476 => "00110111",4477 => "01100100",4478 => "10110100",4479 => "00100110",4480 => "00011010",4481 => "10001001",4482 => "01110101",4483 => "01011000",4484 => "01101111",4485 => "00101011",4486 => "01010101",4487 => "00000100",4488 => "01011110",4489 => "11011101",4490 => "01110101",4491 => "10011110",4492 => "11101100",4493 => "10100110",4494 => "10100101",4495 => "01100001",4496 => "11111001",4497 => "10110101",4498 => "00110010",4499 => "11011110",4500 => "00001011",4501 => "01101110",4502 => "01001110",4503 => "10000010",4504 => "11000001",4505 => "10110001",4506 => "11101111",4507 => "10111100",4508 => "10011000",4509 => "11000110",4510 => "10001001",4511 => "00010110",4512 => "10100000",4513 => "00101111",4514 => "11001000",4515 => "10000001",4516 => "11110010",4517 => "10100010",4518 => "00110101",4519 => "10100110",4520 => "01101110",4521 => "11001110",4522 => "01100110",4523 => "01100001",4524 => "11010010",4525 => "11101110",4526 => "00000000",4527 => "00100000",4528 => "00000011",4529 => "11111110",4530 => "01100110",4531 => "10111011",4532 => "10010100",4533 => "00110000",4534 => "11111111",4535 => "01010110",4536 => "00101111",4537 => "01001000",4538 => "00110010",4539 => "01110110",4540 => "00000000",4541 => "01110011",4542 => "11000111",4543 => "01000000",4544 => "00110001",4545 => "11111101",4546 => "00001111",4547 => "11110000",4548 => "01111000",4549 => "10101110",4550 => "10100010",4551 => "10101010",4552 => "10111101",4553 => "10100111",4554 => "11100010",4555 => "00101111",4556 => "11101010",4557 => "00011110",4558 => "00110011",4559 => "00000111",4560 => "01011001",4561 => "10000101",4562 => "11011011",4563 => "10011111",4564 => "10000111",4565 => "10101101",4566 => "01010100",4567 => "00110010",4568 => "10001010",4569 => "01101110",4570 => "10001111",4571 => "10110101",4572 => "10110111",4573 => "11100111",4574 => "10111101",4575 => "10110011",4576 => "00001011",4577 => "10011110",4578 => "10010110",4579 => "10101110",4580 => "00011101",4581 => "00100000",4582 => "10001010",4583 => "10001000",4584 => "10100101",4585 => "00101011",4586 => "01110000",4587 => "10110011",4588 => "00010100",4589 => "10111110",4590 => "11101100",4591 => "00100100",4592 => "10100001",4593 => "01110101",4594 => "11111001",4595 => "10101101",4596 => "01011000",4597 => "01011110",4598 => "01101001",4599 => "01011000",4600 => "11100101",4601 => "11010100",4602 => "00111001",4603 => "11001110",4604 => "00100010",4605 => "00110111",4606 => "00001001",4607 => "10110001",4608 => "10100110",4609 => "00100101",4610 => "00101101",4611 => "00000101",4612 => "00000001",4613 => "11001011",4614 => "10010100",4615 => "00100000",4616 => "00011011",4617 => "10001001",4618 => "01101101",4619 => "11100001",4620 => "01101101",4621 => "11100111",4622 => "11100111",4623 => "00101101",4624 => "11010100",4625 => "10011100",4626 => "00010101",4627 => "11110100",4628 => "11100001",4629 => "00111000",4630 => "11100101",4631 => "01111111",4632 => "10001000",4633 => "00010110",4634 => "00110111",4635 => "01110100",4636 => "01001110",4637 => "01000011",4638 => "00000000",4639 => "00001101",4640 => "01010101",4641 => "00001011",4642 => "11111111",4643 => "01110111",4644 => "00010110",4645 => "00100101",4646 => "00100110",4647 => "11110011",4648 => "11111100",4649 => "00001001",4650 => "01100010",4651 => "10110010",4652 => "00011011",4653 => "01000000",4654 => "11011111",4655 => "00011001",4656 => "01111001",4657 => "01010100",4658 => "00101011",4659 => "11100001",4660 => "01111010",4661 => "10000001",4662 => "01001010",4663 => "11111101",4664 => "01010110",4665 => "01001111",4666 => "00110011",4667 => "10101111",4668 => "01100011",4669 => "00001101",4670 => "01010111",4671 => "10000100",4672 => "01011000",4673 => "11000011",4674 => "11100000",4675 => "11111110",4676 => "10001101",4677 => "01000100",4678 => "10000010",4679 => "00100010",4680 => "11100001",4681 => "00010010",4682 => "10000000",4683 => "10111011",4684 => "01111111",4685 => "00001001",4686 => "00001001",4687 => "00001101",4688 => "10000101",4689 => "00110001",4690 => "11001111",4691 => "10111011",4692 => "00011110",4693 => "10110100",4694 => "10000000",4695 => "11001010",4696 => "01101111",4697 => "01110100",4698 => "00000101",4699 => "10011010",4700 => "10110110",4701 => "00100111",4702 => "11000000",4703 => "01111101",4704 => "01001000",4705 => "01101010",4706 => "00111011",4707 => "00010010",4708 => "01010110",4709 => "00100101",4710 => "00001100",4711 => "11011001",4712 => "11101010",4713 => "11111001",4714 => "10001100",4715 => "01110100",4716 => "10110111",4717 => "11001000",4718 => "00110001",4719 => "00100110",4720 => "10000000",4721 => "00000010",4722 => "10010101",4723 => "10001101",4724 => "11110100",4725 => "01010010",4726 => "11101000",4727 => "00111101",4728 => "10010011",4729 => "00101101",4730 => "10110110",4731 => "01010001",4732 => "11110010",4733 => "01011110",4734 => "10010111",4735 => "10100010",4736 => "10110010",4737 => "10111000",4738 => "10000101",4739 => "10011001",4740 => "01111001",4741 => "01010110",4742 => "10001111",4743 => "00000000",4744 => "01100100",4745 => "11000001",4746 => "01000011",4747 => "10100100",4748 => "01010001",4749 => "11101100",4750 => "10110010",4751 => "00010000",4752 => "01001000",4753 => "11001100",4754 => "10000001",4755 => "00100101",4756 => "11001001",4757 => "00001001",4758 => "11100111",4759 => "00100011",4760 => "11101001",4761 => "01110111",4762 => "01110100",4763 => "10001110",4764 => "01001000",4765 => "00111011",4766 => "10000101",4767 => "11100010",4768 => "01011100",4769 => "10010010",4770 => "00001110",4771 => "00110110",4772 => "00101111",4773 => "11001101",4774 => "00000001",4775 => "10110010",4776 => "00010101",4777 => "01010010",4778 => "01001111",4779 => "11110010",4780 => "01001110",4781 => "01001110",4782 => "11000000",4783 => "11011010",4784 => "00011000",4785 => "11100111",4786 => "11110101",4787 => "11001101",4788 => "11000000",4789 => "11110110",4790 => "01100000",4791 => "01010001",4792 => "00111110",4793 => "11101111",4794 => "11100010",4795 => "11110001",4796 => "11110010",4797 => "00001101",4798 => "00110101",4799 => "10101010",4800 => "01010110",4801 => "00001111",4802 => "01100101",4803 => "00101111",4804 => "10110100",4805 => "11001010",4806 => "11110111",4807 => "11010000",4808 => "01110011",4809 => "01101100",4810 => "00100111",4811 => "01111111",4812 => "10110011",4813 => "01101110",4814 => "01111101",4815 => "00110100",4816 => "11001011",4817 => "01011001",4818 => "00011101",4819 => "10010000",4820 => "01001111",4821 => "01001110",4822 => "00000111",4823 => "11000111",4824 => "00110100",4825 => "01010101",4826 => "01101010",4827 => "11011011",4828 => "01110010",4829 => "11111000",4830 => "11001010",4831 => "00011001",4832 => "10111111",4833 => "11001011",4834 => "11111010",4835 => "01110101",4836 => "10111000",4837 => "00101010",4838 => "01101010",4839 => "10001110",4840 => "11110000",4841 => "00111111",4842 => "00000010",4843 => "11001000",4844 => "00001101",4845 => "00100000",4846 => "00000001",4847 => "11101010",4848 => "11111011",4849 => "10110100",4850 => "00010010",4851 => "11011010",4852 => "11011011",4853 => "11011100",4854 => "11100000",4855 => "10000010",4856 => "00011111",4857 => "01100100",4858 => "01001011",4859 => "00101101",4860 => "11010010",4861 => "10011000",4862 => "00100011",4863 => "10010001",4864 => "10101010",4865 => "00001100",4866 => "01110001",4867 => "11111100",4868 => "00101111",4869 => "11100101",4870 => "01101010",4871 => "11001101",4872 => "01001000",4873 => "11101110",4874 => "11101011",4875 => "01100101",4876 => "00011000",4877 => "11110110",4878 => "10000101",4879 => "00000000",4880 => "10000011",4881 => "00110110",4882 => "10111000",4883 => "01100100",4884 => "10000000",4885 => "01100001",4886 => "01000111",4887 => "00111010",4888 => "00100100",4889 => "01001011",4890 => "01100111",4891 => "11000011",4892 => "01100101",4893 => "11111011",4894 => "00000010",4895 => "10100011",4896 => "00100011",4897 => "00011001",4898 => "11111100",4899 => "00010010",4900 => "10000011",4901 => "00110100",4902 => "11010111",4903 => "00100011",4904 => "01101110",4905 => "11001000",4906 => "10011010",4907 => "10011001",4908 => "11001111",4909 => "10111001",4910 => "00100100",4911 => "10011100",4912 => "00110101",4913 => "11011111",4914 => "11100110",4915 => "10011011",4916 => "10111110",4917 => "01010011",4918 => "10011111",4919 => "00101110",4920 => "01011101",4921 => "10111111",4922 => "01110011",4923 => "00011011",4924 => "01111001",4925 => "11111110",4926 => "01001100",4927 => "11101110",4928 => "10010111",4929 => "10100001",4930 => "01111011",4931 => "10010100",4932 => "11011001",4933 => "00010010",4934 => "01010111",4935 => "00000101",4936 => "00101100",4937 => "01001101",4938 => "11101111",4939 => "11011100",4940 => "01001000",4941 => "11010001",4942 => "10001001",4943 => "00000000",4944 => "11110011",4945 => "00001010",4946 => "10101110",4947 => "01110101",4948 => "01110111",4949 => "00111010",4950 => "01001110",4951 => "11100111",4952 => "01010110",4953 => "11111110",4954 => "10101110",4955 => "11011111",4956 => "00010010",4957 => "01110111",4958 => "11111101",4959 => "01101000",4960 => "01001111",4961 => "10100001",4962 => "10010100",4963 => "00111010",4964 => "00011101",4965 => "01111010",4966 => "01101010",4967 => "11101101",4968 => "11001001",4969 => "10001111",4970 => "11001000",4971 => "01000101",4972 => "00001111",4973 => "10001000",4974 => "10001111",4975 => "00011111",4976 => "01001111",4977 => "11111011",4978 => "01110010",4979 => "11001010",4980 => "11110100",4981 => "11001000",4982 => "00001100",4983 => "10111001",4984 => "01011110",4985 => "01101111",4986 => "10001000",4987 => "11101100",4988 => "01000000",4989 => "10111001",4990 => "11100001",4991 => "10100110",4992 => "01101100",4993 => "10000110",4994 => "11101100",4995 => "00001001",4996 => "10100000",4997 => "11001010",4998 => "11010110",4999 => "01100101",5000 => "01110000",5001 => "00101000",5002 => "01110000",5003 => "01110111",5004 => "11100000",5005 => "01001110",5006 => "01100101",5007 => "10110100",5008 => "11100101",5009 => "01110100",5010 => "11010011",5011 => "01000101",5012 => "10100100",5013 => "11001010",5014 => "00100111",5015 => "10101111",5016 => "11000110",5017 => "00101010",5018 => "00111001",5019 => "01110010",5020 => "00010001",5021 => "10011111",5022 => "00011100",5023 => "01010010",5024 => "01011010",5025 => "10001010",5026 => "01100001",5027 => "01011001",5028 => "00111100",5029 => "10100000",5030 => "00100011",5031 => "11001000",5032 => "01001011",5033 => "11111000",5034 => "10101000",5035 => "11110011",5036 => "00111000",5037 => "10001110",5038 => "10011001",5039 => "00010010",5040 => "10011010",5041 => "01001100",5042 => "01100011",5043 => "00011100",5044 => "00111001",5045 => "01000111",5046 => "01010100",5047 => "01000011",5048 => "10011001",5049 => "01010101",5050 => "01011111",5051 => "10101000",5052 => "01001100",5053 => "11010100",5054 => "01101110",5055 => "00011000",5056 => "11111010",5057 => "11000101",5058 => "11001001",5059 => "11110110",5060 => "01011111",5061 => "11111111",5062 => "00000010",5063 => "01000000",5064 => "11011111",5065 => "01110111",5066 => "11101001",5067 => "10101011",5068 => "11110011",5069 => "11100001",5070 => "11101100",5071 => "10011011",5072 => "00000110",5073 => "00110000",5074 => "10000011",5075 => "00110101",5076 => "10000010",5077 => "01110101",5078 => "11111010",5079 => "10111100",5080 => "11101001",5081 => "10010011",5082 => "01001000",5083 => "10001101",5084 => "00001001",5085 => "00000101",5086 => "10111101",5087 => "11100011",5088 => "10111011",5089 => "10101100",5090 => "00000110",5091 => "11110110",5092 => "01000111",5093 => "00001010",5094 => "10110111",5095 => "00100001",5096 => "11000000",5097 => "00110001",5098 => "00100000",5099 => "10100110",5100 => "00101011",5101 => "00100010",5102 => "01001011",5103 => "10111101",5104 => "11110101",5105 => "01110001",5106 => "11001101",5107 => "11101000",5108 => "01101110",5109 => "01001111",5110 => "00110110",5111 => "00001111",5112 => "01001101",5113 => "00011100",5114 => "00011000",5115 => "00011100",5116 => "11110011",5117 => "01110001",5118 => "01100111",5119 => "01000011",5120 => "10011011",5121 => "01001100",5122 => "00011111",5123 => "10001001",5124 => "00001011",5125 => "00111111",5126 => "10011111",5127 => "11101100",5128 => "11101111",5129 => "00011001",5130 => "01111101",5131 => "00100000",5132 => "11101001",5133 => "11100000",5134 => "11000011",5135 => "01101110",5136 => "11010100",5137 => "10110100",5138 => "01011011",5139 => "10110100",5140 => "11010101",5141 => "01111101",5142 => "01110001",5143 => "01110111",5144 => "01110110",5145 => "01101110",5146 => "00001001",5147 => "10001011",5148 => "11000010",5149 => "10111100",5150 => "01000110",5151 => "00000010",5152 => "00101110",5153 => "00101101",5154 => "00011100",5155 => "11011110",5156 => "01010110",5157 => "10110101",5158 => "01000110",5159 => "00001001",5160 => "10111011",5161 => "11001101",5162 => "01110010",5163 => "00010001",5164 => "10100111",5165 => "00000111",5166 => "01000000",5167 => "10011111",5168 => "11011100",5169 => "11110100",5170 => "01110000",5171 => "11110100",5172 => "01010101",5173 => "10011111",5174 => "10011010",5175 => "01000100",5176 => "11011111",5177 => "10001100",5178 => "01010110",5179 => "10000000",5180 => "10110010",5181 => "01111011",5182 => "11101101",5183 => "01000010",5184 => "11100100",5185 => "11011010",5186 => "11011101",5187 => "01110001",5188 => "10000011",5189 => "11111101",5190 => "01011100",5191 => "01101111",5192 => "01111110",5193 => "01101011",5194 => "01110101",5195 => "01111001",5196 => "11110110",5197 => "01111011",5198 => "01110111",5199 => "01100010",5200 => "11110111",5201 => "11010011",5202 => "01110010",5203 => "10111110",5204 => "00101101",5205 => "11111100",5206 => "01000111",5207 => "00001111",5208 => "10100110",5209 => "10101101",5210 => "11010110",5211 => "10010000",5212 => "01010100",5213 => "00001110",5214 => "01100111",5215 => "11101110",5216 => "01100011",5217 => "11100101",5218 => "00110001",5219 => "10101111",5220 => "10110010",5221 => "00010111",5222 => "11000111",5223 => "11010110",5224 => "11000111",5225 => "01111010",5226 => "11010011",5227 => "01111011",5228 => "01001011",5229 => "01001100",5230 => "11011011",5231 => "01101010",5232 => "10101010",5233 => "10010010",5234 => "10101100",5235 => "00001100",5236 => "11110111",5237 => "11011001",5238 => "11110100",5239 => "00100111",5240 => "00010010",5241 => "10011110",5242 => "10100011",5243 => "11110110",5244 => "00110100",5245 => "10101001",5246 => "01010100",5247 => "00001010",5248 => "11000000",5249 => "10110101",5250 => "01000100",5251 => "01001100",5252 => "10001010",5253 => "01010010",5254 => "00100011",5255 => "10001011",5256 => "00001100",5257 => "01011111",5258 => "10000011",5259 => "00010000",5260 => "01100111",5261 => "11001000",5262 => "00111100",5263 => "11110011",5264 => "11011100",5265 => "00101011",5266 => "10000001",5267 => "00000001",5268 => "11000001",5269 => "10011000",5270 => "11111001",5271 => "10110000",5272 => "00011001",5273 => "11110111",5274 => "10000101",5275 => "10010110",5276 => "00000001",5277 => "01111011",5278 => "00101010",5279 => "10110101",5280 => "00100010",5281 => "00110101",5282 => "11010010",5283 => "10110101",5284 => "01110001",5285 => "11000000",5286 => "01100100",5287 => "11010101",5288 => "11011011",5289 => "01010001",5290 => "00010011",5291 => "00110110",5292 => "01110000",5293 => "01111101",5294 => "01110111",5295 => "00011100",5296 => "11101101",5297 => "01100000",5298 => "00001011",5299 => "10111111",5300 => "11011101",5301 => "00110011",5302 => "01110101",5303 => "00110110",5304 => "01111011",5305 => "00000000",5306 => "00110000",5307 => "01111100",5308 => "01101010",5309 => "01100111",5310 => "11111111",5311 => "10100000",5312 => "01011111",5313 => "01001001",5314 => "01111111",5315 => "00000110",5316 => "10000101",5317 => "01111110",5318 => "11001111",5319 => "01100101",5320 => "11111010",5321 => "10100101",5322 => "10010001",5323 => "00110101",5324 => "00001101",5325 => "10111000",5326 => "00111111",5327 => "11010010",5328 => "01111100",5329 => "01011001",5330 => "01101101",5331 => "00101101",5332 => "00100110",5333 => "00001000",5334 => "00000101",5335 => "01101011",5336 => "00011001",5337 => "10101111",5338 => "00010011",5339 => "00100101",5340 => "01000011",5341 => "11000101",5342 => "01010010",5343 => "01101101",5344 => "11001100",5345 => "01100000",5346 => "11101000",5347 => "01111111",5348 => "00100011",5349 => "01110111",5350 => "01111100",5351 => "11110011",5352 => "11001100",5353 => "11010101",5354 => "11010100",5355 => "00111101",5356 => "11000000",5357 => "11101000",5358 => "01111000",5359 => "11110000",5360 => "10100110",5361 => "01010101",5362 => "01100111",5363 => "01110011",5364 => "11011100",5365 => "00100110",5366 => "11010011",5367 => "11001100",5368 => "01101111",5369 => "01010010",5370 => "10111111",5371 => "10111001",5372 => "10001101",5373 => "10100011",5374 => "01011010",5375 => "11010001",5376 => "00011001",5377 => "00010110",5378 => "11011110",5379 => "11111000",5380 => "10001111",5381 => "11010000",5382 => "10010011",5383 => "10111011",5384 => "11101011",5385 => "11110011",5386 => "11001101",5387 => "00010000",5388 => "10001101",5389 => "10111101",5390 => "10001011",5391 => "11001101",5392 => "01101100",5393 => "11100101",5394 => "00100110",5395 => "11110110",5396 => "00001100",5397 => "01000010",5398 => "11011000",5399 => "10010111",5400 => "10100010",5401 => "11101011",5402 => "10011100",5403 => "11001011",5404 => "00000101",5405 => "01010101",5406 => "10101110",5407 => "10001010",5408 => "00000001",5409 => "11111001",5410 => "00011001",5411 => "10101010",5412 => "01010110",5413 => "10011000",5414 => "01011101",5415 => "01101110",5416 => "00110110",5417 => "11000111",5418 => "00010011",5419 => "00010110",5420 => "10001101",5421 => "01000111",5422 => "01001001",5423 => "01110001",5424 => "10011111",5425 => "00101010",5426 => "11000100",5427 => "01100101",5428 => "01010111",5429 => "00000011",5430 => "11100000",5431 => "11001111",5432 => "10101111",5433 => "10001000",5434 => "00011111",5435 => "10001111",5436 => "00010010",5437 => "00100100",5438 => "10010110",5439 => "11011100",5440 => "00100110",5441 => "11011011",5442 => "11011000",5443 => "10010101",5444 => "00000100",5445 => "01101001",5446 => "11101101",5447 => "10101011",5448 => "11011101",5449 => "00101101",5450 => "00110101",5451 => "00000000",5452 => "00110011",5453 => "10110010",5454 => "01100010",5455 => "00100101",5456 => "01101111",5457 => "01110001",5458 => "01111101",5459 => "00011001",5460 => "01101110",5461 => "00101010",5462 => "11001110",5463 => "10001101",5464 => "11001101",5465 => "10010011",5466 => "00010100",5467 => "01100010",5468 => "10100111",5469 => "11110101",5470 => "00001110",5471 => "10011100",5472 => "00111110",5473 => "11110100",5474 => "01111111",5475 => "10110001",5476 => "10111001",5477 => "10001000",5478 => "11101110",5479 => "11101011",5480 => "00101100",5481 => "01110000",5482 => "11010010",5483 => "10001110",5484 => "01001011",5485 => "01100011",5486 => "01000111",5487 => "11001100",5488 => "01100111",5489 => "00000010",5490 => "00110000",5491 => "00000011",5492 => "01101110",5493 => "01010001",5494 => "00000011",5495 => "11001101",5496 => "10111010",5497 => "00110010",5498 => "01111000",5499 => "00110010",5500 => "00010010",5501 => "11010010",5502 => "10110101",5503 => "10101101",5504 => "11110000",5505 => "01010000",5506 => "01000101",5507 => "10101000",5508 => "00011010",5509 => "10000010",5510 => "11100000",5511 => "00001001",5512 => "00011000",5513 => "11010011",5514 => "01110100",5515 => "10101110",5516 => "00100110",5517 => "00010100",5518 => "10100100",5519 => "00001000",5520 => "10100000",5521 => "00000101",5522 => "11101001",5523 => "01101011",5524 => "00001110",5525 => "11100000",5526 => "00110110",5527 => "11110001",5528 => "00110110",5529 => "10001110",5530 => "11011100",5531 => "01101001",5532 => "01110011",5533 => "01000011",5534 => "11111110",5535 => "10100100",5536 => "11011010",5537 => "00100011",5538 => "00101010",5539 => "11101101",5540 => "00100101",5541 => "01001001",5542 => "01100001",5543 => "01010100",5544 => "11110000",5545 => "10101011",5546 => "01001011",5547 => "11001010",5548 => "10110100",5549 => "00110000",5550 => "10010010",5551 => "01011101",5552 => "00010000",5553 => "10001010",5554 => "01010110",5555 => "01001001",5556 => "01011001",5557 => "10111100",5558 => "10101111",5559 => "10011010",5560 => "01000010",5561 => "01110100",5562 => "00011001",5563 => "00100110",5564 => "01010000",5565 => "11011000",5566 => "11011100",5567 => "01001011",5568 => "11101101",5569 => "00100010",5570 => "01101000",5571 => "11100101",5572 => "01001000",5573 => "10001100",5574 => "11110000",5575 => "11010001",5576 => "00100000",5577 => "00100111",5578 => "00001100",5579 => "11011011",5580 => "10010101",5581 => "00100101",5582 => "10101100",5583 => "01110110",5584 => "11000011",5585 => "00101000",5586 => "01110011",5587 => "11100110",5588 => "00101101",5589 => "00111010",5590 => "01001011",5591 => "10100010",5592 => "00111100",5593 => "01111001",5594 => "00000011",5595 => "01000100",5596 => "11111100",5597 => "01010001",5598 => "01100011",5599 => "01010010",5600 => "11111011",5601 => "11011100",5602 => "11100010",5603 => "11110110",5604 => "01110010",5605 => "01111011",5606 => "01000100",5607 => "10111110",5608 => "01100001",5609 => "01001111",5610 => "01010111",5611 => "10110010",5612 => "10011001",5613 => "01110110",5614 => "01111101",5615 => "10110101",5616 => "01111100",5617 => "10111100",5618 => "00111011",5619 => "11110011",5620 => "01101101",5621 => "00101001",5622 => "00010010",5623 => "00011001",5624 => "11000011",5625 => "00110001",5626 => "10000001",5627 => "10100101",5628 => "10010000",5629 => "01000101",5630 => "00101110",5631 => "00100110",5632 => "01101011",5633 => "11000001",5634 => "01110110",5635 => "10100110",5636 => "01111101",5637 => "11001010",5638 => "00011101",5639 => "10011010",5640 => "11100001",5641 => "10000100",5642 => "00010000",5643 => "01011101",5644 => "00000000",5645 => "10000000",5646 => "10100101",5647 => "00101111",5648 => "11011001",5649 => "11101011",5650 => "10001000",5651 => "10110100",5652 => "11011001",5653 => "10011100",5654 => "00001100",5655 => "10100111",5656 => "10011001",5657 => "10110000",5658 => "00000011",5659 => "11011100",5660 => "11101111",5661 => "01000010",5662 => "11011101",5663 => "00111101",5664 => "11010011",5665 => "10011110",5666 => "10000101",5667 => "00100000",5668 => "01000101",5669 => "01000001",5670 => "10001110",5671 => "00001100",5672 => "00000110",5673 => "01010111",5674 => "01110101",5675 => "01011100",5676 => "11101011",5677 => "01011111",5678 => "11001000",5679 => "00000100",5680 => "11100000",5681 => "11100010",5682 => "01110001",5683 => "00000011",5684 => "00001110",5685 => "01101111",5686 => "01011110",5687 => "00010101",5688 => "00110101",5689 => "11100011",5690 => "10101011",5691 => "01000011",5692 => "01110010",5693 => "11111011",5694 => "11101111",5695 => "10011000",5696 => "11111101",5697 => "00111010",5698 => "00000000",5699 => "11111100",5700 => "10100111",5701 => "11001110",5702 => "11001100",5703 => "11110000",5704 => "11010001",5705 => "11100000",5706 => "10001101",5707 => "11100011",5708 => "11000111",5709 => "11011000",5710 => "00011101",5711 => "00001001",5712 => "10000111",5713 => "11100101",5714 => "10000110",5715 => "00000000",5716 => "00000011",5717 => "00101000",5718 => "11110001",5719 => "11011111",5720 => "10100010",5721 => "10111000",5722 => "10100000",5723 => "11000100",5724 => "00100101",5725 => "10011011",5726 => "11001010",5727 => "10111001",5728 => "11011101",5729 => "01000100",5730 => "01000000",5731 => "00011110",5732 => "10001110",5733 => "10001110",5734 => "01100001",5735 => "01100000",5736 => "11001000",5737 => "00000001",5738 => "10111011",5739 => "00001101",5740 => "10011111",5741 => "10001101",5742 => "01110010",5743 => "00001010",5744 => "00110100",5745 => "11111011",5746 => "11111101",5747 => "10100011",5748 => "01100111",5749 => "11101011",5750 => "00110111",5751 => "10000001",5752 => "10100101",5753 => "10000010",5754 => "01110101",5755 => "10100000",5756 => "11110011",5757 => "00101011",5758 => "11000111",5759 => "00110000",5760 => "11011000",5761 => "00101001",5762 => "11101101",5763 => "10010101",5764 => "01100010",5765 => "00101100",5766 => "01001110",5767 => "11010000",5768 => "10101011",5769 => "01001111",5770 => "01100100",5771 => "00110100",5772 => "00100100",5773 => "11010011",5774 => "01101011",5775 => "11001110",5776 => "00011100",5777 => "00111111",5778 => "10100100",5779 => "01001100",5780 => "01010001",5781 => "00111111",5782 => "00101110",5783 => "01000111",5784 => "00011100",5785 => "11011001",5786 => "10100011",5787 => "11111100",5788 => "11000101",5789 => "10001011",5790 => "10110100",5791 => "11110110",5792 => "11010101",5793 => "11101101",5794 => "00111100",5795 => "10010100",5796 => "11011010",5797 => "00100101",5798 => "00100001",5799 => "00101100",5800 => "11111100",5801 => "00111111",5802 => "00101000",5803 => "10000110",5804 => "01110110",5805 => "10100110",5806 => "11110111",5807 => "10011011",5808 => "01011110",5809 => "00010010",5810 => "10010100",5811 => "01100000",5812 => "00000010",5813 => "10111100",5814 => "10011010",5815 => "10110000",5816 => "01001001",5817 => "11111010",5818 => "01001100",5819 => "00000100",5820 => "01110101",5821 => "11000100",5822 => "11010100",5823 => "10010111",5824 => "01001010",5825 => "01110011",5826 => "00111011",5827 => "11100101",5828 => "01111000",5829 => "10011101",5830 => "01010000",5831 => "10111000",5832 => "01000000",5833 => "01110110",5834 => "01010001",5835 => "11001010",5836 => "11001111",5837 => "11011111",5838 => "01010010",5839 => "10001111",5840 => "01010001",5841 => "10111111",5842 => "00001110",5843 => "01011011",5844 => "00110001",5845 => "10111010",5846 => "10001010",5847 => "10000101",5848 => "00110000",5849 => "10100011",5850 => "11011001",5851 => "01010001",5852 => "10000000",5853 => "11111100",5854 => "10111111",5855 => "00111110",5856 => "11010001",5857 => "10101001",5858 => "10011001",5859 => "00111111",5860 => "10111001",5861 => "10101011",5862 => "00111011",5863 => "11011001",5864 => "00101101",5865 => "00101100",5866 => "10001111",5867 => "00010010",5868 => "10100101",5869 => "01110001",5870 => "01000001",5871 => "10001101",5872 => "10100011",5873 => "00011011",5874 => "00100001",5875 => "01110011",5876 => "00100001",5877 => "00000111",5878 => "11000110",5879 => "11111011",5880 => "11011000",5881 => "10101001",5882 => "11010011",5883 => "11101000",5884 => "10000100",5885 => "10000000",5886 => "00010001",5887 => "01010111",5888 => "11010100",5889 => "00100010",5890 => "01000010",5891 => "10000101",5892 => "11010111",5893 => "00001100",5894 => "00100110",5895 => "11000100",5896 => "00101110",5897 => "11100001",5898 => "11011010",5899 => "11000110",5900 => "11010111",5901 => "11001110",5902 => "00101010",5903 => "11010001",5904 => "10110011",5905 => "11000011",5906 => "00010111",5907 => "10011000",5908 => "01011000",5909 => "10111011",5910 => "01111010",5911 => "00001001",5912 => "01100110",5913 => "10001011",5914 => "01101110",5915 => "10000001",5916 => "00110100",5917 => "00010011",5918 => "01111010",5919 => "11100111",5920 => "10111000",5921 => "10000001",5922 => "00100001",5923 => "11011010",5924 => "10111011",5925 => "11000010",5926 => "01011111",5927 => "10101100",5928 => "10101111",5929 => "00001101",5930 => "00011101",5931 => "11100001",5932 => "11010101",5933 => "11001010",5934 => "11010101",5935 => "01010101",5936 => "00000011",5937 => "00010100",5938 => "11011000",5939 => "10000001",5940 => "11000110",5941 => "00010010",5942 => "00011101",5943 => "01100010",5944 => "11011010",5945 => "11000001",5946 => "11111001",5947 => "00110001",5948 => "00001001",5949 => "10001000",5950 => "10001101",5951 => "01001010",5952 => "11010011",5953 => "01011011",5954 => "10010001",5955 => "00110011",5956 => "11000010",5957 => "01011111",5958 => "00011111",5959 => "00101010",5960 => "00010101",5961 => "00110010",5962 => "00110000",5963 => "00110110",5964 => "11000111",5965 => "11011110",5966 => "01111101",5967 => "10111001",5968 => "00101100",5969 => "10110001",5970 => "00010111",5971 => "00111001",5972 => "01101000",5973 => "00001100",5974 => "10110011",5975 => "10000011",5976 => "01110011",5977 => "11010000",5978 => "00000111",5979 => "01101001",5980 => "00101010",5981 => "01110100",5982 => "00111111",5983 => "10011101",5984 => "11101111",5985 => "00100100",5986 => "10010000",5987 => "01100010",5988 => "00110011",5989 => "10011100",5990 => "11100010",5991 => "01000001",5992 => "10110010",5993 => "01001110",5994 => "10111011",5995 => "01100101",5996 => "01010111",5997 => "10011110",5998 => "00011101",5999 => "10011100",6000 => "10110011",6001 => "11011010",6002 => "00001010",6003 => "01000010",6004 => "10101010",6005 => "10000011",6006 => "00010010",6007 => "01001111",6008 => "00100010",6009 => "00100010",6010 => "01110011",6011 => "10110000",6012 => "01000010",6013 => "10001101",6014 => "01010010",6015 => "00101111",6016 => "00000110",6017 => "01111010",6018 => "00101000",6019 => "01100010",6020 => "01101100",6021 => "11100010",6022 => "00100101",6023 => "10101110",6024 => "11110001",6025 => "01101001",6026 => "01101111",6027 => "10110010",6028 => "01001100",6029 => "11100000",6030 => "11011101",6031 => "11111001",6032 => "01011011",6033 => "01110101",6034 => "00111100",6035 => "10001100",6036 => "10110011",6037 => "10011100",6038 => "11000000",6039 => "00110001",6040 => "01111110",6041 => "01110110",6042 => "01010001",6043 => "00010100",6044 => "00011001",6045 => "00010010",6046 => "00101110",6047 => "10101101",6048 => "01111101",6049 => "11101110",6050 => "00100111",6051 => "00101111",6052 => "01011100",6053 => "01010110",6054 => "10000011",6055 => "00010100",6056 => "00111110",6057 => "10010010",6058 => "11100011",6059 => "00111110",6060 => "00001110",6061 => "01011010",6062 => "00000000",6063 => "10001110",6064 => "11110110",6065 => "10101001",6066 => "10010010",6067 => "01011110",6068 => "01100011",6069 => "11100011",6070 => "11111101",6071 => "01110111",6072 => "11010100",6073 => "10111001",6074 => "01001101",6075 => "01001011",6076 => "11101000",6077 => "11100100",6078 => "01011111",6079 => "01000110",6080 => "00110110",6081 => "01111001",6082 => "10011110",6083 => "10011000",6084 => "10100001",6085 => "00000000",6086 => "10010111",6087 => "00100101",6088 => "00101111",6089 => "11101011",6090 => "01000011",6091 => "01100111",6092 => "01111010",6093 => "11000011",6094 => "00111100",6095 => "10101100",6096 => "11001100",6097 => "11111001",6098 => "00011000",6099 => "00100010",6100 => "01100100",6101 => "01101011",6102 => "01110100",6103 => "11000001",6104 => "00111000",6105 => "10111100",6106 => "10100010",6107 => "11000100",6108 => "01000110",6109 => "01001011",6110 => "00001111",6111 => "11110111",6112 => "00001110",6113 => "00111011",6114 => "11110010",6115 => "00100001",6116 => "11000011",6117 => "10101100",6118 => "01100011",6119 => "01000001",6120 => "11011111",6121 => "01000100",6122 => "10101011",6123 => "00010000",6124 => "11010001",6125 => "10101101",6126 => "01101011",6127 => "11110000",6128 => "11010100",6129 => "10010100",6130 => "01101110",6131 => "11111100",6132 => "11010000",6133 => "00101010",6134 => "01011010",6135 => "01111001",6136 => "10001100",6137 => "00110000",6138 => "11111110",6139 => "11100101",6140 => "00001000",6141 => "00101100",6142 => "01111001",6143 => "01010110",6144 => "11100101",6145 => "01101011",6146 => "10000101",6147 => "10010010",6148 => "10010100",6149 => "10101010",6150 => "11101110",6151 => "01011100",6152 => "01011100",6153 => "11101010",6154 => "10100000",6155 => "01001010",6156 => "11000000",6157 => "00010010",6158 => "01001010",6159 => "00100100",6160 => "01101101",6161 => "01110101",6162 => "00100100",6163 => "00101010",6164 => "11100100",6165 => "01011000",6166 => "00110100",6167 => "10001001",6168 => "01011001",6169 => "11010111",6170 => "11110110",6171 => "00000101",6172 => "00010111",6173 => "01110011",6174 => "00100000",6175 => "01010101",6176 => "11111010",6177 => "11101101",6178 => "01101001",6179 => "10111101",6180 => "11011111",6181 => "01010011",6182 => "00000000",6183 => "10101110",6184 => "10101101",6185 => "11110010",6186 => "11100111",6187 => "01111100",6188 => "01010001",6189 => "11001000",6190 => "01101010",6191 => "01100100",6192 => "01101110",6193 => "11000000",6194 => "01110001",6195 => "01011111",6196 => "10000001",6197 => "10100001",6198 => "11101000",6199 => "11010011",6200 => "11111000",6201 => "01011110",6202 => "11001011",6203 => "10001011",6204 => "00111000",6205 => "01111011",6206 => "10101011",6207 => "00000100",6208 => "00111010",6209 => "10101100",6210 => "01010010",6211 => "11001011",6212 => "11100011",6213 => "01101000",6214 => "01001101",6215 => "00101001",6216 => "11001111",6217 => "00101110",6218 => "00000100",6219 => "01111000",6220 => "01101011",6221 => "10110010",6222 => "10110011",6223 => "11110000",6224 => "00011101",6225 => "10110010",6226 => "11011101",6227 => "00111011",6228 => "01111001",6229 => "01101001",6230 => "00001101",6231 => "00000001",6232 => "10011101",6233 => "11101101",6234 => "01001111",6235 => "00101011",6236 => "01011001",6237 => "11011101",6238 => "00000101",6239 => "00111110",6240 => "11010100",6241 => "00111010",6242 => "01010110",6243 => "01010101",6244 => "01100000",6245 => "01000101",6246 => "10110001",6247 => "10010101",6248 => "10110010",6249 => "00001100",6250 => "10100111",6251 => "11111010",6252 => "00010011",6253 => "01110001",6254 => "11000011",6255 => "11111010",6256 => "00001011",6257 => "01111100",6258 => "11001011",6259 => "11000110",6260 => "10000101",6261 => "11101110",6262 => "10110011",6263 => "01110110",6264 => "11101100",6265 => "01110000",6266 => "00011011",6267 => "11111101",6268 => "10110011",6269 => "00010011",6270 => "00100011",6271 => "10001010",6272 => "11101101",6273 => "00100100",6274 => "01000001",6275 => "11001010",6276 => "01110100",6277 => "01101111",6278 => "11000000",6279 => "00000111",6280 => "11010111",6281 => "00110110",6282 => "10110100",6283 => "10100010",6284 => "01100011",6285 => "10000110",6286 => "01110101",6287 => "01111011",6288 => "11001101",6289 => "11111011",6290 => "01001010",6291 => "11111111",6292 => "00011110",6293 => "01011011",6294 => "00011001",6295 => "11110011",6296 => "11100110",6297 => "11110100",6298 => "00110001",6299 => "11111100",6300 => "00101000",6301 => "11010110",6302 => "01110001",6303 => "11101001",6304 => "00110011",6305 => "11010111",6306 => "00010000",6307 => "00011000",6308 => "11011110",6309 => "00010010",6310 => "10110011",6311 => "01010000",6312 => "11101111",6313 => "10110110",6314 => "01100001",6315 => "00010000",6316 => "01100100",6317 => "11001111",6318 => "00101011",6319 => "00000011",6320 => "11110111",6321 => "11100010",6322 => "10000101",6323 => "00001110",6324 => "01001001",6325 => "01111101",6326 => "10101000",6327 => "11100011",6328 => "01111011",6329 => "01101001",6330 => "10100000",6331 => "11111101",6332 => "00101101",6333 => "11101010",6334 => "00010010",6335 => "01000110",6336 => "10110010",6337 => "10100110",6338 => "10101100",6339 => "10000010",6340 => "11110100",6341 => "10110100",6342 => "10010001",6343 => "00011000",6344 => "11010110",6345 => "00110011",6346 => "11100101",6347 => "10100001",6348 => "11010011",6349 => "01001000",6350 => "11100100",6351 => "11000111",6352 => "11001011",6353 => "11000101",6354 => "11001001",6355 => "10010011",6356 => "01101110",6357 => "10000011",6358 => "01110010",6359 => "00111111",6360 => "01001011",6361 => "11010110",6362 => "11010110",6363 => "00100010",6364 => "01000010",6365 => "10001101",6366 => "11111100",6367 => "10110111",6368 => "11001100",6369 => "10100100",6370 => "01000000",6371 => "10100110",6372 => "10101101",6373 => "11110110",6374 => "11000000",6375 => "10000110",6376 => "01011110",6377 => "01001000",6378 => "10100110",6379 => "00101101",6380 => "01101111",6381 => "10010010",6382 => "10000111",6383 => "01011111",6384 => "11100010",6385 => "10011010",6386 => "00101110",6387 => "10111100",6388 => "00111001",6389 => "11101101",6390 => "00010000",6391 => "00001010",6392 => "00001011",6393 => "11000011",6394 => "01101000",6395 => "11110000",6396 => "00100101",6397 => "11011001",6398 => "11101000",6399 => "01110111",6400 => "10110110",6401 => "00100110",6402 => "01100111",6403 => "01011001",6404 => "00110001",6405 => "00011010",6406 => "11001000",6407 => "00110100",6408 => "11100111",6409 => "11000111",6410 => "11100101",6411 => "00010110",6412 => "10100101",6413 => "11010101",6414 => "11110101",6415 => "11101110",6416 => "01111011",6417 => "01110010",6418 => "00001110",6419 => "01110001",6420 => "11100010",6421 => "11011100",6422 => "11111101",6423 => "11000001",6424 => "00000111",6425 => "10100011",6426 => "01000001",6427 => "01010100",6428 => "10000101",6429 => "11110101",6430 => "11011001",6431 => "01001000",6432 => "00000000",6433 => "00010111",6434 => "11011001",6435 => "10111010",6436 => "10000001",6437 => "11011101",6438 => "00111110",6439 => "10100111",6440 => "00110001",6441 => "01101010",6442 => "01000111",6443 => "00011011",6444 => "11100000",6445 => "10010010",6446 => "00011101",6447 => "10001110",6448 => "01110110",6449 => "11100001",6450 => "01001111",6451 => "10010110",6452 => "11001101",6453 => "00010100",6454 => "00110101",6455 => "01110101",6456 => "11000110",6457 => "00110010",6458 => "10100101",6459 => "10010100",6460 => "01010111",6461 => "11010111",6462 => "01000101",6463 => "01111001",6464 => "01000000",6465 => "10011110",6466 => "11111011",6467 => "01011100",6468 => "00111000",6469 => "00101001",6470 => "01111101",6471 => "01101000",6472 => "00101110",6473 => "10010011",6474 => "10100101",6475 => "01101110",6476 => "00110001",6477 => "11011101",6478 => "10101111",6479 => "01100010",6480 => "00000011",6481 => "11101101",6482 => "11110010",6483 => "00000000",6484 => "01010010",6485 => "00100111",6486 => "11011101",6487 => "11010000",6488 => "01001111",6489 => "01111001",6490 => "00110110",6491 => "00000001",6492 => "00110001",6493 => "10001000",6494 => "11011000",6495 => "10111100",6496 => "11010011",6497 => "01110011",6498 => "10001010",6499 => "00100001",6500 => "10100111",6501 => "00010011",6502 => "10011110",6503 => "11011101",6504 => "11000111",6505 => "01000110",6506 => "10010111",6507 => "00111011",6508 => "11111011",6509 => "00100010",6510 => "10101100",6511 => "01000110",6512 => "11001111",6513 => "01100011",6514 => "00001111",6515 => "10110111",6516 => "10001100",6517 => "00111100",6518 => "10100000",6519 => "01101010",6520 => "00000001",6521 => "00010110",6522 => "01111100",6523 => "10111111",6524 => "00111101",6525 => "10010101",6526 => "10101101",6527 => "00111001",6528 => "11110111",6529 => "01101010",6530 => "11000011",6531 => "00101011",6532 => "01000001",6533 => "11010011",6534 => "01100101",6535 => "00100010",6536 => "11100001",6537 => "01101100",6538 => "10100010",6539 => "10000110",6540 => "01110111",6541 => "10000010",6542 => "01100000",6543 => "01001010",6544 => "10010010",6545 => "10001010",6546 => "11110001",6547 => "11110110",6548 => "11000001",6549 => "00001010",6550 => "00101000",6551 => "11111000",6552 => "01001000",6553 => "00000000",6554 => "11100101",6555 => "10010111",6556 => "11101110",6557 => "11001100",6558 => "00110110",6559 => "10010111",6560 => "10101110",6561 => "11111011",6562 => "11000100",6563 => "10000001",6564 => "00111111",6565 => "11111111",6566 => "10101110",6567 => "01110011",6568 => "11110000",6569 => "01011110",6570 => "11100101",6571 => "11111011",6572 => "10000111",6573 => "11111000",6574 => "11010111",6575 => "11001101",6576 => "10000000",6577 => "10110110",6578 => "10011010",6579 => "01010111",6580 => "00010110",6581 => "00000111",6582 => "10111010",6583 => "00110101",6584 => "00000000",6585 => "01001111",6586 => "01111010",6587 => "01001100",6588 => "00101100",6589 => "00110101",6590 => "11111111",6591 => "00000001",6592 => "10100000",6593 => "01011011",6594 => "00100101",6595 => "11110011",6596 => "11101000",6597 => "00011001",6598 => "01001100",6599 => "01000010",6600 => "11101100",6601 => "01001100",6602 => "00111010",6603 => "00011001",6604 => "10010001",6605 => "11000110",6606 => "01100010",6607 => "10110111",6608 => "01001000",6609 => "10110001",6610 => "01111111",6611 => "00100100",6612 => "01110110",6613 => "00010000",6614 => "10010010",6615 => "01011000",6616 => "10101000",6617 => "10101010",6618 => "00110010",6619 => "11101110",6620 => "01111001",6621 => "10101000",6622 => "01101010",6623 => "00010001",6624 => "01010000",6625 => "11011000",6626 => "10110001",6627 => "00000001",6628 => "11101100",6629 => "11110101",6630 => "00010111",6631 => "01101001",6632 => "11100100",6633 => "10101111",6634 => "11101101",6635 => "01100011",6636 => "01111010",6637 => "01010101",6638 => "11110101",6639 => "01100010",6640 => "11110001",6641 => "00111001",6642 => "01100000",6643 => "11001000",6644 => "10001101",6645 => "01100001",6646 => "10000010",6647 => "01001001",6648 => "10010110",6649 => "10001101",6650 => "11101010",6651 => "11100000",6652 => "10000101",6653 => "10011010",6654 => "01001011",6655 => "11100000",6656 => "01010010",6657 => "00011111",6658 => "01111011",6659 => "00110001",6660 => "00000000",6661 => "00111100",6662 => "11000011",6663 => "00110101",6664 => "11111100",6665 => "00000111",6666 => "10001010",6667 => "01111011",6668 => "10111101",6669 => "01110100",6670 => "01001111",6671 => "01100001",6672 => "10111011",6673 => "10000100",6674 => "01110110",6675 => "01111101",6676 => "00100010",6677 => "01010101",6678 => "01111011",6679 => "10010100",6680 => "11001001",6681 => "10101111",6682 => "00110111",6683 => "11000001",6684 => "11011110",6685 => "10101110",6686 => "00001010",6687 => "00011100",6688 => "01011010",6689 => "00000011",6690 => "00000010",6691 => "01111100",6692 => "10101011",6693 => "11010110",6694 => "00111000",6695 => "10110011",6696 => "11010110",6697 => "11001110",6698 => "10100101",6699 => "10110010",6700 => "01101100",6701 => "00111111",6702 => "11001010",6703 => "01101110",6704 => "01100010",6705 => "11101001",6706 => "01000101",6707 => "11010110",6708 => "01000110",6709 => "10110001",6710 => "01101110",6711 => "01000011",6712 => "00000001",6713 => "10000011",6714 => "00101001",6715 => "11001101",6716 => "01100100",6717 => "11110100",6718 => "00000001",6719 => "00111000",6720 => "01111001",6721 => "11001111",6722 => "00100101",6723 => "10101101",6724 => "01001110",6725 => "10011000",6726 => "01111001",6727 => "00110000",6728 => "00101101",6729 => "11010100",6730 => "01010111",6731 => "01011011",6732 => "11000101",6733 => "11001000",6734 => "10110011",6735 => "01010011",6736 => "10111101",6737 => "10001100",6738 => "00000100",6739 => "11010000",6740 => "10000100",6741 => "10001111",6742 => "11000000",6743 => "11010011",6744 => "10010010",6745 => "11101110",6746 => "01100110",6747 => "00010100",6748 => "10100111",6749 => "00010100",6750 => "01110001",6751 => "01011010",6752 => "00101101",6753 => "01000001",6754 => "10100100",6755 => "00110010",6756 => "01001011",6757 => "10111101",6758 => "10110101",6759 => "10110101",6760 => "11101011",6761 => "10111100",6762 => "00101101",6763 => "01010001",6764 => "10011100",6765 => "10000110",6766 => "10111011",6767 => "11001001",6768 => "01011000",6769 => "10100000",6770 => "10010000",6771 => "01001101",6772 => "10001110",6773 => "00101101",6774 => "10111000",6775 => "00100000",6776 => "01111111",6777 => "00010000",6778 => "10100101",6779 => "00010000",6780 => "00001100",6781 => "10001010",6782 => "00111000",6783 => "10100001",6784 => "00010101",6785 => "11101111",6786 => "00011111",6787 => "00100000",6788 => "01001100",6789 => "00111000",6790 => "01001111",6791 => "00000001",6792 => "00110101",6793 => "11101011",6794 => "10111010",6795 => "00100101",6796 => "11010000",6797 => "01011011",6798 => "11001100",6799 => "11001000",6800 => "01011010",6801 => "10111011",6802 => "10011000",6803 => "11011001",6804 => "00100010",6805 => "10110111",6806 => "10111111",6807 => "01011011",6808 => "01110110",6809 => "00011101",6810 => "10011111",6811 => "11101110",6812 => "01100100",6813 => "01110011",6814 => "00001010",6815 => "10011101",6816 => "11100110",6817 => "10010101",6818 => "01010001",6819 => "01110000",6820 => "10011101",6821 => "10000010",6822 => "10101011",6823 => "11000011",6824 => "01100110",6825 => "00000100",6826 => "11010110",6827 => "01001111",6828 => "10110010",6829 => "01100010",6830 => "10001000",6831 => "11100100",6832 => "01100000",6833 => "11010100",6834 => "11110101",6835 => "01110010",6836 => "10111100",6837 => "10101000",6838 => "11000010",6839 => "01001110",6840 => "00101000",6841 => "11001111",6842 => "11001111",6843 => "01111110",6844 => "11100001",6845 => "01101101",6846 => "11100011",6847 => "00011101",6848 => "00100110",6849 => "01001000",6850 => "11011000",6851 => "10000010",6852 => "11100011",6853 => "01010100",6854 => "00111101",6855 => "01110101",6856 => "00010111",6857 => "10110110",6858 => "10001001",6859 => "10111101",6860 => "00110110",6861 => "01111100",6862 => "01100101",6863 => "01110011",6864 => "00010101",6865 => "11110111",6866 => "11011000",6867 => "01111000",6868 => "10000100",6869 => "11000101",6870 => "11010101",6871 => "11011001",6872 => "01110001",6873 => "11011100",6874 => "01010000",6875 => "01000000",6876 => "10000000",6877 => "10000000",6878 => "11101000",6879 => "00001100",6880 => "01110010",6881 => "01111100",6882 => "01101100",6883 => "00111011",6884 => "10000010",6885 => "10101010",6886 => "10111111",6887 => "10011010",6888 => "01011110",6889 => "11001010",6890 => "00011101",6891 => "10011100",6892 => "00110000",6893 => "11110000",6894 => "01110010",6895 => "01111110",6896 => "10100011",6897 => "11111001",6898 => "01100000",6899 => "01111001",6900 => "10011000",6901 => "11100101",6902 => "01100000",6903 => "10100111",6904 => "11111100",6905 => "11000010",6906 => "10101100",6907 => "10011010",6908 => "01110011",6909 => "00010010",6910 => "10010010",6911 => "00111011",6912 => "10011010",6913 => "10000001",6914 => "00000001",6915 => "10000010",6916 => "01000000",6917 => "11011111",6918 => "01110010",6919 => "11011100",6920 => "11000000",6921 => "01110100",6922 => "00101000",6923 => "11101011",6924 => "11010111",6925 => "11111011",6926 => "00000010",6927 => "11001010",6928 => "11100111",6929 => "00001000",6930 => "10010101",6931 => "00100110",6932 => "11110101",6933 => "11010000",6934 => "11100100",6935 => "00110001",6936 => "01100000",6937 => "01101111",6938 => "11000110",6939 => "01101110",6940 => "10001001",6941 => "10010010",6942 => "00001001",6943 => "10011110",6944 => "00100001",6945 => "00111000",6946 => "01111011",6947 => "00101000",6948 => "01001101",6949 => "01001010",6950 => "00010111",6951 => "10111011",6952 => "10111011",6953 => "00010111",6954 => "00000100",6955 => "10110110",6956 => "01011001",6957 => "10110001",6958 => "11100100",6959 => "10000000",6960 => "10111001",6961 => "11101010",6962 => "11100011",6963 => "01001100",6964 => "10110111",6965 => "11001000",6966 => "00011001",6967 => "00010010",6968 => "10011110",6969 => "01010110",6970 => "11000010",6971 => "00100101",6972 => "11010011",6973 => "01101010",6974 => "00101010",6975 => "00001100",6976 => "10101011",6977 => "10001101",6978 => "01001100",6979 => "00000101",6980 => "00101010",6981 => "01011110",6982 => "11100001",6983 => "10010010",6984 => "01111000",6985 => "01100101",6986 => "11010001",6987 => "10110010",6988 => "11111100",6989 => "00001010",6990 => "01010111",6991 => "10000111",6992 => "00010101",6993 => "01001000",6994 => "01000100",6995 => "10010111",6996 => "01000101",6997 => "00000101",6998 => "01110101",6999 => "10110100",7000 => "11101011",7001 => "00100001",7002 => "11100011",7003 => "00100001",7004 => "10000110",7005 => "11110000",7006 => "01110111",7007 => "11111001",7008 => "00110010",7009 => "10010110",7010 => "01110110",7011 => "11001001",7012 => "11111110",7013 => "11111101",7014 => "00111100",7015 => "01110001",7016 => "01001011",7017 => "10100011",7018 => "11010011",7019 => "01000011",7020 => "11100101",7021 => "00110101",7022 => "10101110",7023 => "11010111",7024 => "01101000",7025 => "11101011",7026 => "10001010",7027 => "10010011",7028 => "10101101",7029 => "00111011",7030 => "11101011",7031 => "00101010",7032 => "00101011",7033 => "00000111",7034 => "01111010",7035 => "00101001",7036 => "01011111",7037 => "01000100",7038 => "10011110",7039 => "00001011",7040 => "11001010",7041 => "00010101",7042 => "11010001",7043 => "11111000",7044 => "11101000",7045 => "01111000",7046 => "10100011",7047 => "10100110",7048 => "11001100",7049 => "01101101",7050 => "11101110",7051 => "01011000",7052 => "11011001",7053 => "00000010",7054 => "10111010",7055 => "00111010",7056 => "01010101",7057 => "11011101",7058 => "11110010",7059 => "00110010",7060 => "00100110",7061 => "01011100",7062 => "01101110",7063 => "01110011",7064 => "11111110",7065 => "01111111",7066 => "10111110",7067 => "10000100",7068 => "11100001",7069 => "11011000",7070 => "11001011",7071 => "10010011",7072 => "11111110",7073 => "00110110",7074 => "11011101",7075 => "00001011",7076 => "10101101",7077 => "00110010",7078 => "11110010",7079 => "10101011",7080 => "10000000",7081 => "01101011",7082 => "10110111",7083 => "10011001",7084 => "11010011",7085 => "10000001",7086 => "01100011",7087 => "11110101",7088 => "10110010",7089 => "01101001",7090 => "01011010",7091 => "10001010",7092 => "11011011",7093 => "01000011",7094 => "10100111",7095 => "10010111",7096 => "10010100",7097 => "00101100",7098 => "00010100",7099 => "10110110",7100 => "11101000",7101 => "11100110",7102 => "00100101",7103 => "00110101",7104 => "11011011",7105 => "01000001",7106 => "01100000",7107 => "10111101",7108 => "00011110",7109 => "01000100",7110 => "11111100",7111 => "01110111",7112 => "01101111",7113 => "10111011",7114 => "10010010",7115 => "10001010",7116 => "00011101",7117 => "00100110",7118 => "11001010",7119 => "10111011",7120 => "11010100",7121 => "11010101",7122 => "01110111",7123 => "11010101",7124 => "11000000",7125 => "00000100",7126 => "10100100",7127 => "11010010",7128 => "11110000",7129 => "11001110",7130 => "11001011",7131 => "11001011",7132 => "01111010",7133 => "01110010",7134 => "00111001",7135 => "00001101",7136 => "01100000",7137 => "10001101",7138 => "01101010",7139 => "01001111",7140 => "11110000",7141 => "10101111",7142 => "01001101",7143 => "00111010",7144 => "00100101",7145 => "11111110",7146 => "11111011",7147 => "00010001",7148 => "01110111",7149 => "10101010",7150 => "01111010",7151 => "10010001",7152 => "11110001",7153 => "11000110",7154 => "00000001",7155 => "11000101",7156 => "11010111",7157 => "01100101",7158 => "11001101",7159 => "10011010",7160 => "10000100",7161 => "00110100",7162 => "10101110",7163 => "10111000",7164 => "10100101",7165 => "11101000",7166 => "10110110",7167 => "01010001",7168 => "00001110",7169 => "11100100",7170 => "11001010",7171 => "00111010",7172 => "01110011",7173 => "10001101",7174 => "11101110",7175 => "11001111",7176 => "11100111",7177 => "00111010",7178 => "00110010",7179 => "00000000",7180 => "10001111",7181 => "10011001",7182 => "01111010",7183 => "01000110",7184 => "11010010",7185 => "00111011",7186 => "11101101",7187 => "11000111",7188 => "00111101",7189 => "00101000",7190 => "11111111",7191 => "10101011",7192 => "11001001",7193 => "10100111",7194 => "00001110",7195 => "00101011",7196 => "10001101",7197 => "00110100",7198 => "01010111",7199 => "01001011",7200 => "10011110",7201 => "10000011",7202 => "11011001",7203 => "00110101",7204 => "01111100",7205 => "10110001",7206 => "01111101",7207 => "10111001",7208 => "00110000",7209 => "10011101",7210 => "10000100",7211 => "11100011",7212 => "10111010",7213 => "10100101",7214 => "11111100",7215 => "11010010",7216 => "10110100",7217 => "01001101",7218 => "01100101",7219 => "00010001",7220 => "11001010",7221 => "01111001",7222 => "10001111",7223 => "00001111",7224 => "01100111",7225 => "01000000",7226 => "11000110",7227 => "11011000",7228 => "11111011",7229 => "11100110",7230 => "10101111",7231 => "01011010",7232 => "01110110",7233 => "11110010",7234 => "11000100",7235 => "10101101",7236 => "00000111",7237 => "00100100",7238 => "00110100",7239 => "00100001",7240 => "10100000",7241 => "01110010",7242 => "10110011",7243 => "11000100",7244 => "01001001",7245 => "10011110",7246 => "00101100",7247 => "11000011",7248 => "10110010",7249 => "00110011",7250 => "00010100",7251 => "10111001",7252 => "11000011",7253 => "11110101",7254 => "00100000",7255 => "01100010",7256 => "01100001",7257 => "00011111",7258 => "11001111",7259 => "00111001",7260 => "11001011",7261 => "10101000",7262 => "00011111",7263 => "01000001",7264 => "11100000",7265 => "00011101",7266 => "00111010",7267 => "01011010",7268 => "10110111",7269 => "01110011",7270 => "10100011",7271 => "00101001",7272 => "00111001",7273 => "11001100",7274 => "11010001",7275 => "01000001",7276 => "10110111",7277 => "01111110",7278 => "10101000",7279 => "00111110",7280 => "00101111",7281 => "00110001",7282 => "11010010",7283 => "00100011",7284 => "11000100",7285 => "00001001",7286 => "11010010",7287 => "00001101",7288 => "11010001",7289 => "01101111",7290 => "10000001",7291 => "01111011",7292 => "01010100",7293 => "01101010",7294 => "10110111",7295 => "00011011",7296 => "01101101",7297 => "11100101",7298 => "10100010",7299 => "11111000",7300 => "01000101",7301 => "00010111",7302 => "01010010",7303 => "11100111",7304 => "00001011",7305 => "00101100",7306 => "11001111",7307 => "01101011",7308 => "00111100",7309 => "00100010",7310 => "00011000",7311 => "10011111",7312 => "01100111",7313 => "10011111",7314 => "00010011",7315 => "10100101",7316 => "01000110",7317 => "01111101",7318 => "10111100",7319 => "01001000",7320 => "11011100",7321 => "11010010",7322 => "10111111",7323 => "10011001",7324 => "10011100",7325 => "10101001",7326 => "00000000",7327 => "00001100",7328 => "10100011",7329 => "10000100",7330 => "11000100",7331 => "01111100",7332 => "10110101",7333 => "01001101",7334 => "00000000",7335 => "10001100",7336 => "00001101",7337 => "11000001",7338 => "10010000",7339 => "01011110",7340 => "10111010",7341 => "00100010",7342 => "01001000",7343 => "01101111",7344 => "10000010",7345 => "11011001",7346 => "01110011",7347 => "00101101",7348 => "01100111",7349 => "00101111",7350 => "11000000",7351 => "10110100",7352 => "11110010",7353 => "00101011",7354 => "01101100",7355 => "10000110",7356 => "11000011",7357 => "11110101",7358 => "11101011",7359 => "11100011",7360 => "10001001",7361 => "11101001",7362 => "00010011",7363 => "10100110",7364 => "10000110",7365 => "01000101",7366 => "10111111",7367 => "00011011",7368 => "00101111",7369 => "00000111",7370 => "11000001",7371 => "01000110",7372 => "10000111",7373 => "01000101",7374 => "00100011",7375 => "01111110",7376 => "00010100",7377 => "00101101",7378 => "10101110",7379 => "00100100",7380 => "00110110",7381 => "00101101",7382 => "01101000",7383 => "00000000",7384 => "01001111",7385 => "01011001",7386 => "00100110",7387 => "00101101",7388 => "10001111",7389 => "01110010",7390 => "10101010",7391 => "01100100",7392 => "01111101",7393 => "00100000",7394 => "00101001",7395 => "00100001",7396 => "01110000",7397 => "10000000",7398 => "01010110",7399 => "00001100",7400 => "11001111",7401 => "11000100",7402 => "00001111",7403 => "01101000",7404 => "01011000",7405 => "01111101",7406 => "01010010",7407 => "01010101",7408 => "00101010",7409 => "11101011",7410 => "10011101",7411 => "11111110",7412 => "01110111",7413 => "00011110",7414 => "01110111",7415 => "10101110",7416 => "11100101",7417 => "10010101",7418 => "01001111",7419 => "01001001",7420 => "10101111",7421 => "11000011",7422 => "10000001",7423 => "11000110",7424 => "01001001",7425 => "01010111",7426 => "10010001",7427 => "01000100",7428 => "11011110",7429 => "10000010",7430 => "01101010",7431 => "01000010",7432 => "00001010",7433 => "00110011",7434 => "00000000",7435 => "01100001",7436 => "10011010",7437 => "10111111",7438 => "00000111",7439 => "10110111",7440 => "11111000",7441 => "11111001",7442 => "10010100",7443 => "10000011",7444 => "01000001",7445 => "00111011",7446 => "11110110",7447 => "01101001",7448 => "11100100",7449 => "01100111",7450 => "10101011",7451 => "11001110",7452 => "10010101",7453 => "11111101",7454 => "10101100",7455 => "00111110",7456 => "00100111",7457 => "00001101",7458 => "01111111",7459 => "11100101",7460 => "10011110",7461 => "11111110",7462 => "01111010",7463 => "10110101",7464 => "11111110",7465 => "01001000",7466 => "10101111",7467 => "00100000",7468 => "10111100",7469 => "10100011",7470 => "11111101",7471 => "11101001",7472 => "00001000",7473 => "00001101",7474 => "11110010",7475 => "10100010",7476 => "01110111",7477 => "01101011",7478 => "10110000",7479 => "11010001",7480 => "00011111",7481 => "00111000",7482 => "00110000",7483 => "10011000",7484 => "00011011",7485 => "01100100",7486 => "00001110",7487 => "00111110",7488 => "11000100",7489 => "10001000",7490 => "10100001",7491 => "11101011",7492 => "11100010",7493 => "01000001",7494 => "10111000",7495 => "10100110",7496 => "01001100",7497 => "11111001",7498 => "10010101",7499 => "10100110",7500 => "01110011",7501 => "10011011",7502 => "11010111",7503 => "10001101",7504 => "00010110",7505 => "01010010",7506 => "11101111",7507 => "10011001",7508 => "00100111",7509 => "00011000",7510 => "00111011",7511 => "00000100",7512 => "01001101",7513 => "11011000",7514 => "10101001",7515 => "00111011",7516 => "11111101",7517 => "00000010",7518 => "10111000",7519 => "11010001",7520 => "10001101",7521 => "00101111",7522 => "10010000",7523 => "01011100",7524 => "01001000",7525 => "10100100",7526 => "10011001",7527 => "10110100",7528 => "01011010",7529 => "11111101",7530 => "00011010",7531 => "11100110",7532 => "11101100",7533 => "11001100",7534 => "00000100",7535 => "10100011",7536 => "11000101",7537 => "01000001",7538 => "11010100",7539 => "01111100",7540 => "00011000",7541 => "01111101",7542 => "01000000",7543 => "11100110",7544 => "00000010",7545 => "01000001",7546 => "00101110",7547 => "01011011",7548 => "11000010",7549 => "00010000",7550 => "10010001",7551 => "01110110",7552 => "11101010",7553 => "00101001",7554 => "10010010",7555 => "01110110",7556 => "01110001",7557 => "10110001",7558 => "11110100",7559 => "01110101",7560 => "10010110",7561 => "11000101",7562 => "00101110",7563 => "00111100",7564 => "11111011",7565 => "10111111",7566 => "11100001",7567 => "10001111",7568 => "10101000",7569 => "11110000",7570 => "11100100",7571 => "00110010",7572 => "01001011",7573 => "01000000",7574 => "10111111",7575 => "11000001",7576 => "11000000",7577 => "11010000",7578 => "00011010",7579 => "11000011",7580 => "00001001",7581 => "10101010",7582 => "01011001",7583 => "11110000",7584 => "10010111",7585 => "11010101",7586 => "10000101",7587 => "01000100",7588 => "10101111",7589 => "10110011",7590 => "00011110",7591 => "10100010",7592 => "00111011",7593 => "10001001",7594 => "00000010",7595 => "11000000",7596 => "00001001",7597 => "11010001",7598 => "01000111",7599 => "01011101",7600 => "10000111",7601 => "01101100",7602 => "10100101",7603 => "11000011",7604 => "01011101",7605 => "11001001",7606 => "00011011",7607 => "10000001",7608 => "00101101",7609 => "01010110",7610 => "10111010",7611 => "11001010",7612 => "01011110",7613 => "01110011",7614 => "01010011",7615 => "01110111",7616 => "00001001",7617 => "10000100",7618 => "10100101",7619 => "00000111",7620 => "01110011",7621 => "01111010",7622 => "10011100",7623 => "01000011",7624 => "00011010",7625 => "01111011",7626 => "10100111",7627 => "11111110",7628 => "00100110",7629 => "11011100",7630 => "00100111",7631 => "01110100",7632 => "00000111",7633 => "01101011",7634 => "11100110",7635 => "11111001",7636 => "00100100",7637 => "10100011",7638 => "10000100",7639 => "00100010",7640 => "11110000",7641 => "00100010",7642 => "10110011",7643 => "10111100",7644 => "00101010",7645 => "11010110",7646 => "00111110",7647 => "11000001",7648 => "01010111",7649 => "11110011",7650 => "10100111",7651 => "01001101",7652 => "00000011",7653 => "11101001",7654 => "01011010",7655 => "10010001",7656 => "01001110",7657 => "01110101",7658 => "01010101",7659 => "00000000",7660 => "00000000",7661 => "00101000",7662 => "10000011",7663 => "11000000",7664 => "11111011",7665 => "10010010",7666 => "00100001",7667 => "11001000",7668 => "10110101",7669 => "11001100",7670 => "01010010",7671 => "10100001",7672 => "01111011",7673 => "00001001",7674 => "10101001",7675 => "10101100",7676 => "11001101",7677 => "10011011",7678 => "10100000",7679 => "00111010",7680 => "01100110",7681 => "01011100",7682 => "10100111",7683 => "00000011",7684 => "01100111",7685 => "00110010",7686 => "10110111",7687 => "11011000",7688 => "11111011",7689 => "00100011",7690 => "00001100",7691 => "00001111",7692 => "01100101",7693 => "10100110",7694 => "00001011",7695 => "10001000",7696 => "01101000",7697 => "11011110",7698 => "00111100",7699 => "10010000",7700 => "11010111",7701 => "01110000",7702 => "11000000",7703 => "00111010",7704 => "11010011",7705 => "01001110",7706 => "10100110",7707 => "01101111",7708 => "11101101",7709 => "10000101",7710 => "11100111",7711 => "10100000",7712 => "01001110",7713 => "00011000",7714 => "00111110",7715 => "11001011",7716 => "00110001",7717 => "01011001",7718 => "01110011",7719 => "01000100",7720 => "10111100",7721 => "10100010",7722 => "11111101",7723 => "00011110",7724 => "11011000",7725 => "10011010",7726 => "01011110",7727 => "01100100",7728 => "01111111",7729 => "01100000",7730 => "10011001",7731 => "00011101",7732 => "10101010",7733 => "11111110",7734 => "11001110",7735 => "00100101",7736 => "00010111",7737 => "01110110",7738 => "10101011",7739 => "00110011",7740 => "11111011",7741 => "10111010",7742 => "11011101",7743 => "10111000",7744 => "00000100",7745 => "00111101",7746 => "01110101",7747 => "00011100",7748 => "00111011",7749 => "01110110",7750 => "10010110",7751 => "00101010",7752 => "01111010",7753 => "11100101",7754 => "00110011",7755 => "11011100",7756 => "01100111",7757 => "10101000",7758 => "01100000",7759 => "00000111",7760 => "00101000",7761 => "00110110",7762 => "00000011",7763 => "00110011",7764 => "00100000",7765 => "11000010",7766 => "11010010",7767 => "00000110",7768 => "01001110",7769 => "00000011",7770 => "00101010",7771 => "10101011",7772 => "01100011",7773 => "01011101",7774 => "11010100",7775 => "11011001",7776 => "10000000",7777 => "11011110",7778 => "11110011",7779 => "00100001",7780 => "10110001",7781 => "01010101",7782 => "01011011",7783 => "00001100",7784 => "10011100",7785 => "01000010",7786 => "11001001",7787 => "01011000",7788 => "00111110",7789 => "00101111",7790 => "10111010",7791 => "11011110",7792 => "01111111",7793 => "01000001",7794 => "00011100",7795 => "10011110",7796 => "10111001",7797 => "00010000",7798 => "01101100",7799 => "01101101",7800 => "00010010",7801 => "00000000",7802 => "00010001",7803 => "01001001",7804 => "11101010",7805 => "11101001",7806 => "01010111",7807 => "01110110",7808 => "01011011",7809 => "10101110",7810 => "00110110",7811 => "10011101",7812 => "00000110",7813 => "11011010",7814 => "10000011",7815 => "11011111",7816 => "00001101",7817 => "01011100",7818 => "00110111",7819 => "01101101",7820 => "10001010",7821 => "01010010",7822 => "10010001",7823 => "01010111",7824 => "01101100",7825 => "01110000",7826 => "01011100",7827 => "00101011",7828 => "10000011",7829 => "10000010",7830 => "00000011",7831 => "01010100",7832 => "10110001",7833 => "10000110",7834 => "10100101",7835 => "10010111",7836 => "11010101",7837 => "10111001",7838 => "10001010",7839 => "00111000",7840 => "01000100",7841 => "10111101",7842 => "11011011",7843 => "00000101",7844 => "00000011",7845 => "11111010",7846 => "00101010",7847 => "10001111",7848 => "11100000",7849 => "10011111",7850 => "00000000",7851 => "01001010",7852 => "01011000",7853 => "00100010",7854 => "11110001",7855 => "11001111",7856 => "01010011",7857 => "10011011",7858 => "00010101",7859 => "11111110",7860 => "00100000",7861 => "00011011",7862 => "01101110",7863 => "01100100",7864 => "11101000",7865 => "01001100",7866 => "00111111",7867 => "00000000",7868 => "01000010",7869 => "11001010",7870 => "00110101",7871 => "11101110",7872 => "10001010",7873 => "11101111",7874 => "11010111",7875 => "11101111",7876 => "00100000",7877 => "10000010",7878 => "00100000",7879 => "00110000",7880 => "10011011",7881 => "10010111",7882 => "01111110",7883 => "10011011",7884 => "01001000",7885 => "01101110",7886 => "01100001",7887 => "10000010",7888 => "00010101",7889 => "00100010",7890 => "01011111",7891 => "10100100",7892 => "00011011",7893 => "10110100",7894 => "10110101",7895 => "10111100",7896 => "01100000",7897 => "01001001",7898 => "00100100",7899 => "10011110",7900 => "00001101",7901 => "00011100",7902 => "11001000",7903 => "01111000",7904 => "00111000",7905 => "10110011",7906 => "11100101",7907 => "10101101",7908 => "10000111",7909 => "00111111",7910 => "00001001",7911 => "11010111",7912 => "00100000",7913 => "11000101",7914 => "10000010",7915 => "00101111",7916 => "11011111",7917 => "01100101",7918 => "00101001",7919 => "00100101",7920 => "11110011",7921 => "00010110",7922 => "10011111",7923 => "10011111",7924 => "11100100",7925 => "00110101",7926 => "00000010",7927 => "10110000",7928 => "01010100",7929 => "11100011",7930 => "11010001",7931 => "11010101",7932 => "11001011",7933 => "00001101",7934 => "11100011",7935 => "10110001",7936 => "10011000",7937 => "01100101",7938 => "01101101",7939 => "00100010",7940 => "01101011",7941 => "11001100",7942 => "01001101",7943 => "11000100",7944 => "10110110",7945 => "10011101",7946 => "11111111",7947 => "00111101",7948 => "00100101",7949 => "00010100",7950 => "01110011",7951 => "01001111",7952 => "00101011",7953 => "01110100",7954 => "00110010",7955 => "01100100",7956 => "11010111",7957 => "10110100",7958 => "10111110",7959 => "10101011",7960 => "01110011",7961 => "11110001",7962 => "11001000",7963 => "00000001",7964 => "00111000",7965 => "01010011",7966 => "00010001",7967 => "11001100",7968 => "01010011",7969 => "00111110",7970 => "11011000",7971 => "11100000",7972 => "01011000",7973 => "10001100",7974 => "01100011",7975 => "10010110",7976 => "01101001",7977 => "01011100",7978 => "10010110",7979 => "10011100",7980 => "01110100",7981 => "11011010",7982 => "01010011",7983 => "11001000",7984 => "11001101",7985 => "11101000",7986 => "00101010",7987 => "00011010",7988 => "11010001",7989 => "00011010",7990 => "00001100",7991 => "11101101",7992 => "11000011",7993 => "00110100",7994 => "01011101",7995 => "10001111",7996 => "01011011",7997 => "00011010",7998 => "11001011",7999 => "00000110",8000 => "01110111",8001 => "11011101",8002 => "01110001",8003 => "00111100",8004 => "10001101",8005 => "01111100",8006 => "11010110",8007 => "00110110",8008 => "01100001",8009 => "11100111",8010 => "10100111",8011 => "11010101",8012 => "11100001",8013 => "11001100",8014 => "00101000",8015 => "01000111",8016 => "01100011",8017 => "01001000",8018 => "11001110",8019 => "11111001",8020 => "10111101",8021 => "11000010",8022 => "10100010",8023 => "11011000",8024 => "00110101",8025 => "00001001",8026 => "10001110",8027 => "01011010",8028 => "00111111",8029 => "10011011",8030 => "00001011",8031 => "11001110",8032 => "01110101",8033 => "00001110",8034 => "11011111",8035 => "00100110",8036 => "01111101",8037 => "10010101",8038 => "11110110",8039 => "11111001",8040 => "10011010",8041 => "00000101",8042 => "11010110",8043 => "10001111",8044 => "01111000",8045 => "11011000",8046 => "10000011",8047 => "01100001",8048 => "01101010",8049 => "00100111",8050 => "01011010",8051 => "01001011",8052 => "00000110",8053 => "11101101",8054 => "00011111",8055 => "10001110",8056 => "00011101",8057 => "10000101",8058 => "00011000",8059 => "01100110",8060 => "10011010",8061 => "01001010",8062 => "10000111",8063 => "00111111",8064 => "11101110",8065 => "00111110",8066 => "01001110",8067 => "11010011",8068 => "00000110",8069 => "11100111",8070 => "11001001",8071 => "10111100",8072 => "01001011",8073 => "11110011",8074 => "01000100",8075 => "11101000",8076 => "10010011",8077 => "10111000",8078 => "00110100",8079 => "00010000",8080 => "01010110",8081 => "01100011",8082 => "10100101",8083 => "10011011",8084 => "11101010",8085 => "10100110",8086 => "11010010",8087 => "11111010",8088 => "00011101",8089 => "10011001",8090 => "00111111",8091 => "00101010",8092 => "01111010",8093 => "00111000",8094 => "01000101",8095 => "11011100",8096 => "01101001",8097 => "00001010",8098 => "11000000",8099 => "11001110",8100 => "01011010",8101 => "01000000",8102 => "00010011",8103 => "11010011",8104 => "11110101",8105 => "00001100",8106 => "00010101",8107 => "00111011",8108 => "11111010",8109 => "01110110",8110 => "11111010",8111 => "01111101",8112 => "11001111",8113 => "11110110",8114 => "00000001",8115 => "00110101",8116 => "10110000",8117 => "01000101",8118 => "01101100",8119 => "11010100",8120 => "10000101",8121 => "11110000",8122 => "10100000",8123 => "10000001",8124 => "00110000",8125 => "01100011",8126 => "00010011",8127 => "11100100",8128 => "10001100",8129 => "11010010",8130 => "11100101",8131 => "10111000",8132 => "01010110",8133 => "11111000",8134 => "10011010",8135 => "11010101",8136 => "00110010",8137 => "11100000",8138 => "00001001",8139 => "11010100",8140 => "01011111",8141 => "00100000",8142 => "00010010",8143 => "00110000",8144 => "11010110",8145 => "10110100",8146 => "00011101",8147 => "11100101",8148 => "01100111",8149 => "01010010",8150 => "00100011",8151 => "11010000",8152 => "01010001",8153 => "11001100",8154 => "10000111",8155 => "11100000",8156 => "11010010",8157 => "11001101",8158 => "10111001",8159 => "11000111",8160 => "11011011",8161 => "11100001",8162 => "01010000",8163 => "10000110",8164 => "10101101",8165 => "00100010",8166 => "00110100",8167 => "01111000",8168 => "10010111",8169 => "00001011",8170 => "11010011",8171 => "01000111",8172 => "11110111",8173 => "10101011",8174 => "01011011",8175 => "11001001",8176 => "01000111",8177 => "01100110",8178 => "01011111",8179 => "10111010",8180 => "10010111",8181 => "00010010",8182 => "01011001",8183 => "00101110",8184 => "11010101",8185 => "00011101",8186 => "10110110",8187 => "00001111",8188 => "11000110",8189 => "11001010",8190 => "10100011",8191 => "10010010",8192 => "10110011",8193 => "10000010",8194 => "00001010",8195 => "10111110",8196 => "00101100",8197 => "00011101",8198 => "01000111",8199 => "10111001",8200 => "10000001",8201 => "00110101",8202 => "11111101",8203 => "10101101",8204 => "10010101",8205 => "11111110",8206 => "11011110",8207 => "10101001",8208 => "00111001",8209 => "00000010",8210 => "00011110",8211 => "00010100",8212 => "00100001",8213 => "10001010",8214 => "00011100",8215 => "00001010",8216 => "11010010",8217 => "00011010",8218 => "00001000",8219 => "11101111",8220 => "01001001",8221 => "11010001",8222 => "11011111",8223 => "00010000",8224 => "01000101",8225 => "01011111",8226 => "11001011",8227 => "10001000",8228 => "11101000",8229 => "01101101",8230 => "11010001",8231 => "11010011",8232 => "01000111",8233 => "00010000",8234 => "10001001",8235 => "10001101",8236 => "00000000",8237 => "00001111",8238 => "00111000",8239 => "00111000",8240 => "11101011",8241 => "11110101",8242 => "01011011",8243 => "11001101",8244 => "00111110",8245 => "10100101",8246 => "10000100",8247 => "00010101",8248 => "01011101",8249 => "01111011",8250 => "01000100",8251 => "10111010",8252 => "11000100",8253 => "01100111",8254 => "00101010",8255 => "10110101",8256 => "00010101",8257 => "01101010",8258 => "10010011",8259 => "10011100",8260 => "00110011",8261 => "00001001",8262 => "00000110",8263 => "00001010",8264 => "00001000",8265 => "01101011",8266 => "10010100",8267 => "01100011",8268 => "00110001",8269 => "00100000",8270 => "00011101",8271 => "01101010",8272 => "10100110",8273 => "00111010",8274 => "01100001",8275 => "01100111",8276 => "11010101",8277 => "01100101",8278 => "11101111",8279 => "11010101",8280 => "11000100",8281 => "00110111",8282 => "10000100",8283 => "11011000",8284 => "11001011",8285 => "11011101",8286 => "00110101",8287 => "00000001",8288 => "11111001",8289 => "01000111",8290 => "10101001",8291 => "11111111",8292 => "10111000",8293 => "11000101",8294 => "10100011",8295 => "00101111",8296 => "01101000",8297 => "01101001",8298 => "01111011",8299 => "00111111",8300 => "10101001",8301 => "01010111",8302 => "00111000",8303 => "01101111",8304 => "11010011",8305 => "00101100",8306 => "01100110",8307 => "11110001",8308 => "11010100",8309 => "10100001",8310 => "01010001",8311 => "00101000",8312 => "01101100",8313 => "11010011",8314 => "11010101",8315 => "00001001",8316 => "11011011",8317 => "01010001",8318 => "01001010",8319 => "11001000",8320 => "01001010",8321 => "10100101",8322 => "00110010",8323 => "00101011",8324 => "10011010",8325 => "11011000",8326 => "11001100",8327 => "11010101",8328 => "00101010",8329 => "01000111",8330 => "11001100",8331 => "00111111",8332 => "00101001",8333 => "11010111",8334 => "00111100",8335 => "00010000",8336 => "10100010",8337 => "00001000",8338 => "01000101",8339 => "00111101",8340 => "01010010",8341 => "01110111",8342 => "01001110",8343 => "00011101",8344 => "11101110",8345 => "00000001",8346 => "01000110",8347 => "01111011",8348 => "11011001",8349 => "10101000",8350 => "11010100",8351 => "10011001",8352 => "00110100",8353 => "01101001",8354 => "11110000",8355 => "00110111",8356 => "01111110",8357 => "10000010",8358 => "10000100",8359 => "01101010",8360 => "11101110",8361 => "10001010",8362 => "11011111",8363 => "11111001",8364 => "01110101",8365 => "01111011",8366 => "00000101",8367 => "10011000",8368 => "10101001",8369 => "00110000",8370 => "10000010",8371 => "10010011",8372 => "11001110",8373 => "00100000",8374 => "11100010",8375 => "01010011",8376 => "00011100",8377 => "01001111",8378 => "01010001",8379 => "00001000",8380 => "01101010",8381 => "00011011",8382 => "01101011",8383 => "11100101",8384 => "01000001",8385 => "00110011",8386 => "10111000",8387 => "01110010",8388 => "11010011",8389 => "01011100",8390 => "11110110",8391 => "10010100",8392 => "10111111",8393 => "01101100",8394 => "00011101",8395 => "01100100",8396 => "01010101",8397 => "00100111",8398 => "11010001",8399 => "10111010",8400 => "11111100",8401 => "00000000",8402 => "00111111",8403 => "01100111",8404 => "01101000",8405 => "11100011",8406 => "01101101",8407 => "01110011",8408 => "00010101",8409 => "00001001",8410 => "01011111",8411 => "00000110",8412 => "10001110",8413 => "10110001",8414 => "00000101",8415 => "10111111",8416 => "01010111",8417 => "10111111",8418 => "11111001",8419 => "10010100",8420 => "00011101",8421 => "10110100",8422 => "01000110",8423 => "01010000",8424 => "10011110",8425 => "11010111",8426 => "10000010",8427 => "10011011",8428 => "10100100",8429 => "11011001",8430 => "01100101",8431 => "11111100",8432 => "00110011",8433 => "00111010",8434 => "11110111",8435 => "00111010",8436 => "10010111",8437 => "01000101",8438 => "00110010",8439 => "10011001",8440 => "00010110",8441 => "11000110",8442 => "01000001",8443 => "11000011",8444 => "10100101",8445 => "10110110",8446 => "10001100",8447 => "10001010",8448 => "10001001",8449 => "00100101",8450 => "00110100",8451 => "11100110",8452 => "10101111",8453 => "00111010",8454 => "01010001",8455 => "11010000",8456 => "00101010",8457 => "01001100",8458 => "10011100",8459 => "00100101",8460 => "11000001",8461 => "00111000",8462 => "01110000",8463 => "00101110",8464 => "10001011",8465 => "10111010",8466 => "10100000",8467 => "00001000",8468 => "01101001",8469 => "00100000",8470 => "11011011",8471 => "10010110",8472 => "10011011",8473 => "00101101",8474 => "01111001",8475 => "00111010",8476 => "00010110",8477 => "10110101",8478 => "10010110",8479 => "01010011",8480 => "10101001",8481 => "01011001",8482 => "10011111",8483 => "10010100",8484 => "00100111",8485 => "00010100",8486 => "10100000",8487 => "01101011",8488 => "10101111",8489 => "00101011",8490 => "01111000",8491 => "10000001",8492 => "00110010",8493 => "10011111",8494 => "01101111",8495 => "10101111",8496 => "10100010",8497 => "00010010",8498 => "01011010",8499 => "01001000",8500 => "01101101",8501 => "01100111",8502 => "11001111",8503 => "11110110",8504 => "10110100",8505 => "11101101",8506 => "01101111",8507 => "10110101",8508 => "11110111",8509 => "00011101",8510 => "01110101",8511 => "01100000",8512 => "01111010",8513 => "00010111",8514 => "10100100",8515 => "11000111",8516 => "01000001",8517 => "11111111",8518 => "00011000",8519 => "01000111",8520 => "10010111",8521 => "01100110",8522 => "00001011",8523 => "10000111",8524 => "10011011",8525 => "11001001",8526 => "00110111",8527 => "00110100",8528 => "00101001",8529 => "01111100",8530 => "10111110",8531 => "01010001",8532 => "11101110",8533 => "11110110",8534 => "10010100",8535 => "11000011",8536 => "00000101",8537 => "10011110",8538 => "01001001",8539 => "10100101",8540 => "11101110",8541 => "01110010",8542 => "01110010",8543 => "10010001",8544 => "00010001",8545 => "01101111",8546 => "10001000",8547 => "11111011",8548 => "01010101",8549 => "01110001",8550 => "01100000",8551 => "00111111",8552 => "00110000",8553 => "10110011",8554 => "10101010",8555 => "00100101",8556 => "11100101",8557 => "10111101",8558 => "00011000",8559 => "11110100",8560 => "11111010",8561 => "10000010",8562 => "11101100",8563 => "00101010",8564 => "01000100",8565 => "01110101",8566 => "00000000",8567 => "10100011",8568 => "01111000",8569 => "10110110",8570 => "01101010",8571 => "01011011",8572 => "10001110",8573 => "01010110",8574 => "00000100",8575 => "10101010",8576 => "11100100",8577 => "11001111",8578 => "00001011",8579 => "11100100",8580 => "01010001",8581 => "11000110",8582 => "10101110",8583 => "11101111",8584 => "01111111",8585 => "01001111",8586 => "01011011",8587 => "11110010",8588 => "00001101",8589 => "11010001",8590 => "10111000",8591 => "01010100",8592 => "00100000",8593 => "00011001",8594 => "00101100",8595 => "11111110",8596 => "11011110",8597 => "01100001",8598 => "10001010",8599 => "11111001",8600 => "01110011",8601 => "01101000",8602 => "11100101",8603 => "01101000",8604 => "10110110",8605 => "01011010",8606 => "11000100",8607 => "01000000",8608 => "10110000",8609 => "11000101",8610 => "01101001",8611 => "00001000",8612 => "10011101",8613 => "01110110",8614 => "01111011",8615 => "11111111",8616 => "00100100",8617 => "11001011",8618 => "10100000",8619 => "11001111",8620 => "10011100",8621 => "11101011",8622 => "00101001",8623 => "11000010",8624 => "11010110",8625 => "01111011",8626 => "01011110",8627 => "10101001",8628 => "11000001",8629 => "01111001",8630 => "11011100",8631 => "00000100",8632 => "00011001",8633 => "01000110",8634 => "00000000",8635 => "10101000",8636 => "00110101",8637 => "00000101",8638 => "01010110",8639 => "10001110",8640 => "00101110",8641 => "00101111",8642 => "10110100",8643 => "11011111",8644 => "10101000",8645 => "00110100",8646 => "00111010",8647 => "00111111",8648 => "01011011",8649 => "00011111",8650 => "00111100",8651 => "00001101",8652 => "01000000",8653 => "01000000",8654 => "10011101",8655 => "10010101",8656 => "11011111",8657 => "00111000",8658 => "00101001",8659 => "01101001",8660 => "10111111",8661 => "11010001",8662 => "00001011",8663 => "01011100",8664 => "01100111",8665 => "11111110",8666 => "10100000",8667 => "01101010",8668 => "01011001",8669 => "01010101",8670 => "01000011",8671 => "10110100",8672 => "00101011",8673 => "11000100",8674 => "00010000",8675 => "10001110",8676 => "01011110",8677 => "01011001",8678 => "11110010",8679 => "10100101",8680 => "00101010",8681 => "00110100",8682 => "01010111",8683 => "01011000",8684 => "00000010",8685 => "10111010",8686 => "10011010",8687 => "00010100",8688 => "10011001",8689 => "11001011",8690 => "00001101",8691 => "11000010",8692 => "01001001",8693 => "00110001",8694 => "11111001",8695 => "11001100",8696 => "11000101",8697 => "00110011",8698 => "01100010",8699 => "10101001",8700 => "11101111",8701 => "00001000",8702 => "00110110",8703 => "10010100",8704 => "10011111",8705 => "00010000",8706 => "01100000",8707 => "01010110",8708 => "11010010",8709 => "10110011",8710 => "01110011",8711 => "10001100",8712 => "11011111",8713 => "11011100",8714 => "11100010",8715 => "11011001",8716 => "00010010",8717 => "01001010",8718 => "00000110",8719 => "00011010",8720 => "01010001",8721 => "00101000",8722 => "10111000",8723 => "11111001",8724 => "11000001",8725 => "00100011",8726 => "11110101",8727 => "00000011",8728 => "11011011",8729 => "00111110",8730 => "01011110",8731 => "10000101",8732 => "10101111",8733 => "10011100",8734 => "01011110",8735 => "00000110",8736 => "01010111",8737 => "11011010",8738 => "11111101",8739 => "11110010",8740 => "01010011",8741 => "00101101",8742 => "10000111",8743 => "01101110",8744 => "10100011",8745 => "00000100",8746 => "10110110",8747 => "01010011",8748 => "10010101",8749 => "00000000",8750 => "10110110",8751 => "10011101",8752 => "10010010",8753 => "00111011",8754 => "10111100",8755 => "11000011",8756 => "01001000",8757 => "01001100",8758 => "01010111",8759 => "01000001",8760 => "00001011",8761 => "01110010",8762 => "01010001",8763 => "10000001",8764 => "00110001",8765 => "11110101",8766 => "00011000",8767 => "10101010",8768 => "11001110",8769 => "11001101",8770 => "01110000",8771 => "00101100",8772 => "11011110",8773 => "10101010",8774 => "11100100",8775 => "11011110",8776 => "01100011",8777 => "00100101",8778 => "10001010",8779 => "00011110",8780 => "11100010",8781 => "00100101",8782 => "00100011",8783 => "11101101",8784 => "00111001",8785 => "01100110",8786 => "11101011",8787 => "11000101",8788 => "00001110",8789 => "01111111",8790 => "10000110",8791 => "10100101",8792 => "01011000",8793 => "11100010",8794 => "10110010",8795 => "00000010",8796 => "11110111",8797 => "10111100",8798 => "00110101",8799 => "00010011",8800 => "10000101",8801 => "00110101",8802 => "11100000",8803 => "00001110",8804 => "01101100",8805 => "10100111",8806 => "01011011",8807 => "11010000",8808 => "00100101",8809 => "01111010",8810 => "11001110",8811 => "01001000",8812 => "00111011",8813 => "11101101",8814 => "11011011",8815 => "01001010",8816 => "10001110",8817 => "00101000",8818 => "01111011",8819 => "11111001",8820 => "01000000",8821 => "00101010",8822 => "01111001",8823 => "01111011",8824 => "10001001",8825 => "01101101",8826 => "11001110",8827 => "10010001",8828 => "10101010",8829 => "00011000",8830 => "01011100",8831 => "00001010",8832 => "11100101",8833 => "11001010",8834 => "11001011",8835 => "00100010",8836 => "10110111",8837 => "10100001",8838 => "11111100",8839 => "01001001",8840 => "10011001",8841 => "11011110",8842 => "01011001",8843 => "00001101",8844 => "00101011",8845 => "00001110",8846 => "10101111",8847 => "00101110",8848 => "00100001",8849 => "10011110",8850 => "10110001",8851 => "10101100",8852 => "10001111",8853 => "10001101",8854 => "01011100",8855 => "10001011",8856 => "10110110",8857 => "10010010",8858 => "01010110",8859 => "11010111",8860 => "00010101",8861 => "01010011",8862 => "11010111",8863 => "01111001",8864 => "00110011",8865 => "00000000",8866 => "11111011",8867 => "10001010",8868 => "10101101",8869 => "11101011",8870 => "10101010",8871 => "00010000",8872 => "00000010",8873 => "01110011",8874 => "00001111",8875 => "10010101",8876 => "00000111",8877 => "11111100",8878 => "00000101",8879 => "00111101",8880 => "10111011",8881 => "11010011",8882 => "11001100",8883 => "10101001",8884 => "11101110",8885 => "00000110",8886 => "01000111",8887 => "11100011",8888 => "10110001",8889 => "10100101",8890 => "11111111",8891 => "10010011",8892 => "01110010",8893 => "01111010",8894 => "11111111",8895 => "00000011",8896 => "10110101",8897 => "11011001",8898 => "11101000",8899 => "10111001",8900 => "10100001",8901 => "11100000",8902 => "00110001",8903 => "01110011",8904 => "11100000",8905 => "01110100",8906 => "10101000",8907 => "01001110",8908 => "01011001",8909 => "11111100",8910 => "00010011",8911 => "10000101",8912 => "00100011",8913 => "00010101",8914 => "11101010",8915 => "00000100",8916 => "10011011",8917 => "01110000",8918 => "10010011",8919 => "01011000",8920 => "01000100",8921 => "01010001",8922 => "11110011",8923 => "01000100",8924 => "11101111",8925 => "00011100",8926 => "10000100",8927 => "01010011",8928 => "00011010",8929 => "11001010",8930 => "01100010",8931 => "01110101",8932 => "10000011",8933 => "01001010",8934 => "11011100",8935 => "10000110",8936 => "11001011",8937 => "01101001",8938 => "11110001",8939 => "00111010",8940 => "01110111",8941 => "10010111",8942 => "11001101",8943 => "11111000",8944 => "11110000",8945 => "10000101",8946 => "10110111",8947 => "10100110",8948 => "11111001",8949 => "10000101",8950 => "01000001",8951 => "01011100",8952 => "00100111",8953 => "11101110",8954 => "01101110",8955 => "00100100",8956 => "00001101",8957 => "10111001",8958 => "00000000",8959 => "01100011",8960 => "01010011",8961 => "10010011",8962 => "10100000",8963 => "10111111",8964 => "11101110",8965 => "10110000",8966 => "00111101",8967 => "01111000",8968 => "00100010",8969 => "11100110",8970 => "10000010",8971 => "11110110",8972 => "00111110",8973 => "10100011",8974 => "11010011",8975 => "11011100",8976 => "00111000",8977 => "00110011",8978 => "00011001",8979 => "11110110",8980 => "11100011",8981 => "10111100",8982 => "11100000",8983 => "10101101",8984 => "01110100",8985 => "11001111",8986 => "00010110",8987 => "00010111",8988 => "10011110",8989 => "10000110",8990 => "11000111",8991 => "11101100",8992 => "00001100",8993 => "11000010",8994 => "10000100",8995 => "01011011",8996 => "01011010",8997 => "00100010",8998 => "00101011",8999 => "10001001",9000 => "00010110",9001 => "01101011",9002 => "01110010",9003 => "01100001",9004 => "01011110",9005 => "00011111",9006 => "01110100",9007 => "11011111",9008 => "01000101",9009 => "00010001",9010 => "10110001",9011 => "10011101",9012 => "11111101",9013 => "10101010",9014 => "00011001",9015 => "10110100",9016 => "10011011",9017 => "00000001",9018 => "00011100",9019 => "00100001",9020 => "10111110",9021 => "10101110",9022 => "01001100",9023 => "11001101",9024 => "00110011",9025 => "10000011",9026 => "01001111",9027 => "11010001",9028 => "10100110",9029 => "01101100",9030 => "00001010",9031 => "10010011",9032 => "00100010",9033 => "01010111",9034 => "11101000",9035 => "10001100",9036 => "01011110",9037 => "01111101",9038 => "00000100",9039 => "11011011",9040 => "10100000",9041 => "00110000",9042 => "10001000",9043 => "01010011",9044 => "10000111",9045 => "10111011",9046 => "01111001",9047 => "01111000",9048 => "00110010",9049 => "10110110",9050 => "10001011",9051 => "11110110",9052 => "11011011",9053 => "00100100",9054 => "11110101",9055 => "00110101",9056 => "00110110",9057 => "00011011",9058 => "10010100",9059 => "11011100",9060 => "01111110",9061 => "10001010",9062 => "00110111",9063 => "11010101",9064 => "01100101",9065 => "10110000",9066 => "11101001",9067 => "00111101",9068 => "10010011",9069 => "11010001",9070 => "10100100",9071 => "10110011",9072 => "01101111",9073 => "01100101",9074 => "00010110",9075 => "11011001",9076 => "00001000",9077 => "01000111",9078 => "01101110",9079 => "00101110",9080 => "11110010",9081 => "10001010",9082 => "10111101",9083 => "11001111",9084 => "00000001",9085 => "11111110",9086 => "10001100",9087 => "10001001",9088 => "00010001",9089 => "01000010",9090 => "11001101",9091 => "11101100",9092 => "01010011",9093 => "01110111",9094 => "00101010",9095 => "01010011",9096 => "01010010",9097 => "00010001",9098 => "00100100",9099 => "10011100",9100 => "01111101",9101 => "10111100",9102 => "00111100",9103 => "10100100",9104 => "10010001",9105 => "11101001",9106 => "11000010",9107 => "10001001",9108 => "10111001",9109 => "11011000",9110 => "00101011",9111 => "00011001",9112 => "01111011",9113 => "11111000",9114 => "00101110",9115 => "11100000",9116 => "11010111",9117 => "00111100",9118 => "01110011",9119 => "10010101",9120 => "11011000",9121 => "11110000",9122 => "01110111",9123 => "10001000",9124 => "10110011",9125 => "10010011",9126 => "10111000",9127 => "10110101",9128 => "10111011",9129 => "10101100",9130 => "01011110",9131 => "00100010",9132 => "00011010",9133 => "11000001",9134 => "01000000",9135 => "11111100",9136 => "01000110",9137 => "11111010",9138 => "00011010",9139 => "10010011",9140 => "00001111",9141 => "10101101",9142 => "01111000",9143 => "01101011",9144 => "01011010",9145 => "01101110",9146 => "00001101",9147 => "01111010",9148 => "01010101",9149 => "11000100",9150 => "10101000",9151 => "01010100",9152 => "00001111",9153 => "00011011",9154 => "01010010",9155 => "10110001",9156 => "00010111",9157 => "00100001",9158 => "01101100",9159 => "01111101",9160 => "00011100",9161 => "10011011",9162 => "00100110",9163 => "01010001",9164 => "11110101",9165 => "00101010",9166 => "00011101",9167 => "10000100",9168 => "00011101",9169 => "01100000",9170 => "01011101",9171 => "10000000",9172 => "00101010",9173 => "11111110",9174 => "00001111",9175 => "00010010",9176 => "10111110",9177 => "11000000",9178 => "10011000",9179 => "00011001",9180 => "11011100",9181 => "11010100",9182 => "11101000",9183 => "11100110",9184 => "01000100",9185 => "10001100",9186 => "11000110",9187 => "01001110",9188 => "11001110",9189 => "00010000",9190 => "11101011",9191 => "11010001",9192 => "10101111",9193 => "00001010",9194 => "00110111",9195 => "01100110",9196 => "01111001",9197 => "00010001",9198 => "01001111",9199 => "00111001",9200 => "00000111",9201 => "01110011",9202 => "01000011",9203 => "10011100",9204 => "10010110",9205 => "11011010",9206 => "11110101",9207 => "11100011",9208 => "01100101",9209 => "00011011",9210 => "10010101",9211 => "10111011",9212 => "01000111",9213 => "10101001",9214 => "11111000",9215 => "00100100",9216 => "11011110",9217 => "11110000",9218 => "01001110",9219 => "00001001",9220 => "00111100",9221 => "00110110",9222 => "10001010",9223 => "01101101",9224 => "01010110",9225 => "11000101",9226 => "01010000",9227 => "00001110",9228 => "00100001",9229 => "01101101",9230 => "00010000",9231 => "11000100",9232 => "11001111",9233 => "00101001",9234 => "01011000",9235 => "00001100",9236 => "10111000",9237 => "01110111",9238 => "00111101",9239 => "01011011",9240 => "10111000",9241 => "00001001",9242 => "00010000",9243 => "11101111",9244 => "11011101",9245 => "11001100",9246 => "10001000",9247 => "10001010",9248 => "00000111",9249 => "01100011",9250 => "10000000",9251 => "01000110",9252 => "01110111",9253 => "11010010",9254 => "00010100",9255 => "11110111",9256 => "10110111",9257 => "11100000",9258 => "11001110",9259 => "11111110",9260 => "10001000",9261 => "11000000",9262 => "10101100",9263 => "11111110",9264 => "10101101",9265 => "01011000",9266 => "10000111",9267 => "00001100",9268 => "00101100",9269 => "10000100",9270 => "10011001",9271 => "01011100",9272 => "01100010",9273 => "10111110",9274 => "11010010",9275 => "00100001",9276 => "10010110",9277 => "00011100",9278 => "01111100",9279 => "00000111",9280 => "00011100",9281 => "10011110",9282 => "11010001",9283 => "01101001",9284 => "10001100",9285 => "10010111",9286 => "01001110",9287 => "00011011",9288 => "11101100",9289 => "11010010",9290 => "10000011",9291 => "01011011",9292 => "00110000",9293 => "10000001",9294 => "11101000",9295 => "10101100",9296 => "01011111",9297 => "11011011",9298 => "00100010",9299 => "01100011",9300 => "11000110",9301 => "11000111",9302 => "11100001",9303 => "10100100",9304 => "00011111",9305 => "01000001",9306 => "10101100",9307 => "00110011",9308 => "11101110",9309 => "00001111",9310 => "01010000",9311 => "10011001",9312 => "00100001",9313 => "11111110",9314 => "01001101",9315 => "01100001",9316 => "10101001",9317 => "00100010",9318 => "01001011",9319 => "11010000",9320 => "11110100",9321 => "11110011",9322 => "11100110",9323 => "10000001",9324 => "01011110",9325 => "10111111",9326 => "11111010",9327 => "10111010",9328 => "10010011",9329 => "10111111",9330 => "01000010",9331 => "11111111",9332 => "00011101",9333 => "10110100",9334 => "11010111",9335 => "10100010",9336 => "00110100",9337 => "10100011",9338 => "10000111",9339 => "01010100",9340 => "10111010",9341 => "00010001",9342 => "10000110",9343 => "10100001",9344 => "11001011",9345 => "01110010",9346 => "11011101",9347 => "11100001",9348 => "00011101",9349 => "00100100",9350 => "01100110",9351 => "01111111",9352 => "11011000",9353 => "00111101",9354 => "01110101",9355 => "01001010",9356 => "11001000",9357 => "10110101",9358 => "01010100",9359 => "10111011",9360 => "11000110",9361 => "00111101",9362 => "01111001",9363 => "10000100",9364 => "11100000",9365 => "10011011",9366 => "01011111",9367 => "11001111",9368 => "11101100",9369 => "01000111",9370 => "00001010",9371 => "10010011",9372 => "01001110",9373 => "10000001",9374 => "00101111",9375 => "11001010",9376 => "00000001",9377 => "11001101",9378 => "10100111",9379 => "10111111",9380 => "11000011",9381 => "10100001",9382 => "01101011",9383 => "00100100",9384 => "01011110",9385 => "00010100",9386 => "00101111",9387 => "01010001",9388 => "11110001",9389 => "01010011",9390 => "01111010",9391 => "01111000",9392 => "01110011",9393 => "01101111",9394 => "00111110",9395 => "11000010",9396 => "00000100",9397 => "10001110",9398 => "01100001",9399 => "10011001",9400 => "00010101",9401 => "10011000",9402 => "11100011",9403 => "10011110",9404 => "10001000",9405 => "11001001",9406 => "11010100",9407 => "11001011",9408 => "01010011",9409 => "10011011",9410 => "10111110",9411 => "10111100",9412 => "01011110",9413 => "10001001",9414 => "11010011",9415 => "01001110",9416 => "01010010",9417 => "01000100",9418 => "01101000",9419 => "11110011",9420 => "11010100",9421 => "00011010",9422 => "01101100",9423 => "10000110",9424 => "00001001",9425 => "10001000",9426 => "01010000",9427 => "11110011",9428 => "11101000",9429 => "00011001",9430 => "01001101",9431 => "01001100",9432 => "00100001",9433 => "11111110",9434 => "01101000",9435 => "10100011",9436 => "10100010",9437 => "10110001",9438 => "00010001",9439 => "11100001",9440 => "00101110",9441 => "10100101",9442 => "00110110",9443 => "11101111",9444 => "11110001",9445 => "10100010",9446 => "00111010",9447 => "00000000",9448 => "11000110",9449 => "01100001",9450 => "00010110",9451 => "11101100",9452 => "10000010",9453 => "01111110",9454 => "01001101",9455 => "11101101",9456 => "00011010",9457 => "11000110",9458 => "01111001",9459 => "11001101",9460 => "10001110",9461 => "11001100",9462 => "10111111",9463 => "01110100",9464 => "00001100",9465 => "00011000",9466 => "10010110",9467 => "01100111",9468 => "11100110",9469 => "01111100",9470 => "00010100",9471 => "01101110",9472 => "10111010",9473 => "10001100",9474 => "11111100",9475 => "01000110",9476 => "10100100",9477 => "10001010",9478 => "10011111",9479 => "10010110",9480 => "01100000",9481 => "01110110",9482 => "10111111",9483 => "01110011",9484 => "00110100",9485 => "11100100",9486 => "00001001",9487 => "00000111",9488 => "11001111",9489 => "01000100",9490 => "00111110",9491 => "10100111",9492 => "11000000",9493 => "01001011",9494 => "00011101",9495 => "10110100",9496 => "10010111",9497 => "01111011",9498 => "11011110",9499 => "10111011",9500 => "11100000",9501 => "00000000",9502 => "10101111",9503 => "11110111",9504 => "11111110",9505 => "00000000",9506 => "11001111",9507 => "10111010",9508 => "00100111",9509 => "11100100",9510 => "10001011",9511 => "11000100",9512 => "10001101",9513 => "11001110",9514 => "10010011",9515 => "10111100",9516 => "01100001",9517 => "00000001",9518 => "11000010",9519 => "11111111",9520 => "01001110",9521 => "00001000",9522 => "00010000",9523 => "11001001",9524 => "10100001",9525 => "10101111",9526 => "11100001",9527 => "01001101",9528 => "10101101",9529 => "11001101",9530 => "11011111",9531 => "11011101",9532 => "01111001",9533 => "10011101",9534 => "10101001",9535 => "01111011",9536 => "11101110",9537 => "11000010",9538 => "01101110",9539 => "11001111",9540 => "11000000",9541 => "10110000",9542 => "01100011",9543 => "10000110",9544 => "00010001",9545 => "00100010",9546 => "01100110",9547 => "11010111",9548 => "00000011",9549 => "01101110",9550 => "00111111",9551 => "00111000",9552 => "11010011",9553 => "00101010",9554 => "10000100",9555 => "00100111",9556 => "11111001",9557 => "00101110",9558 => "00101110",9559 => "01101011",9560 => "11111010",9561 => "11000011",9562 => "10101010",9563 => "11011110",9564 => "10111001",9565 => "01000000",9566 => "10001101",9567 => "10110011",9568 => "11101010",9569 => "10000011",9570 => "01010110",9571 => "00101101",9572 => "10011101",9573 => "10100110",9574 => "00011011",9575 => "01010101",9576 => "11110111",9577 => "00010110",9578 => "00111100",9579 => "10001010",9580 => "01010001",9581 => "00100001",9582 => "11001110",9583 => "01000010",9584 => "00011011",9585 => "01001101",9586 => "01011110",9587 => "00100111",9588 => "11011101",9589 => "01100111",9590 => "00000100",9591 => "01011101",9592 => "00001100",9593 => "00100101",9594 => "00110000",9595 => "11001010",9596 => "11100001",9597 => "10111110",9598 => "11010011",9599 => "01011101",9600 => "11101101",9601 => "01000101",9602 => "00100101",9603 => "01001110",9604 => "11111100",9605 => "00010010",9606 => "11001111",9607 => "11100100",9608 => "00101001",9609 => "11100111",9610 => "00010101",9611 => "01011110",9612 => "01100011",9613 => "00000011",9614 => "00111101",9615 => "10100001",9616 => "01110000",9617 => "00001110",9618 => "11001000",9619 => "10110011",9620 => "10001000",9621 => "10110001",9622 => "11100000",9623 => "01000011",9624 => "01100100",9625 => "11000010",9626 => "00010000",9627 => "00101100",9628 => "10110111",9629 => "00000101",9630 => "01000110",9631 => "01000000",9632 => "10010111",9633 => "11100010",9634 => "11010101",9635 => "11100000",9636 => "01110010",9637 => "11000010",9638 => "10001001",9639 => "10100010",9640 => "10001101",9641 => "00110001",9642 => "10001010",9643 => "10001110",9644 => "10101001",9645 => "10010000",9646 => "01110110",9647 => "00001001",9648 => "10000100",9649 => "10110110",9650 => "10100101",9651 => "00100111",9652 => "10000100",9653 => "00110111",9654 => "01001000",9655 => "01010010",9656 => "00001110",9657 => "01001110",9658 => "00011111",9659 => "10011100",9660 => "01100011",9661 => "10001010",9662 => "10010000",9663 => "01111101",9664 => "00000111",9665 => "10011010",9666 => "11110101",9667 => "01110101",9668 => "01001001",9669 => "01100011",9670 => "01010110",9671 => "10100010",9672 => "00000001",9673 => "01100111",9674 => "11000111",9675 => "01100010",9676 => "00010000",9677 => "11101011",9678 => "10111000",9679 => "00011000",9680 => "10000100",9681 => "01011000",9682 => "11001111",9683 => "01110110",9684 => "01111000",9685 => "01111100",9686 => "10110001",9687 => "01111010",9688 => "10001010",9689 => "11000010",9690 => "01001011",9691 => "11101011",9692 => "01000000",9693 => "01110101",9694 => "00000010",9695 => "10011011",9696 => "00111000",9697 => "10110100",9698 => "11011010",9699 => "10000100",9700 => "00100110",9701 => "01000010",9702 => "01111000",9703 => "10010100",9704 => "11110011",9705 => "11011011",9706 => "01011000",9707 => "00111110",9708 => "10100011",9709 => "00100011",9710 => "10000001",9711 => "00110001",9712 => "10000101",9713 => "01000001",9714 => "10010110",9715 => "10110111",9716 => "00111011",9717 => "01010110",9718 => "11110110",9719 => "01100011",9720 => "00011001",9721 => "10010000",9722 => "00100101",9723 => "00010111",9724 => "01110101",9725 => "00000101",9726 => "00000010",9727 => "11011100",9728 => "11101101",9729 => "11011110",9730 => "10111101",9731 => "10111111",9732 => "10101011",9733 => "00110101",9734 => "00011011",9735 => "00100110",9736 => "01000000",9737 => "01010100",9738 => "11010001",9739 => "00101010",9740 => "01111000",9741 => "11000110",9742 => "01000100",9743 => "00101111",9744 => "11001010",9745 => "00000111",9746 => "10101101",9747 => "00000001",9748 => "10001010",9749 => "10011001",9750 => "11110100",9751 => "01001010",9752 => "00111110",9753 => "01111000",9754 => "11100010",9755 => "01001001",9756 => "11011110",9757 => "11101011",9758 => "10111000",9759 => "10010000",9760 => "11000000",9761 => "01110101",9762 => "10110010",9763 => "01000110",9764 => "00011000",9765 => "01110010",9766 => "01001111",9767 => "11111101",9768 => "01001111",9769 => "01100001",9770 => "11000000",9771 => "01111110",9772 => "10101001",9773 => "10101100",9774 => "11000000",9775 => "11110001",9776 => "10010001",9777 => "11001110",9778 => "00110110",9779 => "01101101",9780 => "11111000",9781 => "10011000",9782 => "11010110",9783 => "11010010",9784 => "00100101",9785 => "00010000",9786 => "11100110",9787 => "10110000",9788 => "10100001",9789 => "10100011",9790 => "11111000",9791 => "01000011",9792 => "10100010",9793 => "11011110",9794 => "00011001",9795 => "01100010",9796 => "10010010",9797 => "10111100",9798 => "10011000",9799 => "01000000",9800 => "10110010",9801 => "10101001",9802 => "00100000",9803 => "10110100",9804 => "01010010",9805 => "10100100",9806 => "11110111",9807 => "11111000",9808 => "10000111",9809 => "00101110",9810 => "11100011",9811 => "01110100",9812 => "00101010",9813 => "00110100",9814 => "01000010",9815 => "11000001",9816 => "00110100",9817 => "10101000",9818 => "10110001",9819 => "11001011",9820 => "00110101",9821 => "10011100",9822 => "01101100",9823 => "10100110",9824 => "00001100",9825 => "11100001",9826 => "10101001",9827 => "01000110",9828 => "11001111",9829 => "10000101",9830 => "01001001",9831 => "10010101",9832 => "10000100",9833 => "00000101",9834 => "00001011",9835 => "01011100",9836 => "10000100",9837 => "11111011",9838 => "00011110",9839 => "10110001",9840 => "01110000",9841 => "11100100",9842 => "10100000",9843 => "00000110",9844 => "01000010",9845 => "10001011",9846 => "01010100",9847 => "10100011",9848 => "00000111",9849 => "00111000",9850 => "01011011",9851 => "01100001",9852 => "00100000",9853 => "11101001",9854 => "00111000",9855 => "01100011",9856 => "01100111",9857 => "10100111",9858 => "10110001",9859 => "01010010",9860 => "11100111",9861 => "01011011",9862 => "00011100",9863 => "11001110",9864 => "00111000",9865 => "11101100",9866 => "01011010",9867 => "01111100",9868 => "01111001",9869 => "00100011",9870 => "11101011",9871 => "10110110",9872 => "10000000",9873 => "11101110",9874 => "11010011",9875 => "10011011",9876 => "01000011",9877 => "10110000",9878 => "01110011",9879 => "01101001",9880 => "10110000",9881 => "01101101",9882 => "01111110",9883 => "00011110",9884 => "00000000",9885 => "00110010",9886 => "00011001",9887 => "00011111",9888 => "00000101",9889 => "00100101",9890 => "11111111",9891 => "01001100",9892 => "00111100",9893 => "10010011",9894 => "10111011",9895 => "00110110",9896 => "01111110",9897 => "10001100",9898 => "01101001",9899 => "01110111",9900 => "10111011",9901 => "10101111",9902 => "01111010",9903 => "10110110",9904 => "00011000",9905 => "10011101",9906 => "10101101",9907 => "01010000",9908 => "11100011",9909 => "10000001",9910 => "00110000",9911 => "00100100",9912 => "10100011",9913 => "01101100",9914 => "10111101",9915 => "11000010",9916 => "00010001",9917 => "10000101",9918 => "00101011",9919 => "00000101",9920 => "01100100",9921 => "10111010",9922 => "00001000",9923 => "00111010",9924 => "11000100",9925 => "01100010",9926 => "11100000",9927 => "00011000",9928 => "00001111",9929 => "11101110",9930 => "11011101",9931 => "01001101",9932 => "00011111",9933 => "01010010",9934 => "00110011",9935 => "11000100",9936 => "01111101",9937 => "11000000",9938 => "01110001",9939 => "11111101",9940 => "01010110",9941 => "01110101",9942 => "01000000",9943 => "01010110",9944 => "11000100",9945 => "10110000",9946 => "01000011",9947 => "00000101",9948 => "11010110",9949 => "11011101",9950 => "01101111",9951 => "10100100",9952 => "01101011",9953 => "10111110",9954 => "10100011",9955 => "01110011",9956 => "01110010",9957 => "11001011",9958 => "01001111",9959 => "11110100",9960 => "00110110",9961 => "10111111",9962 => "10111111",9963 => "01000100",9964 => "10010111",9965 => "11011100",9966 => "10110010",9967 => "01010101",9968 => "11000010",9969 => "10111001",9970 => "11111010",9971 => "10100010",9972 => "10001111",9973 => "01110111",9974 => "11000111",9975 => "10101010",9976 => "11100001",9977 => "01101011",9978 => "11000001",9979 => "00111010",9980 => "00011011",9981 => "01011010",9982 => "00011000",9983 => "01100011",9984 => "10110011",9985 => "11000011",9986 => "01111110",9987 => "01110111",9988 => "11110101",9989 => "11110011",9990 => "01001101",9991 => "11011100",9992 => "10011011",9993 => "10111000",9994 => "01001010",9995 => "00111000",9996 => "10011001",9997 => "00100101",9998 => "10101101",9999 => "11000100",10000 => "10100000",10001 => "00001011",10002 => "10011011",10003 => "00001010",10004 => "11101101",10005 => "00000001",10006 => "00000101",10007 => "11010001",10008 => "00000000",10009 => "10101011",10010 => "11011001",10011 => "10100111",10012 => "00000011",10013 => "00110000",10014 => "10000011",10015 => "00110000",10016 => "01101010",10017 => "10111110",10018 => "11000011",10019 => "00011111",10020 => "11111110",10021 => "00111100",10022 => "01101100",10023 => "01001100",10024 => "01111101",10025 => "11110110",10026 => "00111100",10027 => "10011111",10028 => "00001010",10029 => "11010110",10030 => "01011100",10031 => "10111111",10032 => "01111001",10033 => "01101011",10034 => "00010110",10035 => "01010110",10036 => "01011011",10037 => "00111110",10038 => "10010001",10039 => "10000001",10040 => "11011010",10041 => "10100011",10042 => "01011001",10043 => "11000111",10044 => "01111010",10045 => "11010010",10046 => "11101011",10047 => "10111001",10048 => "10011011",10049 => "00000001",10050 => "01111110",10051 => "01001001",10052 => "00101011",10053 => "10010001",10054 => "01001110",10055 => "11000101",10056 => "11001011",10057 => "01100100",10058 => "00110111",10059 => "00000111",10060 => "10110101",10061 => "00101101",10062 => "11101100",10063 => "01010100",10064 => "00100000",10065 => "01111001",10066 => "11001001",10067 => "01001010",10068 => "01011101",10069 => "00101000",10070 => "10001111",10071 => "00001101",10072 => "00010011",10073 => "10000010",10074 => "10101101",10075 => "10000101",10076 => "01011011",10077 => "00001101",10078 => "10100011",10079 => "01010100",10080 => "01110111",10081 => "10010111",10082 => "00101000",10083 => "00001110",10084 => "10101011",10085 => "01010100",10086 => "11111111",10087 => "10101101",10088 => "00100000",10089 => "01101100",10090 => "10010100",10091 => "00111000",10092 => "01100010",10093 => "10110110",10094 => "10100110",10095 => "10110110",10096 => "10100100",10097 => "11110010",10098 => "10001100",10099 => "10000100",10100 => "11001111",10101 => "10100101",10102 => "01111011",10103 => "10101100",10104 => "11101100",10105 => "10001000",10106 => "01101100",10107 => "10111101",10108 => "11000100",10109 => "00111110",10110 => "11010110",10111 => "11001100",10112 => "11000111",10113 => "11110000",10114 => "01001111",10115 => "10100110",10116 => "01101101",10117 => "11000101",10118 => "00011001",10119 => "00010110",10120 => "11000000",10121 => "00011010",10122 => "00110010",10123 => "11111010",10124 => "01101110",10125 => "00011010",10126 => "10000011",10127 => "01011111",10128 => "10101011",10129 => "00111101",10130 => "00111010",10131 => "11001100",10132 => "01001100",10133 => "11000101",10134 => "10100100",10135 => "10010101",10136 => "00000000",10137 => "01101111",10138 => "10100010",10139 => "10000011",10140 => "00011100",10141 => "01011101",10142 => "00011100",10143 => "01010001",10144 => "00111111",10145 => "01010010",10146 => "10100001",10147 => "10111010",10148 => "11100001",10149 => "00011111",10150 => "10000000",10151 => "11110000",10152 => "10000101",10153 => "00110110",10154 => "01100100",10155 => "10010111",10156 => "10100011",10157 => "10101000",10158 => "10101011",10159 => "01101010",10160 => "00111101",10161 => "11011101",10162 => "10110110",10163 => "11011011",10164 => "00010011",10165 => "11100000",10166 => "10011111",10167 => "01001011",10168 => "01000001",10169 => "00100111",10170 => "01011011",10171 => "10101001",10172 => "01011010",10173 => "11111101",10174 => "10011101",10175 => "01000000",10176 => "01111010",10177 => "10011000",10178 => "11011010",10179 => "11011101",10180 => "00001110",10181 => "00001110",10182 => "00100111",10183 => "00000000",10184 => "01100110",10185 => "00110101",10186 => "00000001",10187 => "10011001",10188 => "11101110",10189 => "10101010",10190 => "01001001",10191 => "01110100",10192 => "01101011",10193 => "00110010",10194 => "11011010",10195 => "10110101",10196 => "00111100",10197 => "11011000",10198 => "10111101",10199 => "10100101",10200 => "01000111",10201 => "00001101",10202 => "00101110",10203 => "11101000",10204 => "00000000",10205 => "11001100",10206 => "01010101",10207 => "01011011",10208 => "00010111",10209 => "01001100",10210 => "11110111",10211 => "01110101",10212 => "00101110",10213 => "00011101",10214 => "00101001",10215 => "10001011",10216 => "01010000",10217 => "10011011",10218 => "00110001",10219 => "00000001",10220 => "01101100",10221 => "01010111",10222 => "10011000",10223 => "01001111",10224 => "01000110",10225 => "00011000",10226 => "01000010",10227 => "00010000",10228 => "01110100",10229 => "10011000",10230 => "11110111",10231 => "11010010",10232 => "11000101",10233 => "10010111",10234 => "11001011",10235 => "00010011",10236 => "00101000",10237 => "00010111",10238 => "10110110",10239 => "11011111",10240 => "11101001",10241 => "10110111",10242 => "01100001",10243 => "01000001",10244 => "00001110",10245 => "11011100",10246 => "00000100",10247 => "01101001",10248 => "00011010",10249 => "00111101",10250 => "10101100",10251 => "01010010",10252 => "11000010",10253 => "11101101",10254 => "11111001",10255 => "11000111",10256 => "00101001",10257 => "01101010",10258 => "01111111",10259 => "00111101",10260 => "00110011",10261 => "01011111",10262 => "10101011",10263 => "11010110",10264 => "11000000",10265 => "00100100",10266 => "11000010",10267 => "00101000",10268 => "01111110",10269 => "10011101",10270 => "10011010",10271 => "00111110",10272 => "10001011",10273 => "00110011",10274 => "11001100",10275 => "00110000",10276 => "11010011",10277 => "11010000",10278 => "00101011",10279 => "00010101",10280 => "10110001",10281 => "11100001",10282 => "00001000",10283 => "00010100",10284 => "01011110",10285 => "01000111",10286 => "01010011",10287 => "11001100",10288 => "11010100",10289 => "00100110",10290 => "01001001",10291 => "10100011",10292 => "11100001",10293 => "01110000",10294 => "11111000",10295 => "01011000",10296 => "00110010",10297 => "10101110",10298 => "11111001",10299 => "01010010",10300 => "00101010",10301 => "11010101",10302 => "00100011",10303 => "00000101",10304 => "10001111",10305 => "11111101",10306 => "01000110",10307 => "01111000",10308 => "00110011",10309 => "10011001",10310 => "01011100",10311 => "00110101",10312 => "00100101",10313 => "00010100",10314 => "01111000",10315 => "00010001",10316 => "01011110",10317 => "00010001",10318 => "01001010",10319 => "00111001",10320 => "11011000",10321 => "01011001",10322 => "11111100",10323 => "00000111",10324 => "10010110",10325 => "00000100",10326 => "01011010",10327 => "00100101",10328 => "01000110",10329 => "01011111",10330 => "01110000",10331 => "00011110",10332 => "01000111",10333 => "10011101",10334 => "01100011",10335 => "11111100",10336 => "01011111",10337 => "11011001",10338 => "01000010",10339 => "01111110",10340 => "11011110",10341 => "11110001",10342 => "01011100",10343 => "11011000",10344 => "01110110",10345 => "01011111",10346 => "00011101",10347 => "10010000",10348 => "00101000",10349 => "00100111",10350 => "11001111",10351 => "01011100",10352 => "00000010",10353 => "00101001",10354 => "00100111",10355 => "11100111",10356 => "10111100",10357 => "10101101",10358 => "01001101",10359 => "00101001",10360 => "01011000",10361 => "01000111",10362 => "10000000",10363 => "10110010",10364 => "11100100",10365 => "00110000",10366 => "10000110",10367 => "01000111",10368 => "01100011",10369 => "00100000",10370 => "00101101",10371 => "01111001",10372 => "01000101",10373 => "11001001",10374 => "11011100",10375 => "00000100",10376 => "11101101",10377 => "00011101",10378 => "11111000",10379 => "11010011",10380 => "01110110",10381 => "10111010",10382 => "00100010",10383 => "00111101",10384 => "10110111",10385 => "11000101",10386 => "10010011",10387 => "00101110",10388 => "00100110",10389 => "10010101",10390 => "10010001",10391 => "00011110",10392 => "10110011",10393 => "10010111",10394 => "00101010",10395 => "10010001",10396 => "01100010",10397 => "11000010",10398 => "10001101",10399 => "00110010",10400 => "01001010",10401 => "00010110",10402 => "01000010",10403 => "10011000",10404 => "11100001",10405 => "01000001",10406 => "00101011",10407 => "01000001",10408 => "01111000",10409 => "10100100",10410 => "11110100",10411 => "10011101",10412 => "10001111",10413 => "10101111",10414 => "10010101",10415 => "10100010",10416 => "10001001",10417 => "11001111",10418 => "11110100",10419 => "11011100",10420 => "10110010",10421 => "00100100",10422 => "01011100",10423 => "10010111",10424 => "11111000",10425 => "01100111",10426 => "01110100",10427 => "01111001",10428 => "11000111",10429 => "10011001",10430 => "11111110",10431 => "10000101",10432 => "11000100",10433 => "00111111",10434 => "10000010",10435 => "10101100",10436 => "11001011",10437 => "10110111",10438 => "00000111",10439 => "11011100",10440 => "11001000",10441 => "10111100",10442 => "11000011",10443 => "10110110",10444 => "00111001",10445 => "10001101",10446 => "10100010",10447 => "01010010",10448 => "01111010",10449 => "00110010",10450 => "00010010",10451 => "01101001",10452 => "01010101",10453 => "00010100",10454 => "11101110",10455 => "00111000",10456 => "10110010",10457 => "01110110",10458 => "00111111",10459 => "01110010",10460 => "10000000",10461 => "11101011",10462 => "01001010",10463 => "00011100",10464 => "01001101",10465 => "11001100",10466 => "10100011",10467 => "10011001",10468 => "10011001",10469 => "01111011",10470 => "00101110",10471 => "01000011",10472 => "01111010",10473 => "01101011",10474 => "10110011",10475 => "00101110",10476 => "00010100",10477 => "01011111",10478 => "01011111",10479 => "01001111",10480 => "10001010",10481 => "10010001",10482 => "10110010",10483 => "10101000",10484 => "00111110",10485 => "11001011",10486 => "10011100",10487 => "01010001",10488 => "00011100",10489 => "01001111",10490 => "00110110",10491 => "10110111",10492 => "10001000",10493 => "00101111",10494 => "10011001",10495 => "01001111",10496 => "11001100",10497 => "11110110",10498 => "10101011",10499 => "10101101",10500 => "10101000",10501 => "01000100",10502 => "11101100",10503 => "01111001",10504 => "10100011",10505 => "01010100",10506 => "10010001",10507 => "01110111",10508 => "10100100",10509 => "00011010",10510 => "00000000",10511 => "11010000",10512 => "11000001",10513 => "01001110",10514 => "10111110",10515 => "00101011",10516 => "01011100",10517 => "10000001",10518 => "10100011",10519 => "10000110",10520 => "10011111",10521 => "11000001",10522 => "01111100",10523 => "10010011",10524 => "10011110",10525 => "10011011",10526 => "10000100",10527 => "10011000",10528 => "10111010",10529 => "11110010",10530 => "00101100",10531 => "11101101",10532 => "00111001",10533 => "11011000",10534 => "01001111",10535 => "11011111",10536 => "10110000",10537 => "00011011",10538 => "10111100",10539 => "11001001",10540 => "01111011",10541 => "10110110",10542 => "00001111",10543 => "11001110",10544 => "10101100",10545 => "00110001",10546 => "01101000",10547 => "10010110",10548 => "10100101",10549 => "10110000",10550 => "10111100",10551 => "01100001",10552 => "01010011",10553 => "11011011",10554 => "11011000",10555 => "10011100",10556 => "11110011",10557 => "01100100",10558 => "01111111",10559 => "00100100",10560 => "00100000",10561 => "10001000",10562 => "00111111",10563 => "10101000",10564 => "01010101",10565 => "01010110",10566 => "01110001",10567 => "11010111",10568 => "10011010",10569 => "00110011",10570 => "10001011",10571 => "10011110",10572 => "10101111",10573 => "00111110",10574 => "01111100",10575 => "01110010",10576 => "11000101",10577 => "11100011",10578 => "11011101",10579 => "01110110",10580 => "01000001",10581 => "01100011",10582 => "10010000",10583 => "00101111",10584 => "10110001",10585 => "00000100",10586 => "10001001",10587 => "00100101",10588 => "01010001",10589 => "01010010",10590 => "11000010",10591 => "00110110",10592 => "00110101",10593 => "10111110",10594 => "11001100",10595 => "11010010",10596 => "11111001",10597 => "01001010",10598 => "10100001",10599 => "00010111",10600 => "01010000",10601 => "11001000",10602 => "01010100",10603 => "10110011",10604 => "10011010",10605 => "01101101",10606 => "11000101",10607 => "10010000",10608 => "10011001",10609 => "00010010",10610 => "11011110",10611 => "00010000",10612 => "00011000",10613 => "00101101",10614 => "11101010",10615 => "10101010",10616 => "11100001",10617 => "11011100",10618 => "01111010",10619 => "01110110",10620 => "11101000",10621 => "10011001",10622 => "11110000",10623 => "01001000",10624 => "10110101",10625 => "11011111",10626 => "01111000",10627 => "01000110",10628 => "00100101",10629 => "00011100",10630 => "00011111",10631 => "01001001",10632 => "01000001",10633 => "11001010",10634 => "01000111",10635 => "00100101",10636 => "00101010",10637 => "10101000",10638 => "10100000",10639 => "00111100",10640 => "11000111",10641 => "11001111",10642 => "00011100",10643 => "11110111",10644 => "10000011",10645 => "11011110",10646 => "10001010",10647 => "00011010",10648 => "00010101",10649 => "01101010",10650 => "11111010",10651 => "00111110",10652 => "10001110",10653 => "11010100",10654 => "11101001",10655 => "00100000",10656 => "00001000",10657 => "00011111",10658 => "11011010",10659 => "10110111",10660 => "00010110",10661 => "11110101",10662 => "01110100",10663 => "10111101",10664 => "11010110",10665 => "11110110",10666 => "10001110",10667 => "00010110",10668 => "00101110",10669 => "10111100",10670 => "10000001",10671 => "10000101",10672 => "11101100",10673 => "00010110",10674 => "10111001",10675 => "10101111",10676 => "00111010",10677 => "01001010",10678 => "10100001",10679 => "00111011",10680 => "11010000",10681 => "01101111",10682 => "01101001",10683 => "10010101",10684 => "00110011",10685 => "01110110",10686 => "01011010",10687 => "01100001",10688 => "11101011",10689 => "00010101",10690 => "10000010",10691 => "01000100",10692 => "10111000",10693 => "01111011",10694 => "10110101",10695 => "10111100",10696 => "11111011",10697 => "00000110",10698 => "00100111",10699 => "01100111",10700 => "00110101",10701 => "11001101",10702 => "00000010",10703 => "10111000",10704 => "00101011",10705 => "01000100",10706 => "11010000",10707 => "01010010",10708 => "10110100",10709 => "10001110",10710 => "00111100",10711 => "00100001",10712 => "00111000",10713 => "00110010",10714 => "11110111",10715 => "00000101",10716 => "10110010",10717 => "01001100",10718 => "10011101",10719 => "11010110",10720 => "01101101",10721 => "10010011",10722 => "11010100",10723 => "00001000",10724 => "00000011",10725 => "01010100",10726 => "10000011",10727 => "10100111",10728 => "00111111",10729 => "10010011",10730 => "10110010",10731 => "01111111",10732 => "01001111",10733 => "10100110",10734 => "11111011",10735 => "00110110",10736 => "10111101",10737 => "11010111",10738 => "11000100",10739 => "10111100",10740 => "11111001",10741 => "10000101",10742 => "00010100",10743 => "10101000",10744 => "10011111",10745 => "01111010",10746 => "10100001",10747 => "11001001",10748 => "10000111",10749 => "01111000",10750 => "01111010",10751 => "10111101",10752 => "01110101",10753 => "01100000",10754 => "11010001",10755 => "11001001",10756 => "01100011",10757 => "00100010",10758 => "10000001",10759 => "10011101",10760 => "01011100",10761 => "00101011",10762 => "11101110",10763 => "10111010",10764 => "11110111",10765 => "01011110",10766 => "01111010",10767 => "11001111",10768 => "11111110",10769 => "10010000",10770 => "00100001",10771 => "00111010",10772 => "01011110",10773 => "01000010",10774 => "01111000",10775 => "11100001",10776 => "01100001",10777 => "10100001",10778 => "00011110",10779 => "11111101",10780 => "11100011",10781 => "10101011",10782 => "10001110",10783 => "00111111",10784 => "11010101",10785 => "01100110",10786 => "10101010",10787 => "11011001",10788 => "11100010",10789 => "11110010",10790 => "10000010",10791 => "11001010",10792 => "11100001",10793 => "01110110",10794 => "10110001",10795 => "01011011",10796 => "10110101",10797 => "01111110",10798 => "01000010",10799 => "10110101",10800 => "10111111",10801 => "01111100",10802 => "11101011",10803 => "11001011",10804 => "01100000",10805 => "01110101",10806 => "10101000",10807 => "10010001",10808 => "11010101",10809 => "10010000",10810 => "01110000",10811 => "01110101",10812 => "01101110",10813 => "10010111",10814 => "01100110",10815 => "11000101",10816 => "11011110",10817 => "01101011",10818 => "00110100",10819 => "01100101",10820 => "01100110",10821 => "10111101",10822 => "10000101",10823 => "00110010",10824 => "10000101",10825 => "00001010",10826 => "00110011",10827 => "00111010",10828 => "01100001",10829 => "01000101",10830 => "01110100",10831 => "10011100",10832 => "10001111",10833 => "01011100",10834 => "00010000",10835 => "00110011",10836 => "10101111",10837 => "10101011",10838 => "10011011",10839 => "01010000",10840 => "01110001",10841 => "11101011",10842 => "10010101",10843 => "00110100",10844 => "00010001",10845 => "01110001",10846 => "10010010",10847 => "10111100",10848 => "01001010",10849 => "01100111",10850 => "01010000",10851 => "11110011",10852 => "10010010",10853 => "00101011",10854 => "10101101",10855 => "00111000",10856 => "01011101",10857 => "01001100",10858 => "11011110",10859 => "11000011",10860 => "00100100",10861 => "11000011",10862 => "10110100",10863 => "10011011",10864 => "01001001",10865 => "11100110",10866 => "00000011",10867 => "00010100",10868 => "01101000",10869 => "01110110",10870 => "00100001",10871 => "11011000",10872 => "10001010",10873 => "11001011",10874 => "11010101",10875 => "01000010",10876 => "00111001",10877 => "01001001",10878 => "00100111",10879 => "01000100",10880 => "11111110",10881 => "00011000",10882 => "00000101",10883 => "10100101",10884 => "11100110",10885 => "11000110",10886 => "11111001",10887 => "01100010",10888 => "01100110",10889 => "10100001",10890 => "00010001",10891 => "10101111",10892 => "00111101",10893 => "10010010",10894 => "00100000",10895 => "01011110",10896 => "11100111",10897 => "11100010",10898 => "00011100",10899 => "10000000",10900 => "10111101",10901 => "00000100",10902 => "10101000",10903 => "10110011",10904 => "10111100",10905 => "01101110",10906 => "00110110",10907 => "01011010",10908 => "10001100",10909 => "01000100",10910 => "11111100",10911 => "11110001",10912 => "10001101",10913 => "01101010",10914 => "00110101",10915 => "11110110",10916 => "00101110",10917 => "11101010",10918 => "01011011",10919 => "11011000",10920 => "01111111",10921 => "11001010",10922 => "10000111",10923 => "10101001",10924 => "10000010",10925 => "11011100",10926 => "00010101",10927 => "01011100",10928 => "11011000",10929 => "11010010",10930 => "00101000",10931 => "01100010",10932 => "10101001",10933 => "10011111",10934 => "00010011",10935 => "11000010",10936 => "01101000",10937 => "10010000",10938 => "01010110",10939 => "01101101",10940 => "00111000",10941 => "01011000",10942 => "00110000",10943 => "00100001",10944 => "10110100",10945 => "00001111",10946 => "01011010",10947 => "10110101",10948 => "01111000",10949 => "00101100",10950 => "11001000",10951 => "10101101",10952 => "11110001",10953 => "10000001",10954 => "11000110",10955 => "00100111",10956 => "01100110",10957 => "11100000",10958 => "00110000",10959 => "11100001",10960 => "11101011",10961 => "00010011",10962 => "11010100",10963 => "10001001",10964 => "00010101",10965 => "01011101",10966 => "00101000",10967 => "00001101",10968 => "10010011",10969 => "10110011",10970 => "00101001",10971 => "10101101",10972 => "10101000",10973 => "00111011",10974 => "11100111",10975 => "00111101",10976 => "01110011",10977 => "10111101",10978 => "01101100",10979 => "01010011",10980 => "01011110",10981 => "01000111",10982 => "11100110",10983 => "00100011",10984 => "11100010",10985 => "11001110",10986 => "10101100",10987 => "00101011",10988 => "01010011",10989 => "00100001",10990 => "01110100",10991 => "01001011",10992 => "01001011",10993 => "01110101",10994 => "01011100",10995 => "10100100",10996 => "10100100",10997 => "00001011",10998 => "10110011",10999 => "10010111",11000 => "00001010",11001 => "01100100",11002 => "01111111",11003 => "10100100",11004 => "01010000",11005 => "00001111",11006 => "01001111",11007 => "11000110",11008 => "00010101",11009 => "00100101",11010 => "11100011",11011 => "11110110",11012 => "11011110",11013 => "10010111",11014 => "11000110",11015 => "00111100",11016 => "10011111",11017 => "01011111",11018 => "00101100",11019 => "10111111",11020 => "10110011",11021 => "11010001",11022 => "11000000",11023 => "10010111",11024 => "11110001",11025 => "00010000",11026 => "00110100",11027 => "00010101",11028 => "00100011",11029 => "01100110",11030 => "11011010",11031 => "10111010",11032 => "01011001",11033 => "11111101",11034 => "11000011",11035 => "11001010",11036 => "11101000",11037 => "01101111",11038 => "11001001",11039 => "01011110",11040 => "10100011",11041 => "11010100",11042 => "10111101",11043 => "10001101",11044 => "10100100",11045 => "00111101",11046 => "10110000",11047 => "00110101",11048 => "11010110",11049 => "00010111",11050 => "10101001",11051 => "00111010",11052 => "00000000",11053 => "00001000",11054 => "00000101",11055 => "00010011",11056 => "11100001",11057 => "00101010",11058 => "00100101",11059 => "00001100",11060 => "01100111",11061 => "01000010",11062 => "00100011",11063 => "11111110",11064 => "10110110",11065 => "01011100",11066 => "00000100",11067 => "00001101",11068 => "11100101",11069 => "11011000",11070 => "01011010",11071 => "01111000",11072 => "10000111",11073 => "10110100",11074 => "01101000",11075 => "10011111",11076 => "00000101",11077 => "01000000",11078 => "10010100",11079 => "01001100",11080 => "01101111",11081 => "01111000",11082 => "00010100",11083 => "10001011",11084 => "11111001",11085 => "10010111",11086 => "11001111",11087 => "00011101",11088 => "10111110",11089 => "01101001",11090 => "10000011",11091 => "10101011",11092 => "01000011",11093 => "00011010",11094 => "01000101",11095 => "00111000",11096 => "11101010",11097 => "11100100",11098 => "00101000",11099 => "00100010",11100 => "01110010",11101 => "11010010",11102 => "11000100",11103 => "00011011",11104 => "01001100",11105 => "01000000",11106 => "11101111",11107 => "11011110",11108 => "00001110",11109 => "00111010",11110 => "11111010",11111 => "01010000",11112 => "11100110",11113 => "10111101",11114 => "01000010",11115 => "10010011",11116 => "11011100",11117 => "00000011",11118 => "01100000",11119 => "11100100",11120 => "10110101",11121 => "11011010",11122 => "11101101",11123 => "11010010",11124 => "01010100",11125 => "01110100",11126 => "10001011",11127 => "01011110",11128 => "00000000",11129 => "10111100",11130 => "11101001",11131 => "00101101",11132 => "01110110",11133 => "00101101",11134 => "00010101",11135 => "01011010",11136 => "00011100",11137 => "00111110",11138 => "11110110",11139 => "11100000",11140 => "00010010",11141 => "11111101",11142 => "01001111",11143 => "00101100",11144 => "01110010",11145 => "00110111",11146 => "01111110",11147 => "00110000",11148 => "11111001",11149 => "01111100",11150 => "11001111",11151 => "10101110",11152 => "11011001",11153 => "01001101",11154 => "01101001",11155 => "11001101",11156 => "00001000",11157 => "10100001",11158 => "10000111",11159 => "01010011",11160 => "11001011",11161 => "10111110",11162 => "11011100",11163 => "01111000",11164 => "10101111",11165 => "10000001",11166 => "11011001",11167 => "11011010",11168 => "11111000",11169 => "11101110",11170 => "01001001",11171 => "10111110",11172 => "11100000",11173 => "00001101",11174 => "00001101",11175 => "11111010",11176 => "00111100",11177 => "10111000",11178 => "10111000",11179 => "01010001",11180 => "01110011",11181 => "01000011",11182 => "10101001",11183 => "11111000",11184 => "10011110",11185 => "10101100",11186 => "01000001",11187 => "10010000",11188 => "11001000",11189 => "11100100",11190 => "11010010",11191 => "10111001",11192 => "01110000",11193 => "10001001",11194 => "00010010",11195 => "00011001",11196 => "11111001",11197 => "10000011",11198 => "10100011",11199 => "10000101",11200 => "10000111",11201 => "01111101",11202 => "01011001",11203 => "10001110",11204 => "00101000",11205 => "01001100",11206 => "01011011",11207 => "10010101",11208 => "11100110",11209 => "00011100",11210 => "10100101",11211 => "00110010",11212 => "11110101",11213 => "10010110",11214 => "01110101",11215 => "00010111",11216 => "00111001",11217 => "10010111",11218 => "11000000",11219 => "11100000",11220 => "10111000",11221 => "00011001",11222 => "11111000",11223 => "00000101",11224 => "11101010",11225 => "01000000",11226 => "01001101",11227 => "11010000",11228 => "11110110",11229 => "01101010",11230 => "01000100",11231 => "10010001",11232 => "00101010",11233 => "01000100",11234 => "10000110",11235 => "01100110",11236 => "10111100",11237 => "00101101",11238 => "00101011",11239 => "11001101",11240 => "00010010",11241 => "10001010",11242 => "10001011",11243 => "01111011",11244 => "10101000",11245 => "10100101",11246 => "10011001",11247 => "10100011",11248 => "00100010",11249 => "10001011",11250 => "11110010",11251 => "10000101",11252 => "01100000",11253 => "00000010",11254 => "00001100",11255 => "00001100",11256 => "11000110",11257 => "01011001",11258 => "00001110",11259 => "01111011",11260 => "01110010",11261 => "11111100",11262 => "11100110",11263 => "11011011",11264 => "10011001",11265 => "10000111",11266 => "00110000",11267 => "01111010",11268 => "01100001",11269 => "11010010",11270 => "01001001",11271 => "00000110",11272 => "11001001",11273 => "11000000",11274 => "01100010",11275 => "01100101",11276 => "11111001",11277 => "00110001",11278 => "00010100",11279 => "00000111",11280 => "00010000",11281 => "00111001",11282 => "11000100",11283 => "01010100",11284 => "10110101",11285 => "00010011",11286 => "10111000",11287 => "00110000",11288 => "11000010",11289 => "00101110",11290 => "10011010",11291 => "00100110",11292 => "11100001",11293 => "10101000",11294 => "00001010",11295 => "01000010",11296 => "11011111",11297 => "01111101",11298 => "00111111",11299 => "10110110",11300 => "00011101",11301 => "11111000",11302 => "01010001",11303 => "00010010",11304 => "01010110",11305 => "10010001",11306 => "00111110",11307 => "00001100",11308 => "10101011",11309 => "00011100",11310 => "11100001",11311 => "11000010",11312 => "10000101",11313 => "00111011",11314 => "01000100",11315 => "11000111",11316 => "10100010",11317 => "01110111",11318 => "01011001",11319 => "11000111",11320 => "01111000",11321 => "01111100",11322 => "01010111",11323 => "11100111",11324 => "00011101",11325 => "00111011",11326 => "11101010",11327 => "00100101",11328 => "10110001",11329 => "10011111",11330 => "00010010",11331 => "00001001",11332 => "01101011",11333 => "10000110",11334 => "00011011",11335 => "00000101",11336 => "11010110",11337 => "10111001",11338 => "11001010",11339 => "01110111",11340 => "01011011",11341 => "11001101",11342 => "10100001",11343 => "10101100",11344 => "10101111",11345 => "11010111",11346 => "00001111",11347 => "00001000",11348 => "01110000",11349 => "11001110",11350 => "01010100",11351 => "01101001",11352 => "11101000",11353 => "11001100",11354 => "01111101",11355 => "10100000",11356 => "01101100",11357 => "01000001",11358 => "10101100",11359 => "00100101",11360 => "11010101",11361 => "01110101",11362 => "01101110",11363 => "10100000",11364 => "01100001",11365 => "01011001",11366 => "00011000",11367 => "10000100",11368 => "00111011",11369 => "00000010",11370 => "00101110",11371 => "01111010",11372 => "11001111",11373 => "01011101",11374 => "00111000",11375 => "11100001",11376 => "11001111",11377 => "00101100",11378 => "10101110",11379 => "10101001",11380 => "00000110",11381 => "11000000",11382 => "00011000",11383 => "11000111",11384 => "10110110",11385 => "01101111",11386 => "10001001",11387 => "01110111",11388 => "10110100",11389 => "10101100",11390 => "00000100",11391 => "00101000",11392 => "11110110",11393 => "10111000",11394 => "11100010",11395 => "10010111",11396 => "00111010",11397 => "11010100",11398 => "01100000",11399 => "11101110",11400 => "00101011",11401 => "01010001",11402 => "01100011",11403 => "00010000",11404 => "00101111",11405 => "10011110",11406 => "00100110",11407 => "10010100",11408 => "01101011",11409 => "01110110",11410 => "10000000",11411 => "10111110",11412 => "10101111",11413 => "00000101",11414 => "00010000",11415 => "00010000",11416 => "00011010",11417 => "11100100",11418 => "01011101",11419 => "01011001",11420 => "01001101",11421 => "11111001",11422 => "00110011",11423 => "10110110",11424 => "11001000",11425 => "10001110",11426 => "01011011",11427 => "00001100",11428 => "11001001",11429 => "11001010",11430 => "00010110",11431 => "01101110",11432 => "11011111",11433 => "01000101",11434 => "00111101",11435 => "10001001",11436 => "01111111",11437 => "11000010",11438 => "01111110",11439 => "10110100",11440 => "01001101",11441 => "00011111",11442 => "01001011",11443 => "10111011",11444 => "11011010",11445 => "10001011",11446 => "10001010",11447 => "00101001",11448 => "01111101",11449 => "01110011",11450 => "10111001",11451 => "10110110",11452 => "00110001",11453 => "00111110",11454 => "01010001",11455 => "11101010",11456 => "10011000",11457 => "10110011",11458 => "10010100",11459 => "00010011",11460 => "01111111",11461 => "00101100",11462 => "00001100",11463 => "00111101",11464 => "01011001",11465 => "01110110",11466 => "11001000",11467 => "00101101",11468 => "11100001",11469 => "11000101",11470 => "01100100",11471 => "11001111",11472 => "00111001",11473 => "01010110",11474 => "01010011",11475 => "11001100",11476 => "11000001",11477 => "00010010",11478 => "11101011",11479 => "00110000",11480 => "00111101",11481 => "01011010",11482 => "10001111",11483 => "10100011",11484 => "11110011",11485 => "01101111",11486 => "01001101",11487 => "10101101",11488 => "10010110",11489 => "10010111",11490 => "01010101",11491 => "11010100",11492 => "01101010",11493 => "01000010",11494 => "00101001",11495 => "00001001",11496 => "11111100",11497 => "01000001",11498 => "11100011",11499 => "11010100",11500 => "01110111",11501 => "01110010",11502 => "10111011",11503 => "01101010",11504 => "01011111",11505 => "00111100",11506 => "01001011",11507 => "00000010",11508 => "11100110",11509 => "00100110",11510 => "10010110",11511 => "01010010",11512 => "11011101",11513 => "11001011",11514 => "00100010",11515 => "11101110",11516 => "00010011",11517 => "11001100",11518 => "11000001",11519 => "00011000",11520 => "01110101",11521 => "01000111",11522 => "10011001",11523 => "00100000",11524 => "11010001",11525 => "00110101",11526 => "00001111",11527 => "01010001",11528 => "11110110",11529 => "01110010",11530 => "11100011",11531 => "01101011",11532 => "10000010",11533 => "10101100",11534 => "10111110",11535 => "00001001",11536 => "11110110",11537 => "11011100",11538 => "10111110",11539 => "01101110",11540 => "00100110",11541 => "01101101",11542 => "01011110",11543 => "10010100",11544 => "11110011",11545 => "11100000",11546 => "10011101",11547 => "00000101",11548 => "10000010",11549 => "10001001",11550 => "11001111",11551 => "10111010",11552 => "00000011",11553 => "10110100",11554 => "00010011",11555 => "01001110",11556 => "10111001",11557 => "01111010",11558 => "10010101",11559 => "10010011",11560 => "01111011",11561 => "00111110",11562 => "11110111",11563 => "10010111",11564 => "01000100",11565 => "01001010",11566 => "10100000",11567 => "11101100",11568 => "00101100",11569 => "10011011",11570 => "01011101",11571 => "11101111",11572 => "11111100",11573 => "01100101",11574 => "11001000",11575 => "10110111",11576 => "11111011",11577 => "00001011",11578 => "11001001",11579 => "11110111",11580 => "10000010",11581 => "01000100",11582 => "10010001",11583 => "11110001",11584 => "11000010",11585 => "00100101",11586 => "01110011",11587 => "11000110",11588 => "10011011",11589 => "11001010",11590 => "00101000",11591 => "01101110",11592 => "11001001",11593 => "11101110",11594 => "11011010",11595 => "01010111",11596 => "11111101",11597 => "10010100",11598 => "10111101",11599 => "00110111",11600 => "00010101",11601 => "11101011",11602 => "00110101",11603 => "10110110",11604 => "10010100",11605 => "01011100",11606 => "00101000",11607 => "11010101",11608 => "00011001",11609 => "00111111",11610 => "01000000",11611 => "10001010",11612 => "01100101",11613 => "00010110",11614 => "01000100",11615 => "01000111",11616 => "11001011",11617 => "01101110",11618 => "00111101",11619 => "10101100",11620 => "01111001",11621 => "11100100",11622 => "00011110",11623 => "00011001",11624 => "01011110",11625 => "11100010",11626 => "10101010",11627 => "00010101",11628 => "10011101",11629 => "01100010",11630 => "00110100",11631 => "00100000",11632 => "11000100",11633 => "00011010",11634 => "11010111",11635 => "11101101",11636 => "01000111",11637 => "10010000",11638 => "11010111",11639 => "01101110",11640 => "10001001",11641 => "10001010",11642 => "00010100",11643 => "01100111",11644 => "11110100",11645 => "11101101",11646 => "10011001",11647 => "01000011",11648 => "11011110",11649 => "00001001",11650 => "10101001",11651 => "00010010",11652 => "11000101",11653 => "00111000",11654 => "10000000",11655 => "10010100",11656 => "00000110",11657 => "10101010",11658 => "01011011",11659 => "11111010",11660 => "11110000",11661 => "01001101",11662 => "00001111",11663 => "00101011",11664 => "00011111",11665 => "10100100",11666 => "11100110",11667 => "00010010",11668 => "01011001",11669 => "11010111",11670 => "11100011",11671 => "10001100",11672 => "10101010",11673 => "01010111",11674 => "10010001",11675 => "11100010",11676 => "10001111",11677 => "10101010",11678 => "01010101",11679 => "10110100",11680 => "10100110",11681 => "11010110",11682 => "00110101",11683 => "00101110",11684 => "00010100",11685 => "11101110",11686 => "00110110",11687 => "01010001",11688 => "00101011",11689 => "11110100",11690 => "00111000",11691 => "01001010",11692 => "00001011",11693 => "00111111",11694 => "00100000",11695 => "01100010",11696 => "11101100",11697 => "11000010",11698 => "10101000",11699 => "11011001",11700 => "00110100",11701 => "00000011",11702 => "11011110",11703 => "00000010",11704 => "10110111",11705 => "10100001",11706 => "11000000",11707 => "10100010",11708 => "10000000",11709 => "11001111",11710 => "10010010",11711 => "00100011",11712 => "00000110",11713 => "11101001",11714 => "01110110",11715 => "01001001",11716 => "10100110",11717 => "10000101",11718 => "10100110",11719 => "00111011",11720 => "01000111",11721 => "10000001",11722 => "01000011",11723 => "11100100",11724 => "10100100",11725 => "01000010",11726 => "00011010",11727 => "00111100",11728 => "01110110",11729 => "10100001",11730 => "01101011",11731 => "00000001",11732 => "10100000",11733 => "11001011",11734 => "00100110",11735 => "11010110",11736 => "10001110",11737 => "01000100",11738 => "11000001",11739 => "10100010",11740 => "10101010",11741 => "10100001",11742 => "11110111",11743 => "11110010",11744 => "00000011",11745 => "00111111",11746 => "01100010",11747 => "01011111",11748 => "11110100",11749 => "01011000",11750 => "11110110",11751 => "10001100",11752 => "10111100",11753 => "11100100",11754 => "10001001",11755 => "00101110",11756 => "11101010",11757 => "00000011",11758 => "11010010",11759 => "10110110",11760 => "00010010",11761 => "01101000",11762 => "01000010",11763 => "01011001",11764 => "00110111",11765 => "01111011",11766 => "01011001",11767 => "00110110",11768 => "11110101",11769 => "00001110",11770 => "10011011",11771 => "00010010",11772 => "11011100",11773 => "11011011",11774 => "10101010",11775 => "11000010",11776 => "00111001",11777 => "10011000",11778 => "10011010",11779 => "11010010",11780 => "00101001",11781 => "11101000",11782 => "10100111",11783 => "10000000",11784 => "01110101",11785 => "01111010",11786 => "00010010",11787 => "01010011",11788 => "00000100",11789 => "11100000",11790 => "01011011",11791 => "01111011",11792 => "01111100",11793 => "11011111",11794 => "00001100",11795 => "00111111",11796 => "01011111",11797 => "01010111",11798 => "10000110",11799 => "01011011",11800 => "00100101",11801 => "11010000",11802 => "00100100",11803 => "11100000",11804 => "00100001",11805 => "10111101",11806 => "11111000",11807 => "10101110",11808 => "00101010",11809 => "01111100",11810 => "00110101",11811 => "11111011",11812 => "00000011",11813 => "00110011",11814 => "11101010",11815 => "10101000",11816 => "10111110",11817 => "10011111",11818 => "00101100",11819 => "01100110",11820 => "10111110",11821 => "11110010",11822 => "10110110",11823 => "10000100",11824 => "00000000",11825 => "10111111",11826 => "10110011",11827 => "10011111",11828 => "01110000",11829 => "01000111",11830 => "11010011",11831 => "01101110",11832 => "10001000",11833 => "01110011",11834 => "10101111",11835 => "10100010",11836 => "11111110",11837 => "11001011",11838 => "11010100",11839 => "11000110",11840 => "11011000",11841 => "10011000",11842 => "01100000",11843 => "01110001",11844 => "11010011",11845 => "01110010",11846 => "11001110",11847 => "10100001",11848 => "10001110",11849 => "10110010",11850 => "10100011",11851 => "00000001",11852 => "10101111",11853 => "01001000",11854 => "00111000",11855 => "10110011",11856 => "11110111",11857 => "10011100",11858 => "00110101",11859 => "10010011",11860 => "00100101",11861 => "11111010",11862 => "01101011",11863 => "01101101",11864 => "11110101",11865 => "10011000",11866 => "01001010",11867 => "01010111",11868 => "01111001",11869 => "00001101",11870 => "10110101",11871 => "11000011",11872 => "11100110",11873 => "01000001",11874 => "11111010",11875 => "00011010",11876 => "00100101",11877 => "10000101",11878 => "10010011",11879 => "01101101",11880 => "11001010",11881 => "00000000",11882 => "11101011",11883 => "10110000",11884 => "10110000",11885 => "01000101",11886 => "10001010",11887 => "11101010",11888 => "11000010",11889 => "01000001",11890 => "10011001",11891 => "10001111",11892 => "01010100",11893 => "01000011",11894 => "01010010",11895 => "00111001",11896 => "11011101",11897 => "00101000",11898 => "01000111",11899 => "11101111",11900 => "01101000",11901 => "01010010",11902 => "11001111",11903 => "10101101",11904 => "11101011",11905 => "01100010",11906 => "10100000",11907 => "00010000",11908 => "10111011",11909 => "00110011",11910 => "10101110",11911 => "11000100",11912 => "00001001",11913 => "10010101",11914 => "10011011",11915 => "10111100",11916 => "10111001",11917 => "00111011",11918 => "10011111",11919 => "11110110",11920 => "00010100",11921 => "10011111",11922 => "00100010",11923 => "10100101",11924 => "11010101",11925 => "10110001",11926 => "10111111",11927 => "00001010",11928 => "00101011",11929 => "00011111",11930 => "10010001",11931 => "10110100",11932 => "01010000",11933 => "10010110",11934 => "11011100",11935 => "00001001",11936 => "11100111",11937 => "11111000",11938 => "10000101",11939 => "00000000",11940 => "01000000",11941 => "00100000",11942 => "11001000",11943 => "10101010",11944 => "11100010",11945 => "00111110",11946 => "10101101",11947 => "11110111",11948 => "01101100",11949 => "10101001",11950 => "11011001",11951 => "01100011",11952 => "01010011",11953 => "00100011",11954 => "10000101",11955 => "01000100",11956 => "01000000",11957 => "11001000",11958 => "01111011",11959 => "00010001",11960 => "10000110",11961 => "10010011",11962 => "01111000",11963 => "01000100",11964 => "00000001",11965 => "00101010",11966 => "11011000",11967 => "11011110",11968 => "10001100",11969 => "10100101",11970 => "00111111",11971 => "11011111",11972 => "00000101",11973 => "01001100",11974 => "10010010",11975 => "01001111",11976 => "11010110",11977 => "10001000",11978 => "00101100",11979 => "00000101",11980 => "01101101",11981 => "10101110",11982 => "00111100",11983 => "01011100",11984 => "00110100",11985 => "01001011",11986 => "11010000",11987 => "00111010",11988 => "11010110",11989 => "00110101",11990 => "11010111",11991 => "00010110",11992 => "11011100",11993 => "11110110",11994 => "11010100",11995 => "00010011",11996 => "00100100",11997 => "01010011",11998 => "00110100",11999 => "11110010",12000 => "00001000",12001 => "11110001",12002 => "00100110",12003 => "00100100",12004 => "11000001",12005 => "11010001",12006 => "11111010",12007 => "00101011",12008 => "11110101",12009 => "01000111",12010 => "10101010",12011 => "10001001",12012 => "11011000",12013 => "01000010",12014 => "01110001",12015 => "01011000",12016 => "10101110",12017 => "01100001",12018 => "11011000",12019 => "00101111",12020 => "00010101",12021 => "10011110",12022 => "00100111",12023 => "00000010",12024 => "11100110",12025 => "10010011",12026 => "10101010",12027 => "10001010",12028 => "11011100",12029 => "00001010",12030 => "00000000",12031 => "01000111",12032 => "01110010",12033 => "01010001",12034 => "01010010",12035 => "11100001",12036 => "10110000",12037 => "10111000",12038 => "11110110",12039 => "10010011",12040 => "11001110",12041 => "10111111",12042 => "01010110",12043 => "00001110",12044 => "11111011",12045 => "01110000",12046 => "11000100",12047 => "10011110",12048 => "11000001",12049 => "00101110",12050 => "01000011",12051 => "01010111",12052 => "10001010",12053 => "00011111",12054 => "00111101",12055 => "11100000",12056 => "10000010",12057 => "10010111",12058 => "11011110",12059 => "00110010",12060 => "10010101",12061 => "00001001",12062 => "01111000",12063 => "10100011",12064 => "00001101",12065 => "00001100",12066 => "01001010",12067 => "11101001",12068 => "00011001",12069 => "11111101",12070 => "10100101",12071 => "10111110",12072 => "11010100",12073 => "01101111",12074 => "01000011",12075 => "01010100",12076 => "11101011",12077 => "01000010",12078 => "00000101",12079 => "11010110",12080 => "01010110",12081 => "01001110",12082 => "00000001",12083 => "01100010",12084 => "11011101",12085 => "00100011",12086 => "01100110",12087 => "01010100",12088 => "10111000",12089 => "11000101",12090 => "11111100",12091 => "01011010",12092 => "10010100",12093 => "10100100",12094 => "11001101",12095 => "11101011",12096 => "00100000",12097 => "01101110",12098 => "01000101",12099 => "01000111",12100 => "00000011",12101 => "11011010",12102 => "00110101",12103 => "01001100",12104 => "10000111",12105 => "01000000",12106 => "00110000",12107 => "11000001",12108 => "01100101",12109 => "10000010",12110 => "10101000",12111 => "11101010",12112 => "11000010",12113 => "11000101",12114 => "10110010",12115 => "10001100",12116 => "10000101",12117 => "11000111",12118 => "01000100",12119 => "10101101",12120 => "11010101",12121 => "10001011",12122 => "10010011",12123 => "10001101",12124 => "00010001",12125 => "00011011",12126 => "01011001",12127 => "01001101",12128 => "00101001",12129 => "10110001",12130 => "10100100",12131 => "10011100",12132 => "11101001",12133 => "00010011",12134 => "11100010",12135 => "01101000",12136 => "01011011",12137 => "11001010",12138 => "01111110",12139 => "00000001",12140 => "01001000",12141 => "11101110",12142 => "11001010",12143 => "10110001",12144 => "01000001",12145 => "10011110",12146 => "00011110",12147 => "10111101",12148 => "11101001",12149 => "00011000",12150 => "10100100",12151 => "10101110",12152 => "01011100",12153 => "10111001",12154 => "10101000",12155 => "10101001",12156 => "00011010",12157 => "00001010",12158 => "01000001",12159 => "10100011",12160 => "01001100",12161 => "11101000",12162 => "10011110",12163 => "01111011",12164 => "00001100",12165 => "01011111",12166 => "01100010",12167 => "11001101",12168 => "11011001",12169 => "11001111",12170 => "01011110",12171 => "10000011",12172 => "00011001",12173 => "11111000",12174 => "00110101",12175 => "01100011",12176 => "11010110",12177 => "11110111",12178 => "10101110",12179 => "11001100",12180 => "00001000",12181 => "10110001",12182 => "01010100",12183 => "11010010",12184 => "10001110",12185 => "01111110",12186 => "10110000",12187 => "01010010",12188 => "11001010",12189 => "11100101",12190 => "11111111",12191 => "00101010",12192 => "11001011",12193 => "11010111",12194 => "01010000",12195 => "00100110",12196 => "01001010",12197 => "00011100",12198 => "11001111",12199 => "11101110",12200 => "10010101",12201 => "11011001",12202 => "11100011",12203 => "11110110",12204 => "00111110",12205 => "01101011",12206 => "11001110",12207 => "11001111",12208 => "10111111",12209 => "11101111",12210 => "01000101",12211 => "00110101",12212 => "00001100",12213 => "11000100",12214 => "11101010",12215 => "00011011",12216 => "10111001",12217 => "10000000",12218 => "00110101",12219 => "00011001",12220 => "01100000",12221 => "10000101",12222 => "01000010",12223 => "01011110",12224 => "00110010",12225 => "11011101",12226 => "10111011",12227 => "01000000",12228 => "10001011",12229 => "00101110",12230 => "10110111",12231 => "00000001",12232 => "01001101",12233 => "00010110",12234 => "10000011",12235 => "10000011",12236 => "10111000",12237 => "11100010",12238 => "00100000",12239 => "00100001",12240 => "11101010",12241 => "00110000",12242 => "00010100",12243 => "01000000",12244 => "01110111",12245 => "00100001",12246 => "00111100",12247 => "00010000",12248 => "00010111",12249 => "01000001",12250 => "11000100",12251 => "11011011",12252 => "01000100",12253 => "11110111",12254 => "10111100",12255 => "11001110",12256 => "00111010",12257 => "11000011",12258 => "00100110",12259 => "00010011",12260 => "00011101",12261 => "11001000",12262 => "11010001",12263 => "00011110",12264 => "00001010",12265 => "10101001",12266 => "01001011",12267 => "01110001",12268 => "00011110",12269 => "01110011",12270 => "11100010",12271 => "01110110",12272 => "11001000",12273 => "00010111",12274 => "01001000",12275 => "10110010",12276 => "00101101",12277 => "10000111",12278 => "11011100",12279 => "01111000",12280 => "11011111",12281 => "00000101",12282 => "01101101",12283 => "01110011",12284 => "10100011",12285 => "00111001",12286 => "00000001",12287 => "00100101",12288 => "01100100",12289 => "10001010",12290 => "11001111",12291 => "10001010",12292 => "10011111",12293 => "11101111",12294 => "10111111",12295 => "10110101",12296 => "10011101",12297 => "11101100",12298 => "11110111",12299 => "11110100",12300 => "01100100",12301 => "01100011",12302 => "00100000",12303 => "01100000",12304 => "11011101",12305 => "11110100",12306 => "01110010",12307 => "01010010",12308 => "11101000",12309 => "01110011",12310 => "10010101",12311 => "11000101",12312 => "01000111",12313 => "11101100",12314 => "10101000",12315 => "00001100",12316 => "11101011",12317 => "00011100",12318 => "00100001",12319 => "00010110",12320 => "00001101",12321 => "11101001",12322 => "01011001",12323 => "00001010",12324 => "00101000",12325 => "11011110",12326 => "10011000",12327 => "00111000",12328 => "01010111",12329 => "11110010",12330 => "10111110",12331 => "10000111",12332 => "00110111",12333 => "11110101",12334 => "10010101",12335 => "01011110",12336 => "00010011",12337 => "10101011",12338 => "11010110",12339 => "01001100",12340 => "00000011",12341 => "10000100",12342 => "01001000",12343 => "01100010",12344 => "00000001",12345 => "11001110",12346 => "11110100",12347 => "01101110",12348 => "01110011",12349 => "10000111",12350 => "00110011",12351 => "11011111",12352 => "11111100",12353 => "11001011",12354 => "00111101",12355 => "01000000",12356 => "00100101",12357 => "10101101",12358 => "01001100",12359 => "10110000",12360 => "00000110",12361 => "00101100",12362 => "01000111",12363 => "11010011",12364 => "10110010",12365 => "00111101",12366 => "10000011",12367 => "01001110",12368 => "10111000",12369 => "11001111",12370 => "10010011",12371 => "00111000",12372 => "00011110",12373 => "10111000",12374 => "10001000",12375 => "01100101",12376 => "10110101",12377 => "10100111",12378 => "00110001",12379 => "00011001",12380 => "01100100",12381 => "11010110",12382 => "10000100",12383 => "00010001",12384 => "11011001",12385 => "01011110",12386 => "10111011",12387 => "00101001",12388 => "01110100",12389 => "10111011",12390 => "00001101",12391 => "00110101",12392 => "01111111",12393 => "11001100",12394 => "01001010",12395 => "00100101",12396 => "11010000",12397 => "00100000",12398 => "00110101",12399 => "00000111",12400 => "00111101",12401 => "01101111",12402 => "00000101",12403 => "01111111",12404 => "10101001",12405 => "01111101",12406 => "11101110",12407 => "00100001",12408 => "11100101",12409 => "10111101",12410 => "11100000",12411 => "00011100",12412 => "00011010",12413 => "01100010",12414 => "01100110",12415 => "10010101",12416 => "01000101",12417 => "01001000",12418 => "11110101",12419 => "10001111",12420 => "01010001",12421 => "10100110",12422 => "00100011",12423 => "00110001",12424 => "10100001",12425 => "01011001",12426 => "10010100",12427 => "10110100",12428 => "01000100",12429 => "01001101",12430 => "10100011",12431 => "01000101",12432 => "00000001",12433 => "10111010",12434 => "00111110",12435 => "11100110",12436 => "10000010",12437 => "00111010",12438 => "10110000",12439 => "10101001",12440 => "00111110",12441 => "01010111",12442 => "11000100",12443 => "10000101",12444 => "00000110",12445 => "01110100",12446 => "00110000",12447 => "00101001",12448 => "11101001",12449 => "00110001",12450 => "01000100",12451 => "01010001",12452 => "00101111",12453 => "11011001",12454 => "01111001",12455 => "00010111",12456 => "00101010",12457 => "01001100",12458 => "00011011",12459 => "00011010",12460 => "00110100",12461 => "00010001",12462 => "00100100",12463 => "01000100",12464 => "10011111",12465 => "01111110",12466 => "11001110",12467 => "10100011",12468 => "01110111",12469 => "00001110",12470 => "10100110",12471 => "01100010",12472 => "01110101",12473 => "00001010",12474 => "10110101",12475 => "11101110",12476 => "01010111",12477 => "00000111",12478 => "01101100",12479 => "01011110",12480 => "11101000",12481 => "10110011",12482 => "01110011",12483 => "10000100",12484 => "01111000",12485 => "00101110",12486 => "01100010",12487 => "10010010",12488 => "11001010",12489 => "10110010",12490 => "11011110",12491 => "11011111",12492 => "00111011",12493 => "01101000",12494 => "01101110",12495 => "11100001",12496 => "11100001",12497 => "01000110",12498 => "00011100",12499 => "11100110",12500 => "10000110",12501 => "11010001",12502 => "01100100",12503 => "10101111",12504 => "10011011",12505 => "10010001",12506 => "01000101",12507 => "10011010",12508 => "00011000",12509 => "00010110",12510 => "00010101",12511 => "10011101",12512 => "00111111",12513 => "11000110",12514 => "10110100",12515 => "11001100",12516 => "10011100",12517 => "11000111",12518 => "10001110",12519 => "11100110",12520 => "10111010",12521 => "01000010",12522 => "00011110",12523 => "10001101",12524 => "01000110",12525 => "00101001",12526 => "00101010",12527 => "00011000",12528 => "11001010",12529 => "00111100",12530 => "01101111",12531 => "10111001",12532 => "00111101",12533 => "10000001",12534 => "01100011",12535 => "00111011",12536 => "10101000",12537 => "01010011",12538 => "11110111",12539 => "10000110",12540 => "11011101",12541 => "11000001",12542 => "11101110",12543 => "01001101",12544 => "10101100",12545 => "00111101",12546 => "01000000",12547 => "10111110",12548 => "10100110",12549 => "00010111",12550 => "11010001",12551 => "11101110",12552 => "00101101",12553 => "11110001",12554 => "11000001",12555 => "00100111",12556 => "11011000",12557 => "01101110",12558 => "11011001",12559 => "00111000",12560 => "00111100",12561 => "10111011",12562 => "11100000",12563 => "00100111",12564 => "10101111",12565 => "10000111",12566 => "00000100",12567 => "10100010",12568 => "10000011",12569 => "00101110",12570 => "10100001",12571 => "10000101",12572 => "10001111",12573 => "11000011",12574 => "11000110",12575 => "01100111",12576 => "10001011",12577 => "11000010",12578 => "11111001",12579 => "11000000",12580 => "10001010",12581 => "01100010",12582 => "10001010",12583 => "10010001",12584 => "10011001",12585 => "01100110",12586 => "01010101",12587 => "00110011",12588 => "10101010",12589 => "10100000",12590 => "10011100",12591 => "11110100",12592 => "00000011",12593 => "01100011",12594 => "10111111",12595 => "00001110",12596 => "00111101",12597 => "01101010",12598 => "01000001",12599 => "01111001",12600 => "10011100",12601 => "00100110",12602 => "01001010",12603 => "01100010",12604 => "00101000",12605 => "11110001",12606 => "11101110",12607 => "00101011",12608 => "11001010",12609 => "11000101",12610 => "10001100",12611 => "10011110",12612 => "10001101",12613 => "11110010",12614 => "11111111",12615 => "00111110",12616 => "00111011",12617 => "00100101",12618 => "00000001",12619 => "00101001",12620 => "10100010",12621 => "10011101",12622 => "00010100",12623 => "00111011",12624 => "10010000",12625 => "10000000",12626 => "00000110",12627 => "10100011",12628 => "11011010",12629 => "00101101",12630 => "11011100",12631 => "01100000",12632 => "00110001",12633 => "10110100",12634 => "01100100",12635 => "00111010",12636 => "01010100",12637 => "10101111",12638 => "11011001",12639 => "11110101",12640 => "11110001",12641 => "11000100",12642 => "10000001",12643 => "11110000",12644 => "01011101",12645 => "10101011",12646 => "10011001",12647 => "00000101",12648 => "00110101",12649 => "01011000",12650 => "11010101",12651 => "01111000",12652 => "11110100",12653 => "01101100",12654 => "01000001",12655 => "00111111",12656 => "01000011",12657 => "11101001",12658 => "10001011",12659 => "00110010",12660 => "10000100",12661 => "10101000",12662 => "00100111",12663 => "11111001",12664 => "10000011",12665 => "11010101",12666 => "10010101",12667 => "11000011",12668 => "01100010",12669 => "00001010",12670 => "10001101",12671 => "01001100",12672 => "10101011",12673 => "10100100",12674 => "01111110",12675 => "00101101",12676 => "10001101",12677 => "11100101",12678 => "11101110",12679 => "01101011",12680 => "00111000",12681 => "01110111",12682 => "10000100",12683 => "00111101",12684 => "01000011",12685 => "11100000",12686 => "11011001",12687 => "01001100",12688 => "01011100",12689 => "11100101",12690 => "10110100",12691 => "11010011",12692 => "11110101",12693 => "01010100",12694 => "10100001",12695 => "01111101",12696 => "11100011",12697 => "10000001",12698 => "00101010",12699 => "11011100",12700 => "10010011",12701 => "00011100",12702 => "00101010",12703 => "00111000",12704 => "11101101",12705 => "01111011",12706 => "01010110",12707 => "01011000",12708 => "11001101",12709 => "11100100",12710 => "01011010",12711 => "11111001",12712 => "10010110",12713 => "10110111",12714 => "11110110",12715 => "11100110",12716 => "10000110",12717 => "10100010",12718 => "00011010",12719 => "11011111",12720 => "00001100",12721 => "10101011",12722 => "00100111",12723 => "11000111",12724 => "01101001",12725 => "00011000",12726 => "01011001",12727 => "10100001",12728 => "10100010",12729 => "00000101",12730 => "11101000",12731 => "11000010",12732 => "01110110",12733 => "00001011",12734 => "11101000",12735 => "00000010",12736 => "00110100",12737 => "11011111",12738 => "10010010",12739 => "11110000",12740 => "11101011",12741 => "10010100",12742 => "10001001",12743 => "01000110",12744 => "10100011",12745 => "00011110",12746 => "10100101",12747 => "11000101",12748 => "00110111",12749 => "10100010",12750 => "01011010",12751 => "00011111",12752 => "10001101",12753 => "11011100",12754 => "10001001",12755 => "01011010",12756 => "10010010",12757 => "01011100",12758 => "11011001",12759 => "11111010",12760 => "01100100",12761 => "00110011",12762 => "01110011",12763 => "01001000",12764 => "10000001",12765 => "10011110",12766 => "01100000",12767 => "00001010",12768 => "10001101",12769 => "10111111",12770 => "00011100",12771 => "01010011",12772 => "01011110",12773 => "01101100",12774 => "00010010",12775 => "10101010",12776 => "00111001",12777 => "01111001",12778 => "11010111",12779 => "01100110",12780 => "01010110",12781 => "10001101",12782 => "00010011",12783 => "11111001",12784 => "10010011",12785 => "10100011",12786 => "01111011",12787 => "10110111",12788 => "00110011",12789 => "11001111",12790 => "10001101",12791 => "11011010",12792 => "10110010",12793 => "00000101",12794 => "00110100",12795 => "01000101",12796 => "01000011",12797 => "00101010",12798 => "01110001",12799 => "01100001",12800 => "01010011",12801 => "01101110",12802 => "00011100",12803 => "11101111",12804 => "00111100",12805 => "11001011",12806 => "00010000",12807 => "10011111",12808 => "01011000",12809 => "00111001",12810 => "01011000",12811 => "00111110",12812 => "00100000",12813 => "00001011",12814 => "10011100",12815 => "01100011",12816 => "10111101",12817 => "11001110",12818 => "01100001",12819 => "01101110",12820 => "10111101",12821 => "11101110",12822 => "01110011",12823 => "10010110",12824 => "10110100",12825 => "10100100",12826 => "10010110",12827 => "10001001",12828 => "01010101",12829 => "01011100",12830 => "00111010",12831 => "01110100",12832 => "01010011",12833 => "01100111",12834 => "00111111",12835 => "01000101",12836 => "10111111",12837 => "10010110",12838 => "00001110",12839 => "10001101",12840 => "10011000",12841 => "00001000",12842 => "10111000",12843 => "10010110",12844 => "10000000",12845 => "01001101",12846 => "11110001",12847 => "00000101",12848 => "01110011",12849 => "01010000",12850 => "01011101",12851 => "11110011",12852 => "00010111",12853 => "01110010",12854 => "10111101",12855 => "11100000",12856 => "00111000",12857 => "01001100",12858 => "00000000",12859 => "11010101",12860 => "00011100",12861 => "01010101",12862 => "01110100",12863 => "10000101",12864 => "01001000",12865 => "10001100",12866 => "11000000",12867 => "10011001",12868 => "10100010",12869 => "01100101",12870 => "01001010",12871 => "11111000",12872 => "11110001",12873 => "01001101",12874 => "11111001",12875 => "10110011",12876 => "01111111",12877 => "01000100",12878 => "11001011",12879 => "01101101",12880 => "00111001",12881 => "00010010",12882 => "11100000",12883 => "00101101",12884 => "10000000",12885 => "00110000",12886 => "00011011",12887 => "01010000",12888 => "11111011",12889 => "00110001",12890 => "11001000",12891 => "00011011",12892 => "00011101",12893 => "01111000",12894 => "01100000",12895 => "00101000",12896 => "11111110",12897 => "11111101",12898 => "11101101",12899 => "10101001",12900 => "01110010",12901 => "01011011",12902 => "01101010",12903 => "10011110",12904 => "01101000",12905 => "10111110",12906 => "00010101",12907 => "01111000",12908 => "11111111",12909 => "11110010",12910 => "10111000",12911 => "01011000",12912 => "11001000",12913 => "10000000",12914 => "01101111",12915 => "01011101",12916 => "10101110",12917 => "01000010",12918 => "01011110",12919 => "00001010",12920 => "00000100",12921 => "00011001",12922 => "11101011",12923 => "00001000",12924 => "01010001",12925 => "00111101",12926 => "01111000",12927 => "01000100",12928 => "11111110",12929 => "10011110",12930 => "10001011",12931 => "10010111",12932 => "11000011",12933 => "00101011",12934 => "01100000",12935 => "10110100",12936 => "00001100",12937 => "10001001",12938 => "11010110",12939 => "01011010",12940 => "11110010",12941 => "11110010",12942 => "00001101",12943 => "11101001",12944 => "11110000",12945 => "11000010",12946 => "01000101",12947 => "00011000",12948 => "11101111",12949 => "01000100",12950 => "10011010",12951 => "11001100",12952 => "01010000",12953 => "01100010",12954 => "10110001",12955 => "01101011",12956 => "00111010",12957 => "01011010",12958 => "11010111",12959 => "10001000",12960 => "01110101",12961 => "11100110",12962 => "00010011",12963 => "00110111",12964 => "11011100",12965 => "00001001",12966 => "01110011",12967 => "10100001",12968 => "01100110",12969 => "01001001",12970 => "01110100",12971 => "10010101",12972 => "01000110",12973 => "10000110",12974 => "01000111",12975 => "01010000",12976 => "11110001",12977 => "11111001",12978 => "11110101",12979 => "00001010",12980 => "00111011",12981 => "00110010",12982 => "10001011",12983 => "11111111",12984 => "01110110",12985 => "11110010",12986 => "10010101",12987 => "01110001",12988 => "11010110",12989 => "10110001",12990 => "11001110",12991 => "10011000",12992 => "10000101",12993 => "01010000",12994 => "11100001",12995 => "00100110",12996 => "11111001",12997 => "01111100",12998 => "01101011",12999 => "10100011",13000 => "01111110",13001 => "01110100",13002 => "00101110",13003 => "00111100",13004 => "11010111",13005 => "11100011",13006 => "01011011",13007 => "00101010",13008 => "01000011",13009 => "00001111",13010 => "10100100",13011 => "11001011",13012 => "01101111",13013 => "01100010",13014 => "10110011",13015 => "10001000",13016 => "11001011",13017 => "00100010",13018 => "01111001",13019 => "00101101",13020 => "11011110",13021 => "11011111",13022 => "10010100",13023 => "11011110",13024 => "00110001",13025 => "10000111",13026 => "00011000",13027 => "11011101",13028 => "10000010",13029 => "00101111",13030 => "01111010",13031 => "00010000",13032 => "11000110",13033 => "10100011",13034 => "00010001",13035 => "00001011",13036 => "00010101",13037 => "10000011",13038 => "00101010",13039 => "00101001",13040 => "01111101",13041 => "01000101",13042 => "11001111",13043 => "11100001",13044 => "01101111",13045 => "00011001",13046 => "11100010",13047 => "01000011",13048 => "01001101",13049 => "11010100",13050 => "11000111",13051 => "01001000",13052 => "11100010",13053 => "10011001",13054 => "11011100",13055 => "10111111",13056 => "00001100",13057 => "11100011",13058 => "11000011",13059 => "11110110",13060 => "10100011",13061 => "10100100",13062 => "11110010",13063 => "10001100",13064 => "01011100",13065 => "11001000",13066 => "11111111",13067 => "10111110",13068 => "00101100",13069 => "00001000",13070 => "01110100",13071 => "00010111",13072 => "10111100",13073 => "11011010",13074 => "11111111",13075 => "01100010",13076 => "11010001",13077 => "11101100",13078 => "11000111",13079 => "10100101",13080 => "00100011",13081 => "10011111",13082 => "01001011",13083 => "11100000",13084 => "10110110",13085 => "00001101",13086 => "11111110",13087 => "01000111",13088 => "10111010",13089 => "10010110",13090 => "01000000",13091 => "00111111",13092 => "10011011",13093 => "11111110",13094 => "00011011",13095 => "10101111",13096 => "01010100",13097 => "01101100",13098 => "11011001",13099 => "01111111",13100 => "11000100",13101 => "01011010",13102 => "01010101",13103 => "00000001",13104 => "00000101",13105 => "01001101",13106 => "11010011",13107 => "11111101",13108 => "01001101",13109 => "11111001",13110 => "10100100",13111 => "11110001",13112 => "01111000",13113 => "11010000",13114 => "00101110",13115 => "00100000",13116 => "10001100",13117 => "11100110",13118 => "11110111",13119 => "10010100",13120 => "11110010",13121 => "11101100",13122 => "11010000",13123 => "01110110",13124 => "01110110",13125 => "00111111",13126 => "11011100",13127 => "10100110",13128 => "10100110",13129 => "01111001",13130 => "01000001",13131 => "00000011",13132 => "00010110",13133 => "11101101",13134 => "11011011",13135 => "01111010",13136 => "00010000",13137 => "10011111",13138 => "11001011",13139 => "00100101",13140 => "01000011",13141 => "00010010",13142 => "10111011",13143 => "10100000",13144 => "00000001",13145 => "10001101",13146 => "11111100",13147 => "01011011",13148 => "00010010",13149 => "01011111",13150 => "10010100",13151 => "01011000",13152 => "00000011",13153 => "01111000",13154 => "01110111",13155 => "11111001",13156 => "01101001",13157 => "01000110",13158 => "00000010",13159 => "01001101",13160 => "10011110",13161 => "00000000",13162 => "10001110",13163 => "00110001",13164 => "00010111",13165 => "10001001",13166 => "11000110",13167 => "00001000",13168 => "11010111",13169 => "10110001",13170 => "01011110",13171 => "10101111",13172 => "01001001",13173 => "11101000",13174 => "10101010",13175 => "11110101",13176 => "10111001",13177 => "00111100",13178 => "01000100",13179 => "01001101",13180 => "01001100",13181 => "00111001",13182 => "10110001",13183 => "01111110",13184 => "11011100",13185 => "01100110",13186 => "11101001",13187 => "01000101",13188 => "11101000",13189 => "01001001",13190 => "01000010",13191 => "00111000",13192 => "00111101",13193 => "11101010",13194 => "00010010",13195 => "01010110",13196 => "01011000",13197 => "10101101",13198 => "11000000",13199 => "11101001",13200 => "11001100",13201 => "00010110",13202 => "11110001",13203 => "01001101",13204 => "00000000",13205 => "11111011",13206 => "00001011",13207 => "01111110",13208 => "10000100",13209 => "01001111",13210 => "00001101",13211 => "10010001",13212 => "10000011",13213 => "01111000",13214 => "01110111",13215 => "11010001",13216 => "01011000",13217 => "10000110",13218 => "01111101",13219 => "10110110",13220 => "01011101",13221 => "10011101",13222 => "01000110",13223 => "11100010",13224 => "11000000",13225 => "10111010",13226 => "11111111",13227 => "00001100",13228 => "11000110",13229 => "10001111",13230 => "01011001",13231 => "01110110",13232 => "01111011",13233 => "01111100",13234 => "01111111",13235 => "10110100",13236 => "00000101",13237 => "01100100",13238 => "10000010",13239 => "10101000",13240 => "11110100",13241 => "10011011",13242 => "11101111",13243 => "11111101",13244 => "00111101",13245 => "10101001",13246 => "01001000",13247 => "10100000",13248 => "01001010",13249 => "10001000",13250 => "01011011",13251 => "00111100",13252 => "11010001",13253 => "01101000",13254 => "10100101",13255 => "01011101",13256 => "10101110",13257 => "00011100",13258 => "10111001",13259 => "10010010",13260 => "01100101",13261 => "10110011",13262 => "10010110",13263 => "00111011",13264 => "10110101",13265 => "00000111",13266 => "00110010",13267 => "11000111",13268 => "10111111",13269 => "01110111",13270 => "01011111",13271 => "00111100",13272 => "01110101",13273 => "11111001",13274 => "11111110",13275 => "00001001",13276 => "00000001",13277 => "01111111",13278 => "01101001",13279 => "01100001",13280 => "10101110",13281 => "00000101",13282 => "01001100",13283 => "10101101",13284 => "01110101",13285 => "11010110",13286 => "11101000",13287 => "00110001",13288 => "11001001",13289 => "10110001",13290 => "00100011",13291 => "11110011",13292 => "01111011",13293 => "11100101",13294 => "11000100",13295 => "01011001",13296 => "01011011",13297 => "01101001",13298 => "01011011",13299 => "00001001",13300 => "10011100",13301 => "01010110",13302 => "10101001",13303 => "00111000",13304 => "10010110",13305 => "01000100",13306 => "11001110",13307 => "11010110",13308 => "01001111",13309 => "00000010",13310 => "10011101",13311 => "11111110",13312 => "11000110",13313 => "01101101",13314 => "11111001",13315 => "01111100",13316 => "01010010",13317 => "11010110",13318 => "01100001",13319 => "00100101",13320 => "01010111",13321 => "11101111",13322 => "11011101",13323 => "00000011",13324 => "01100101",13325 => "00111000",13326 => "11000000",13327 => "10111010",13328 => "01101010",13329 => "10101000",13330 => "01001000",13331 => "10010001",13332 => "10011110",13333 => "00100000",13334 => "01111011",13335 => "10100000",13336 => "10000010",13337 => "00111100",13338 => "11111110",13339 => "10101011",13340 => "01110010",13341 => "00101010",13342 => "00010001",13343 => "10101001",13344 => "10111011",13345 => "10010011",13346 => "00011111",13347 => "10010100",13348 => "01000000",13349 => "01001111",13350 => "10101111",13351 => "11110001",13352 => "01011000",13353 => "00010111",13354 => "00001101",13355 => "01010010",13356 => "00111011",13357 => "01011100",13358 => "10110010",13359 => "11011101",13360 => "01100010",13361 => "10111010",13362 => "00011110",13363 => "00101111",13364 => "01110011",13365 => "01011000",13366 => "00101011",13367 => "11010110",13368 => "11111000",13369 => "10101111",13370 => "00011101",13371 => "11100110",13372 => "10010011",13373 => "00001110",13374 => "11010111",13375 => "00110011",13376 => "00111101",13377 => "10110011",13378 => "10100111",13379 => "10111111",13380 => "10010000",13381 => "01111100",13382 => "10010000",13383 => "10101100",13384 => "10000010",13385 => "01000001",13386 => "10100010",13387 => "10100011",13388 => "00010011",13389 => "00010010",13390 => "11010000",13391 => "11110000",13392 => "00010000",13393 => "00010000",13394 => "10111011",13395 => "11010011",13396 => "10101101",13397 => "00110110",13398 => "00110111",13399 => "00110011",13400 => "00011110",13401 => "01100101",13402 => "01010100",13403 => "10100001",13404 => "01111101",13405 => "00001010",13406 => "10011011",13407 => "00001111",13408 => "00110000",13409 => "11111110",13410 => "00111000",13411 => "01111001",13412 => "10011110",13413 => "11001101",13414 => "01100000",13415 => "01110100",13416 => "01110010",13417 => "11001010",13418 => "10111101",13419 => "10100010",13420 => "11001001",13421 => "01101011",13422 => "01111101",13423 => "00100110",13424 => "11101111",13425 => "01111011",13426 => "11110100",13427 => "10001010",13428 => "10111101",13429 => "11110110",13430 => "00000001",13431 => "01111010",13432 => "11001001",13433 => "11101110",13434 => "11001111",13435 => "00010100",13436 => "01000000",13437 => "01100011",13438 => "01001110",13439 => "11000110",13440 => "00000000",13441 => "10110111",13442 => "10001011",13443 => "01000011",13444 => "11100111",13445 => "11100010",13446 => "00000001",13447 => "11000101",13448 => "11000110",13449 => "10001000",13450 => "01011110",13451 => "11101110",13452 => "11100111",13453 => "01001101",13454 => "11110110",13455 => "00010100",13456 => "10011110",13457 => "10100000",13458 => "01000001",13459 => "00000100",13460 => "00000011",13461 => "01110010",13462 => "01001101",13463 => "00111001",13464 => "00011000",13465 => "11010110",13466 => "00010111",13467 => "01001100",13468 => "10100011",13469 => "00110110",13470 => "01010101",13471 => "10101011",13472 => "11111100",13473 => "00111001",13474 => "10111001",13475 => "00001101",13476 => "01010000",13477 => "01100011",13478 => "00100001",13479 => "11111010",13480 => "00010010",13481 => "11101010",13482 => "10000000",13483 => "10001010",13484 => "10101010",13485 => "00000100",13486 => "00101100",13487 => "01000101",13488 => "00110011",13489 => "11111001",13490 => "00111111",13491 => "01011101",13492 => "10000011",13493 => "10000001",13494 => "10101000",13495 => "00011000",13496 => "11000010",13497 => "10111000",13498 => "10000001",13499 => "01100001",13500 => "10111000",13501 => "00111011",13502 => "00011001",13503 => "00110001",13504 => "01010101",13505 => "01011010",13506 => "00001001",13507 => "11000011",13508 => "10011101",13509 => "11011010",13510 => "11110101",13511 => "01000011",13512 => "10001111",13513 => "11010110",13514 => "10101010",13515 => "00101100",13516 => "00010110",13517 => "11001101",13518 => "00001101",13519 => "11110111",13520 => "11110000",13521 => "11000000",13522 => "10100010",13523 => "11100001",13524 => "00000010",13525 => "11111111",13526 => "00001110",13527 => "00101000",13528 => "00111001",13529 => "01000110",13530 => "10110110",13531 => "10111000",13532 => "11010110",13533 => "10010001",13534 => "11010111",13535 => "00100000",13536 => "10100100",13537 => "01011011",13538 => "01110100",13539 => "01001000",13540 => "11110010",13541 => "11111010",13542 => "11000001",13543 => "10111110",13544 => "11100010",13545 => "10111101",13546 => "00001011",13547 => "10101101",13548 => "11001110",13549 => "01110101",13550 => "10110100",13551 => "01101000",13552 => "11100100",13553 => "11111000",13554 => "10001110",13555 => "10010110",13556 => "01100110",13557 => "11101100",13558 => "01010001",13559 => "10111101",13560 => "11111100",13561 => "00110000",13562 => "10111110",13563 => "01000001",13564 => "11100101",13565 => "01001001",13566 => "01010100",13567 => "00011100",13568 => "10111101",13569 => "01110011",13570 => "10010010",13571 => "01000111",13572 => "11011101",13573 => "10111000",13574 => "00011001",13575 => "01011001",13576 => "10001001",13577 => "10110110",13578 => "00110011",13579 => "00000111",13580 => "00011100",13581 => "10101111",13582 => "10001001",13583 => "01101010",13584 => "00000110",13585 => "00111110",13586 => "11011011",13587 => "10100100",13588 => "01010011",13589 => "11010010",13590 => "00001110",13591 => "10100000",13592 => "00101001",13593 => "10010100",13594 => "10111101",13595 => "10100001",13596 => "11110011",13597 => "11001110",13598 => "10100011",13599 => "00010001",13600 => "00101010",13601 => "00100100",13602 => "11010111",13603 => "11010110",13604 => "01110001",13605 => "10101000",13606 => "11011111",13607 => "00000110",13608 => "01000011",13609 => "10110010",13610 => "11011011",13611 => "10000011",13612 => "10011100",13613 => "00100111",13614 => "11111100",13615 => "11011110",13616 => "10000110",13617 => "10000101",13618 => "11101010",13619 => "10011000",13620 => "11111010",13621 => "01111111",13622 => "00100011",13623 => "00111001",13624 => "01100100",13625 => "11010101",13626 => "10100000",13627 => "11011000",13628 => "00000101",13629 => "10110001",13630 => "11101001",13631 => "10010111",13632 => "00011110",13633 => "00001101",13634 => "00101111",13635 => "00001010",13636 => "11010111",13637 => "11011100",13638 => "00100001",13639 => "10001000",13640 => "01010011",13641 => "10101010",13642 => "10010010",13643 => "11100011",13644 => "00101010",13645 => "00101011",13646 => "01110000",13647 => "00110111",13648 => "11000010",13649 => "11011101",13650 => "10011100",13651 => "10111000",13652 => "10100011",13653 => "01000000",13654 => "11010100",13655 => "10010011",13656 => "11100111",13657 => "01011011",13658 => "00000011",13659 => "10001010",13660 => "11001011",13661 => "11111101",13662 => "00001100",13663 => "10110101",13664 => "00100100",13665 => "00110101",13666 => "01100010",13667 => "01101101",13668 => "01010110",13669 => "00001000",13670 => "00001100",13671 => "00000011",13672 => "01010010",13673 => "11001100",13674 => "11011001",13675 => "00001000",13676 => "11100001",13677 => "11100100",13678 => "11010111",13679 => "00100001",13680 => "00100001",13681 => "01110000",13682 => "01010110",13683 => "00100011",13684 => "00010010",13685 => "11111011",13686 => "01100001",13687 => "11100001",13688 => "00110001",13689 => "10011110",13690 => "11101010",13691 => "10101001",13692 => "11000100",13693 => "10101111",13694 => "01001111",13695 => "01000111",13696 => "11011000",13697 => "01010010",13698 => "11111100",13699 => "00001000",13700 => "11010010",13701 => "10010100",13702 => "01111111",13703 => "10111000",13704 => "11110001",13705 => "11001010",13706 => "00111101",13707 => "11011001",13708 => "10111010",13709 => "00110010",13710 => "10001101",13711 => "10110110",13712 => "00110101",13713 => "11100000",13714 => "00111011",13715 => "01101011",13716 => "01101100",13717 => "01001101",13718 => "01100101",13719 => "00000101",13720 => "10110010",13721 => "11111100",13722 => "00111001",13723 => "10001110",13724 => "10000011",13725 => "10011101",13726 => "00010110",13727 => "11110101",13728 => "10100100",13729 => "11010010",13730 => "10100101",13731 => "01010111",13732 => "10001001",13733 => "00000010",13734 => "00011100",13735 => "10101100",13736 => "01110110",13737 => "00010000",13738 => "10011101",13739 => "00000111",13740 => "11010010",13741 => "11111001",13742 => "11000110",13743 => "10001001",13744 => "01011010",13745 => "01001101",13746 => "00101100",13747 => "00011111",13748 => "11011111",13749 => "01011110",13750 => "10111110",13751 => "01111001",13752 => "00110001",13753 => "00110010",13754 => "00110011",13755 => "10001101",13756 => "10100101",13757 => "01101111",13758 => "10101000",13759 => "00001011",13760 => "00010001",13761 => "01011001",13762 => "00000010",13763 => "01110111",13764 => "00000000",13765 => "10110111",13766 => "00011110",13767 => "10111101",13768 => "00101011",13769 => "01100100",13770 => "01000000",13771 => "11110100",13772 => "01111000",13773 => "00111011",13774 => "00100110",13775 => "01011111",13776 => "11110010",13777 => "10000100",13778 => "11011110",13779 => "00011100",13780 => "01111100",13781 => "10000000",13782 => "01010011",13783 => "11110100",13784 => "11000111",13785 => "11011010",13786 => "01110000",13787 => "11001100",13788 => "10001011",13789 => "11110011",13790 => "10010001",13791 => "01100000",13792 => "11000001",13793 => "00011111",13794 => "00001110",13795 => "00010010",13796 => "11101110",13797 => "00010100",13798 => "01111110",13799 => "00100110",13800 => "10110100",13801 => "10101001",13802 => "01010110",13803 => "01011011",13804 => "01110011",13805 => "00111010",13806 => "00111101",13807 => "10101000",13808 => "11110111",13809 => "00111101",13810 => "11010010",13811 => "10101011",13812 => "01001001",13813 => "01111000",13814 => "11101010",13815 => "01100000",13816 => "11010001",13817 => "11110100",13818 => "01110111",13819 => "11010100",13820 => "01100101",13821 => "10111011",13822 => "01000010",13823 => "10100011",13824 => "10111101",13825 => "10110100",13826 => "11010111",13827 => "10110011",13828 => "10110100",13829 => "01011010",13830 => "01101011",13831 => "00001010",13832 => "10101100",13833 => "00111101",13834 => "00001000",13835 => "00000101",13836 => "10111010",13837 => "10111000",13838 => "00101111",13839 => "00101111",13840 => "11011001",13841 => "10101001",13842 => "01010001",13843 => "11110101",13844 => "01100110",13845 => "10100001",13846 => "00000000",13847 => "10101111",13848 => "01001010",13849 => "11001010",13850 => "10010010",13851 => "10010101",13852 => "11001110",13853 => "00110111",13854 => "10000010",13855 => "10011101",13856 => "10001110",13857 => "10010011",13858 => "00111011",13859 => "11110000",13860 => "00101011",13861 => "00111001",13862 => "01100100",13863 => "10011100",13864 => "11111001",13865 => "10111000",13866 => "10111001",13867 => "00110100",13868 => "01101000",13869 => "10011010",13870 => "11010111",13871 => "11101010",13872 => "10110110",13873 => "01110100",13874 => "10100100",13875 => "01001011",13876 => "01001110",13877 => "01110110",13878 => "10001100",13879 => "01001001",13880 => "01001000",13881 => "10011100",13882 => "01100011",13883 => "10001000",13884 => "00000111",13885 => "01101100",13886 => "00111010",13887 => "00100000",13888 => "01010010",13889 => "01010101",13890 => "00011100",13891 => "01001010",13892 => "11110011",13893 => "01110100",13894 => "10101110",13895 => "10011110",13896 => "00000000",13897 => "00100001",13898 => "10111000",13899 => "10111111",13900 => "10010111",13901 => "10010001",13902 => "00011000",13903 => "00000101",13904 => "00001111",13905 => "11001010",13906 => "11100000",13907 => "01110001",13908 => "01000111",13909 => "11111101",13910 => "00111001",13911 => "00110111",13912 => "11010100",13913 => "11011101",13914 => "01011110",13915 => "01011101",13916 => "01000000",13917 => "01100110",13918 => "01111011",13919 => "01011110",13920 => "01110000",13921 => "00000110",13922 => "01011000",13923 => "00001001",13924 => "11011000",13925 => "11011101",13926 => "11101010",13927 => "10010000",13928 => "10100001",13929 => "10001100",13930 => "11011101",13931 => "11011011",13932 => "00111001",13933 => "10100011",13934 => "01100100",13935 => "10011000",13936 => "01110110",13937 => "01110100",13938 => "00101101",13939 => "01011001",13940 => "01010001",13941 => "11101111",13942 => "00100001",13943 => "00000010",13944 => "10001001",13945 => "00111100",13946 => "11000110",13947 => "11000011",13948 => "11111011",13949 => "11011011",13950 => "00111010",13951 => "01000110",13952 => "01111101",13953 => "10001100",13954 => "01101000",13955 => "10100101",13956 => "01010000",13957 => "01100000",13958 => "01011000",13959 => "11000000",13960 => "00110010",13961 => "01110000",13962 => "01000000",13963 => "00011110",13964 => "11111101",13965 => "11110001",13966 => "01010101",13967 => "01100110",13968 => "11111100",13969 => "01110110",13970 => "11101011",13971 => "11000101",13972 => "00011101",13973 => "00100011",13974 => "00101001",13975 => "11101110",13976 => "10111111",13977 => "00101111",13978 => "10101110",13979 => "00111110",13980 => "10001000",13981 => "00011010",13982 => "01101000",13983 => "11000110",13984 => "11101010",13985 => "00111000",13986 => "00111001",13987 => "01111011",13988 => "00100101",13989 => "10011011",13990 => "11110010",13991 => "01110000",13992 => "00111100",13993 => "01000100",13994 => "01011010",13995 => "00101110",13996 => "10111110",13997 => "00001000",13998 => "01110100",13999 => "00110010",14000 => "11100011",14001 => "01000010",14002 => "10101011",14003 => "11001111",14004 => "11001100",14005 => "01011011",14006 => "00110000",14007 => "10100111",14008 => "01010100",14009 => "10110010",14010 => "10110011",14011 => "11011111",14012 => "10011010",14013 => "00011100",14014 => "10000111",14015 => "10011101",14016 => "00011010",14017 => "11111011",14018 => "11011111",14019 => "10001111",14020 => "10011011",14021 => "01110001",14022 => "00100101",14023 => "01001011",14024 => "10110010",14025 => "10001100",14026 => "11010001",14027 => "11000000",14028 => "11101001",14029 => "11110110",14030 => "10101101",14031 => "00101111",14032 => "00010111",14033 => "10001101",14034 => "00010101",14035 => "11110000",14036 => "00000101",14037 => "00100010",14038 => "11000001",14039 => "11101001",14040 => "11011010",14041 => "10001000",14042 => "01001011",14043 => "01111010",14044 => "11100001",14045 => "01111001",14046 => "10011111",14047 => "11101010",14048 => "10100011",14049 => "01000110",14050 => "00111010",14051 => "11010100",14052 => "01110010",14053 => "01011001",14054 => "00110001",14055 => "00000001",14056 => "01100001",14057 => "10100111",14058 => "10011010",14059 => "11111001",14060 => "01100011",14061 => "10100011",14062 => "01111011",14063 => "11111011",14064 => "10011001",14065 => "00100110",14066 => "00000010",14067 => "10011000",14068 => "01111000",14069 => "11100110",14070 => "11101110",14071 => "01111001",14072 => "11010011",14073 => "10111100",14074 => "11001111",14075 => "01010110",14076 => "00000001",14077 => "11111010",14078 => "11010011",14079 => "10100100",14080 => "01101110",14081 => "00011010",14082 => "00000111",14083 => "11000000",14084 => "00011001",14085 => "00101101",14086 => "00010111",14087 => "01000100",14088 => "01101010",14089 => "00000100",14090 => "10101100",14091 => "00110101",14092 => "11000110",14093 => "10011011",14094 => "01000111",14095 => "01111111",14096 => "00110110",14097 => "01001110",14098 => "10010111",14099 => "00000001",14100 => "00110111",14101 => "01101110",14102 => "11111001",14103 => "10100011",14104 => "11010110",14105 => "01110010",14106 => "11101000",14107 => "11110110",14108 => "01001001",14109 => "01110100",14110 => "01111011",14111 => "10110111",14112 => "11001100",14113 => "00010001",14114 => "11111111",14115 => "10001100",14116 => "00111010",14117 => "11101000",14118 => "01100110",14119 => "10001001",14120 => "11111100",14121 => "01110011",14122 => "01011010",14123 => "11100110",14124 => "11000011",14125 => "11111100",14126 => "11101101",14127 => "11111100",14128 => "00001110",14129 => "00011000",14130 => "11110111",14131 => "00010000",14132 => "00100100",14133 => "01111111",14134 => "01111101",14135 => "11000101",14136 => "00110001",14137 => "11011110",14138 => "00011100",14139 => "01011101",14140 => "11110000",14141 => "10111101",14142 => "00011000",14143 => "11101111",14144 => "10100110",14145 => "01011100",14146 => "10000011",14147 => "01100000",14148 => "11111111",14149 => "11011110",14150 => "10110101",14151 => "10110100",14152 => "11000010",14153 => "00110100",14154 => "11000000",14155 => "11001011",14156 => "10011000",14157 => "01111111",14158 => "01111100",14159 => "00000000",14160 => "01110100",14161 => "11101011",14162 => "01101010",14163 => "10011101",14164 => "01101110",14165 => "01000111",14166 => "00010010",14167 => "01011111",14168 => "00111000",14169 => "11101011",14170 => "11001011",14171 => "00010100",14172 => "00000111",14173 => "00110000",14174 => "10101101",14175 => "01011111",14176 => "10100111",14177 => "10011001",14178 => "10110010",14179 => "11111101",14180 => "01100011",14181 => "11111010",14182 => "10000010",14183 => "11011001",14184 => "11001001",14185 => "11011100",14186 => "11101011",14187 => "10001100",14188 => "00100010",14189 => "01100000",14190 => "01111100",14191 => "11000010",14192 => "10001111",14193 => "01110000",14194 => "01111111",14195 => "01101010",14196 => "11010000",14197 => "10011010",14198 => "10110010",14199 => "10001101",14200 => "00101011",14201 => "10001111",14202 => "01110101",14203 => "11010111",14204 => "00001101",14205 => "11011000",14206 => "10111111",14207 => "11001010",14208 => "00010010",14209 => "10000011",14210 => "00100111",14211 => "10010001",14212 => "01001110",14213 => "00000110",14214 => "11011010",14215 => "00010111",14216 => "11101001",14217 => "11000111",14218 => "11000010",14219 => "11101100",14220 => "10010001",14221 => "01011010",14222 => "01101010",14223 => "01000110",14224 => "10111110",14225 => "01100101",14226 => "00000111",14227 => "01111010",14228 => "00101101",14229 => "00111010",14230 => "11000001",14231 => "00100100",14232 => "10100110",14233 => "00110001",14234 => "11000001",14235 => "11000110",14236 => "00011100",14237 => "00110011",14238 => "11100011",14239 => "11010101",14240 => "11100100",14241 => "11111110",14242 => "00010111",14243 => "11110010",14244 => "10110000",14245 => "11100011",14246 => "00001100",14247 => "00001100",14248 => "01100110",14249 => "10011100",14250 => "00000010",14251 => "01110100",14252 => "00100011",14253 => "10101010",14254 => "11100100",14255 => "01100101",14256 => "10110111",14257 => "00100110",14258 => "00100001",14259 => "01000001",14260 => "10001001",14261 => "01111011",14262 => "01100110",14263 => "10011111",14264 => "11011010",14265 => "01100000",14266 => "00100011",14267 => "01010011",14268 => "11001000",14269 => "00100101",14270 => "01011010",14271 => "10110110",14272 => "01000100",14273 => "01110010",14274 => "01011101",14275 => "00101100",14276 => "00101010",14277 => "10101111",14278 => "10001101",14279 => "10011001",14280 => "11000101",14281 => "11100010",14282 => "11110110",14283 => "00111101",14284 => "11100100",14285 => "00101000",14286 => "10011110",14287 => "10011010",14288 => "10100001",14289 => "01000000",14290 => "00001000",14291 => "10110111",14292 => "00010010",14293 => "11001010",14294 => "00001000",14295 => "10110001",14296 => "10100001",14297 => "10111111",14298 => "11100111",14299 => "00111110",14300 => "11001001",14301 => "01101101",14302 => "01110011",14303 => "01110010",14304 => "00011101",14305 => "11001101",14306 => "11010100",14307 => "10011111",14308 => "11000101",14309 => "11100111",14310 => "00000000",14311 => "01000000",14312 => "01010011",14313 => "11101110",14314 => "01110111",14315 => "10100000",14316 => "00001011",14317 => "11011000",14318 => "01010100",14319 => "10010001",14320 => "10000011",14321 => "00000001",14322 => "11101101",14323 => "00011101",14324 => "01001100",14325 => "11010010",14326 => "11111001",14327 => "00101010",14328 => "11111000",14329 => "01010001",14330 => "00011110",14331 => "01111011",14332 => "01011110",14333 => "11001011",14334 => "00010001",14335 => "01101001",14336 => "01101111",14337 => "00001101",14338 => "01011001",14339 => "01100010",14340 => "11011100",14341 => "10100110",14342 => "10010101",14343 => "01110110",14344 => "11100001",14345 => "01111101",14346 => "11000110",14347 => "11111100",14348 => "00111011",14349 => "01111101",14350 => "01111110",14351 => "01111100",14352 => "10011011",14353 => "10101000",14354 => "11001101",14355 => "11010111",14356 => "10101110",14357 => "11110100",14358 => "10101001",14359 => "10111001",14360 => "11010101",14361 => "11001011",14362 => "01011011",14363 => "01000110",14364 => "10000001",14365 => "00110011",14366 => "00001110",14367 => "11101000",14368 => "11010100",14369 => "10110110",14370 => "00000001",14371 => "11001100",14372 => "11010011",14373 => "00001011",14374 => "00111111",14375 => "01011101",14376 => "11000010",14377 => "01011111",14378 => "00011001",14379 => "10010101",14380 => "00100000",14381 => "10110010",14382 => "01100000",14383 => "01110110",14384 => "10000000",14385 => "10110111",14386 => "01110010",14387 => "00001010",14388 => "10100001",14389 => "01000101",14390 => "01001110",14391 => "11101100",14392 => "00011001",14393 => "10001110",14394 => "10110011",14395 => "00011000",14396 => "11101000",14397 => "01000100",14398 => "00010011",14399 => "00000101",14400 => "01110100",14401 => "01111000",14402 => "01111110",14403 => "11010101",14404 => "01011000",14405 => "01010010",14406 => "10011110",14407 => "00000010",14408 => "01011111",14409 => "11110011",14410 => "10001010",14411 => "01010010",14412 => "00010010",14413 => "11100110",14414 => "10001101",14415 => "01111001",14416 => "11010011",14417 => "10010100",14418 => "00111110",14419 => "11100111",14420 => "11001010",14421 => "10110100",14422 => "00011110",14423 => "11011011",14424 => "10000101",14425 => "10101001",14426 => "11011000",14427 => "00101101",14428 => "11010111",14429 => "10111110",14430 => "11001111",14431 => "10010010",14432 => "01101101",14433 => "00111111",14434 => "00010101",14435 => "10001111",14436 => "01001110",14437 => "10001001",14438 => "01011001",14439 => "11010110",14440 => "10011010",14441 => "11010111",14442 => "11011100",14443 => "10101010",14444 => "10111011",14445 => "10000100",14446 => "11001110",14447 => "00110001",14448 => "00011010",14449 => "00110011",14450 => "11011110",14451 => "10010100",14452 => "00111101",14453 => "01000011",14454 => "00110010",14455 => "00111011",14456 => "11111110",14457 => "10010000",14458 => "10000101",14459 => "01111010",14460 => "01010011",14461 => "11000100",14462 => "10110010",14463 => "01110011",14464 => "00101100",14465 => "00110101",14466 => "11100110",14467 => "10001000",14468 => "00001110",14469 => "01000001",14470 => "11000111",14471 => "00101011",14472 => "11000100",14473 => "01001110",14474 => "10101010",14475 => "01110111",14476 => "10110001",14477 => "00000101",14478 => "01001111",14479 => "10110001",14480 => "00000100",14481 => "11001111",14482 => "01110010",14483 => "00011101",14484 => "01100100",14485 => "11100001",14486 => "10001111",14487 => "11010101",14488 => "11000001",14489 => "11011001",14490 => "10101000",14491 => "10110100",14492 => "01100111",14493 => "10111001",14494 => "10111010",14495 => "01010011",14496 => "01011100",14497 => "00110111",14498 => "10010100",14499 => "11010100",14500 => "00110011",14501 => "01011110",14502 => "11010010",14503 => "00101010",14504 => "00010010",14505 => "10100111",14506 => "01100001",14507 => "11100001",14508 => "11001001",14509 => "11011100",14510 => "10101001",14511 => "01000001",14512 => "10100101",14513 => "11000000",14514 => "10001001",14515 => "00000001",14516 => "01011001",14517 => "11111110",14518 => "00101001",14519 => "10101011",14520 => "01111010",14521 => "01011101",14522 => "01100100",14523 => "11011000",14524 => "11100001",14525 => "11100011",14526 => "10000000",14527 => "01000010",14528 => "10011101",14529 => "01011010",14530 => "11101110",14531 => "01101100",14532 => "01001110",14533 => "00010010",14534 => "10110111",14535 => "01001111",14536 => "11010101",14537 => "11011100",14538 => "00001100",14539 => "01010111",14540 => "11000001",14541 => "01001111",14542 => "11000000",14543 => "11001111",14544 => "10001101",14545 => "10011100",14546 => "00010011",14547 => "11110101",14548 => "01010001",14549 => "11111101",14550 => "00010000",14551 => "10101111",14552 => "01110000",14553 => "10000111",14554 => "00110111",14555 => "10001001",14556 => "01001111",14557 => "00001011",14558 => "10001111",14559 => "01101000",14560 => "01100011",14561 => "01010000",14562 => "10011011",14563 => "00010001",14564 => "11110110",14565 => "10110101",14566 => "01001100",14567 => "00111111",14568 => "01110000",14569 => "00101101",14570 => "00100010",14571 => "10111101",14572 => "01000011",14573 => "01111010",14574 => "01000110",14575 => "11010010",14576 => "10110111",14577 => "11100100",14578 => "10000010",14579 => "10110010",14580 => "01101101",14581 => "10100000",14582 => "10011010",14583 => "01100100",14584 => "11101100",14585 => "10101001",14586 => "00100111",14587 => "11010111",14588 => "00100010",14589 => "00000011",14590 => "00111110",14591 => "10011101",14592 => "00100000",14593 => "11000011",14594 => "11001111",14595 => "01110101",14596 => "01010011",14597 => "10000000",14598 => "00010010",14599 => "00001001",14600 => "01101111",14601 => "01100010",14602 => "01011110",14603 => "11101111",14604 => "10100110",14605 => "00001110",14606 => "01000001",14607 => "10011011",14608 => "11111101",14609 => "01100000",14610 => "10110111",14611 => "01010001",14612 => "11000100",14613 => "10110101",14614 => "00101110",14615 => "10110101",14616 => "11010110",14617 => "10101111",14618 => "01111101",14619 => "11010001",14620 => "01010000",14621 => "10110011",14622 => "11101111",14623 => "00110001",14624 => "10111011",14625 => "00001111",14626 => "10110000",14627 => "10110001",14628 => "10011101",14629 => "11011011",14630 => "01001100",14631 => "00100100",14632 => "11001110",14633 => "11101100",14634 => "00110110",14635 => "11111110",14636 => "00011101",14637 => "00110001",14638 => "10100110",14639 => "00111110",14640 => "01000000",14641 => "10101001",14642 => "11010111",14643 => "01101101",14644 => "10111100",14645 => "00010110",14646 => "10110001",14647 => "01001110",14648 => "01011001",14649 => "00111110",14650 => "11110101",14651 => "00001010",14652 => "00100000",14653 => "00010100",14654 => "01101110",14655 => "00011001",14656 => "00000101",14657 => "00001101",14658 => "00011011",14659 => "01001010",14660 => "00001111",14661 => "10001110",14662 => "00101001",14663 => "11111001",14664 => "11010100",14665 => "01011110",14666 => "01101010",14667 => "01111011",14668 => "01010011",14669 => "00000000",14670 => "10011011",14671 => "10110111",14672 => "11100010",14673 => "01000100",14674 => "00010100",14675 => "00010110",14676 => "11000011",14677 => "11101100",14678 => "00011010",14679 => "10010010",14680 => "01001001",14681 => "01000101",14682 => "00001010",14683 => "11001011",14684 => "11001100",14685 => "01000100",14686 => "00110000",14687 => "10000010",14688 => "01111000",14689 => "01000000",14690 => "10100101",14691 => "00000010",14692 => "11101001",14693 => "00101101",14694 => "01111111",14695 => "01010110",14696 => "11100000",14697 => "10000000",14698 => "10111111",14699 => "00010001",14700 => "00100010",14701 => "01010010",14702 => "10011101",14703 => "11110010",14704 => "11010010",14705 => "00110111",14706 => "11010101",14707 => "10101101",14708 => "01010110",14709 => "01111101",14710 => "11000010",14711 => "00110000",14712 => "10101000",14713 => "10011100",14714 => "10010100",14715 => "10011010",14716 => "00100001",14717 => "10011011",14718 => "01101011",14719 => "10110011",14720 => "10010011",14721 => "11110010",14722 => "00001110",14723 => "10110000",14724 => "10110100",14725 => "10100110",14726 => "11000011",14727 => "00010010",14728 => "00000001",14729 => "00001111",14730 => "11100010",14731 => "00111001",14732 => "11101100",14733 => "00110010",14734 => "01110000",14735 => "00111010",14736 => "00010001",14737 => "01001000",14738 => "01011000",14739 => "11111110",14740 => "00010001",14741 => "11110100",14742 => "00111110",14743 => "10000101",14744 => "10010101",14745 => "10110101",14746 => "01001001",14747 => "10110100",14748 => "10011111",14749 => "01011001",14750 => "00101111",14751 => "01011010",14752 => "01010010",14753 => "01110110",14754 => "00110111",14755 => "00011110",14756 => "01100101",14757 => "00000010",14758 => "10101111",14759 => "11010111",14760 => "10110111",14761 => "00001101",14762 => "01001100",14763 => "10011100",14764 => "11001010",14765 => "10001001",14766 => "11110010",14767 => "00101010",14768 => "01010000",14769 => "00010110",14770 => "10001100",14771 => "00111101",14772 => "10111001",14773 => "11000000",14774 => "11010100",14775 => "00000001",14776 => "00101100",14777 => "11101100",14778 => "01101011",14779 => "11011001",14780 => "10001101",14781 => "11110101",14782 => "00011110",14783 => "10101101",14784 => "10001001",14785 => "00011010",14786 => "11110100",14787 => "10110000",14788 => "10101001",14789 => "10011100",14790 => "11110000",14791 => "11111000",14792 => "00101010",14793 => "01110110",14794 => "01111000",14795 => "00111000",14796 => "01001010",14797 => "10110111",14798 => "00100000",14799 => "10100000",14800 => "01001101",14801 => "11000111",14802 => "00010001",14803 => "10110111",14804 => "10101110",14805 => "11001011",14806 => "10111010",14807 => "10110101",14808 => "00100000",14809 => "11101100",14810 => "00111101",14811 => "10100011",14812 => "00110100",14813 => "11111111",14814 => "11110100",14815 => "01100011",14816 => "11001011",14817 => "01011001",14818 => "01101101",14819 => "10101111",14820 => "01000001",14821 => "00110011",14822 => "00110100",14823 => "11001101",14824 => "01001010",14825 => "00001111",14826 => "01111100",14827 => "10110100",14828 => "10101000",14829 => "01000010",14830 => "11110010",14831 => "01101010",14832 => "11010001",14833 => "00010100",14834 => "11000000",14835 => "00010111",14836 => "11101100",14837 => "00100001",14838 => "00100000",14839 => "00111101",14840 => "10101001",14841 => "01110011",14842 => "00111011",14843 => "11100101",14844 => "01011010",14845 => "01111110",14846 => "11000101",14847 => "01100101",14848 => "01111111",14849 => "00001000",14850 => "11001011",14851 => "10011100",14852 => "00010100",14853 => "11110110",14854 => "01110110",14855 => "01101000",14856 => "00110000",14857 => "01110110",14858 => "11001101",14859 => "11001111",14860 => "01101001",14861 => "00000101",14862 => "11100111",14863 => "00110010",14864 => "01111101",14865 => "11010111",14866 => "01001011",14867 => "10001101",14868 => "11101100",14869 => "11010001",14870 => "11000000",14871 => "00100101",14872 => "11010101",14873 => "10110111",14874 => "00000000",14875 => "10110011",14876 => "10000001",14877 => "01100110",14878 => "10010011",14879 => "11111110",14880 => "00010101",14881 => "00110111",14882 => "01110100",14883 => "11110101",14884 => "01011101",14885 => "11110101",14886 => "01110000",14887 => "00110110",14888 => "00111101",14889 => "11100000",14890 => "00011110",14891 => "11011101",14892 => "00001110",14893 => "00001111",14894 => "01000101",14895 => "11110011",14896 => "10111100",14897 => "11000111",14898 => "01111111",14899 => "11010000",14900 => "10011000",14901 => "00000000",14902 => "01000011",14903 => "11101101",14904 => "00110101",14905 => "01111000",14906 => "11100001",14907 => "01011011",14908 => "11111100",14909 => "00110110",14910 => "01011100",14911 => "01101001",14912 => "01010101",14913 => "11001010",14914 => "01110101",14915 => "11101011",14916 => "01011010",14917 => "10111110",14918 => "01001101",14919 => "00100000",14920 => "00110000",14921 => "11011100",14922 => "00000111",14923 => "01101111",14924 => "10001100",14925 => "01100010",14926 => "11001110",14927 => "01011110",14928 => "11110001",14929 => "11001100",14930 => "01110100",14931 => "00100011",14932 => "10010100",14933 => "10110111",14934 => "01010110",14935 => "00100000",14936 => "00100000",14937 => "10000010",14938 => "01101001",14939 => "11111001",14940 => "01100100",14941 => "11100001",14942 => "11001111",14943 => "01101010",14944 => "00011111",14945 => "11100101",14946 => "10000110",14947 => "11101010",14948 => "00000110",14949 => "10001101",14950 => "10110110",14951 => "01010111",14952 => "11001011",14953 => "10100011",14954 => "00110011",14955 => "10001011",14956 => "11111111",14957 => "10010010",14958 => "01110111",14959 => "00011101",14960 => "11011011",14961 => "00000101",14962 => "00101100",14963 => "10100101",14964 => "00100010",14965 => "01101101",14966 => "00010011",14967 => "11110100",14968 => "10000010",14969 => "10010101",14970 => "11011011",14971 => "11011111",14972 => "11111000",14973 => "01001010",14974 => "10011110",14975 => "10010101",14976 => "01011111",14977 => "00110111",14978 => "11100100",14979 => "10100001",14980 => "10110010",14981 => "00010111",14982 => "11011100",14983 => "10101110",14984 => "01011000",14985 => "11110000",14986 => "01110001",14987 => "00010001",14988 => "11011001",14989 => "01001101",14990 => "00001111",14991 => "00001101",14992 => "11010110",14993 => "10000101",14994 => "11011110",14995 => "11010000",14996 => "01111111",14997 => "11011001",14998 => "01010000",14999 => "01011100",15000 => "01100001",15001 => "01111001",15002 => "01111110",15003 => "10111100",15004 => "01001000",15005 => "11111100",15006 => "01100110",15007 => "10111011",15008 => "01000001",15009 => "10001111",15010 => "11100111",15011 => "11110100",15012 => "01110100",15013 => "00011010",15014 => "11010010",15015 => "00110010",15016 => "01001110",15017 => "00011111",15018 => "10100100",15019 => "01010000",15020 => "10110101",15021 => "10110011",15022 => "01111000",15023 => "11101101",15024 => "00000111",15025 => "10000011",15026 => "00101100",15027 => "01101011",15028 => "10100100",15029 => "00000010",15030 => "00111000",15031 => "11011101",15032 => "11101001",15033 => "11110111",15034 => "00110011",15035 => "11000011",15036 => "11010100",15037 => "10101100",15038 => "00110011",15039 => "01001011",15040 => "00011010",15041 => "00010110",15042 => "00000000",15043 => "01110100",15044 => "00101100",15045 => "10010010",15046 => "11010000",15047 => "10000100",15048 => "01100001",15049 => "00010100",15050 => "10011001",15051 => "11011110",15052 => "11110001",15053 => "10100101",15054 => "01000000",15055 => "00010110",15056 => "11001110",15057 => "00010110",15058 => "11110000",15059 => "10011111",15060 => "01101001",15061 => "01111010",15062 => "11001011",15063 => "01010000",15064 => "01111101",15065 => "01011101",15066 => "11001010",15067 => "01100110",15068 => "10100100",15069 => "11110000",15070 => "10101110",15071 => "10001000",15072 => "11100100",15073 => "01001100",15074 => "00100010",15075 => "01100001",15076 => "00111010",15077 => "11000101",15078 => "11000001",15079 => "01011000",15080 => "00010000",15081 => "11101001",15082 => "10110010",15083 => "11011000",15084 => "11001011",15085 => "10101011",15086 => "00101000",15087 => "01001101",15088 => "01011000",15089 => "00111110",15090 => "11111110",15091 => "11100111",15092 => "10100010",15093 => "11000110",15094 => "10010101",15095 => "11101010",15096 => "10111111",15097 => "00101110",15098 => "10110111",15099 => "00010011",15100 => "10101100",15101 => "00101000",15102 => "11001110",15103 => "01111010",15104 => "00001011",15105 => "00001110",15106 => "10111110",15107 => "01010010",15108 => "00000100",15109 => "01001101",15110 => "00010000",15111 => "01110100",15112 => "11000100",15113 => "00001000",15114 => "10010101",15115 => "00100101",15116 => "11100110",15117 => "11111101",15118 => "01000011",15119 => "01101111",15120 => "00011011",15121 => "00110001",15122 => "10101111",15123 => "00101100",15124 => "01000110",15125 => "00101001",15126 => "01101100",15127 => "01010101",15128 => "10001101",15129 => "11100111",15130 => "00111000",15131 => "00111100",15132 => "00010101",15133 => "10110000",15134 => "10000101",15135 => "00110111",15136 => "01100110",15137 => "11001010",15138 => "01111111",15139 => "10111110",15140 => "10111000",15141 => "01010101",15142 => "11110000",15143 => "00001011",15144 => "00110000",15145 => "01101011",15146 => "10100010",15147 => "10111011",15148 => "01010000",15149 => "10111110",15150 => "11100101",15151 => "10100100",15152 => "10111111",15153 => "01011100",15154 => "11101001",15155 => "10001110",15156 => "10100111",15157 => "01000011",15158 => "01000010",15159 => "11100001",15160 => "10010100",15161 => "00111110",15162 => "10001100",15163 => "11010101",15164 => "00001110",15165 => "01000001",15166 => "00010010",15167 => "10011110",15168 => "00010000",15169 => "10111000",15170 => "00011111",15171 => "01001011",15172 => "10100001",15173 => "01001001",15174 => "10000010",15175 => "10001100",15176 => "01111110",15177 => "01101110",15178 => "00011111",15179 => "11000110",15180 => "11111110",15181 => "10111101",15182 => "01101110",15183 => "01111011",15184 => "01101010",15185 => "10110001",15186 => "01001011",15187 => "01110010",15188 => "10000101",15189 => "11111011",15190 => "00000101",15191 => "00101001",15192 => "01110100",15193 => "10001101",15194 => "01010101",15195 => "11101101",15196 => "01001101",15197 => "01000001",15198 => "00000111",15199 => "01011101",15200 => "00001010",15201 => "00100110",15202 => "10000101",15203 => "11100001",15204 => "01100000",15205 => "01101001",15206 => "10111010",15207 => "11011011",15208 => "01010111",15209 => "01111011",15210 => "01000110",15211 => "00111000",15212 => "10011101",15213 => "01111000",15214 => "11010011",15215 => "01010011",15216 => "01100010",15217 => "10100001",15218 => "11011000",15219 => "10111010",15220 => "01101010",15221 => "10000111",15222 => "01101100",15223 => "11010011",15224 => "01100000",15225 => "01110101",15226 => "00111100",15227 => "11011100",15228 => "11011111",15229 => "00110110",15230 => "00101111",15231 => "01111111",15232 => "01001010",15233 => "00000010",15234 => "11111111",15235 => "01001000",15236 => "11001111",15237 => "11000101",15238 => "00010011",15239 => "01000111",15240 => "00100101",15241 => "00001100",15242 => "01011110",15243 => "00011000",15244 => "01010100",15245 => "00000111",15246 => "11000101",15247 => "01101000",15248 => "11100011",15249 => "00001001",15250 => "01001110",15251 => "11110001",15252 => "01000001",15253 => "01011101",15254 => "01011011",15255 => "01001111",15256 => "00010010",15257 => "11100010",15258 => "10011111",15259 => "01101011",15260 => "11111010",15261 => "01100001",15262 => "10000110",15263 => "11001001",15264 => "01010010",15265 => "00110000",15266 => "00100001",15267 => "01111000",15268 => "00110010",15269 => "01111001",15270 => "11110010",15271 => "11110010",15272 => "01110111",15273 => "01110101",15274 => "00001011",15275 => "10011000",15276 => "10100111",15277 => "11100111",15278 => "11101000",15279 => "00110011",15280 => "10101011",15281 => "00111000",15282 => "10001011",15283 => "10010101",15284 => "10001100",15285 => "01000110",15286 => "01111001",15287 => "11110011",15288 => "01011000",15289 => "11100010",15290 => "01000110",15291 => "01101100",15292 => "01001011",15293 => "00101001",15294 => "01000100",15295 => "01001101",15296 => "01110110",15297 => "01100111",15298 => "01110111",15299 => "00011100",15300 => "00001010",15301 => "11100011",15302 => "01001010",15303 => "10110101",15304 => "01111010",15305 => "00110111",15306 => "11000110",15307 => "11101100",15308 => "01101011",15309 => "10000101",15310 => "01010111",15311 => "00000010",15312 => "10100011",15313 => "10011001",15314 => "11111010",15315 => "10110011",15316 => "10101110",15317 => "00110110",15318 => "11000100",15319 => "01010010",15320 => "11001111",15321 => "11101000",15322 => "01100001",15323 => "11111000",15324 => "11011000",15325 => "00110010",15326 => "11110110",15327 => "01110100",15328 => "11000111",15329 => "11010111",15330 => "11011010",15331 => "10111110",15332 => "11101011",15333 => "11111101",15334 => "10111110",15335 => "11111101",15336 => "00011010",15337 => "10010101",15338 => "01000011",15339 => "11010100",15340 => "01000001",15341 => "11010101",15342 => "11111111",15343 => "00100010",15344 => "01010111",15345 => "11011010",15346 => "01011111",15347 => "11101111",15348 => "10010110",15349 => "01110100",15350 => "10011001",15351 => "11101100",15352 => "11010100",15353 => "11010010",15354 => "01100001",15355 => "11100000",15356 => "11000110",15357 => "11010001",15358 => "00100111",15359 => "00110110",15360 => "01111110",15361 => "00110000",15362 => "01010001",15363 => "00010101",15364 => "10011111",15365 => "01000100",15366 => "10011100",15367 => "00111100",15368 => "00001101",15369 => "11100110",15370 => "10011111",15371 => "00110110",15372 => "11110101",15373 => "01100010",15374 => "01011010",15375 => "00001001",15376 => "11000011",15377 => "01000110",15378 => "10101000",15379 => "01001001",15380 => "01010111",15381 => "00011010",15382 => "00000100",15383 => "00010011",15384 => "10001110",15385 => "00101000",15386 => "00000010",15387 => "01101010",15388 => "01100001",15389 => "11000101",15390 => "00111101",15391 => "11011110",15392 => "01111011",15393 => "00100111",15394 => "11100011",15395 => "01001111",15396 => "00110110",15397 => "01111000",15398 => "10110010",15399 => "10010000",15400 => "00010111",15401 => "11110011",15402 => "11000100",15403 => "10001110",15404 => "01011100",15405 => "10100101",15406 => "01000000",15407 => "11101001",15408 => "11010100",15409 => "01110101",15410 => "11111110",15411 => "00101000",15412 => "00101011",15413 => "11011111",15414 => "10010101",15415 => "01000110",15416 => "10011011",15417 => "00101110",15418 => "10100111",15419 => "00101111",15420 => "00011011",15421 => "01000111",15422 => "11101001",15423 => "10001010",15424 => "10100001",15425 => "11110100",15426 => "10101010",15427 => "11110011",15428 => "10011010",15429 => "01100010",15430 => "10110100",15431 => "10101010",15432 => "11011000",15433 => "11110011",15434 => "01000010",15435 => "00111001",15436 => "11101100",15437 => "10001101",15438 => "11100100",15439 => "00100100",15440 => "01000101",15441 => "00010110",15442 => "10011101",15443 => "01100010",15444 => "00000001",15445 => "01110000",15446 => "10101010",15447 => "01101010",15448 => "10000001",15449 => "10100011",15450 => "11100101",15451 => "10110110",15452 => "01010000",15453 => "01101101",15454 => "01111001",15455 => "10011110",15456 => "11001111",15457 => "11110011",15458 => "01010101",15459 => "10101101",15460 => "00101011",15461 => "10010101",15462 => "10100011",15463 => "00111111",15464 => "00101011",15465 => "00110111",15466 => "01000010",15467 => "01100001",15468 => "00110110",15469 => "11000000",15470 => "00111110",15471 => "01110111",15472 => "11000001",15473 => "00100000",15474 => "10000110",15475 => "11001011",15476 => "10010101",15477 => "00100000",15478 => "10011110",15479 => "11101111",15480 => "00101010",15481 => "00011010",15482 => "11011101",15483 => "01111000",15484 => "10100111",15485 => "01011011",15486 => "01001110",15487 => "01101101",15488 => "11001101",15489 => "10001010",15490 => "11001111",15491 => "11000110",15492 => "10101011",15493 => "10011111",15494 => "01100011",15495 => "10001011",15496 => "11110101",15497 => "10000001",15498 => "10100110",15499 => "01111000",15500 => "00111001",15501 => "01100000",15502 => "01101101",15503 => "10011010",15504 => "00011010",15505 => "00111000",15506 => "11110101",15507 => "10100100",15508 => "00100100",15509 => "11010101",15510 => "10101010",15511 => "10010110",15512 => "00111011",15513 => "10110011",15514 => "11110001",15515 => "01000000",15516 => "11101101",15517 => "10001001",15518 => "10010100",15519 => "11101111",15520 => "01010101",15521 => "10101100",15522 => "00010111",15523 => "01100011",15524 => "00001010",15525 => "00010101",15526 => "10001010",15527 => "00011110",15528 => "00100101",15529 => "00100100",15530 => "10111111",15531 => "00010101",15532 => "10111110",15533 => "01001000",15534 => "11101101",15535 => "01010000",15536 => "00001000",15537 => "00100101",15538 => "10010001",15539 => "01110110",15540 => "11010000",15541 => "10001000",15542 => "10010101",15543 => "01100011",15544 => "10111101",15545 => "00001011",15546 => "10100110",15547 => "01011100",15548 => "10111010",15549 => "00101100",15550 => "11011100",15551 => "01101111",15552 => "10000101",15553 => "00110010",15554 => "10111001",15555 => "01101010",15556 => "00000000",15557 => "11110001",15558 => "01111101",15559 => "01100001",15560 => "10001011",15561 => "01100001",15562 => "01110101",15563 => "01110111",15564 => "10101110",15565 => "11000111",15566 => "01001100",15567 => "01110000",15568 => "00110000",15569 => "00000111",15570 => "00111111",15571 => "00101000",15572 => "11111101",15573 => "11101010",15574 => "01110100",15575 => "01101010",15576 => "10100001",15577 => "11101000",15578 => "11100001",15579 => "10011110",15580 => "11011100",15581 => "00011001",15582 => "01101110",15583 => "01101011",15584 => "11100100",15585 => "00010000",15586 => "10011111",15587 => "11100010",15588 => "10111100",15589 => "00010110",15590 => "01100100",15591 => "10010010",15592 => "11000010",15593 => "00101011",15594 => "00110011",15595 => "11110110",15596 => "10110110",15597 => "11011101",15598 => "00110100",15599 => "10010100",15600 => "01010011",15601 => "01100010",15602 => "01101011",15603 => "11110110",15604 => "10111001",15605 => "10111011",15606 => "10101011",15607 => "00011010",15608 => "11101010",15609 => "10100110",15610 => "01000111",15611 => "00011011",15612 => "00111111",15613 => "00100011",15614 => "11000000",15615 => "11110010",15616 => "01111111",15617 => "01111001",15618 => "10010111",15619 => "00100000",15620 => "10011100",15621 => "00010101",15622 => "01101010",15623 => "11001101",15624 => "11001000",15625 => "11101001",15626 => "10010000",15627 => "11011110",15628 => "00011000",15629 => "10000011",15630 => "00101111",15631 => "00110000",15632 => "01111011",15633 => "10000110",15634 => "01000111",15635 => "11111100",15636 => "01111100",15637 => "01100000",15638 => "01000010",15639 => "00000110",15640 => "11000000",15641 => "01101100",15642 => "11100111",15643 => "11110110",15644 => "00010111",15645 => "10010100",15646 => "11110010",15647 => "11010111",15648 => "10001010",15649 => "00001000",15650 => "00000011",15651 => "01110101",15652 => "00001111",15653 => "01101010",15654 => "10111101",15655 => "11111110",15656 => "00100010",15657 => "01010101",15658 => "00101000",15659 => "01111000",15660 => "11011110",15661 => "11100111",15662 => "10001000",15663 => "01001100",15664 => "00110110",15665 => "11101111",15666 => "00011000",15667 => "11100011",15668 => "10110000",15669 => "11100111",15670 => "00010001",15671 => "00000010",15672 => "10011010",15673 => "10000010",15674 => "01100110",15675 => "11010011",15676 => "00000011",15677 => "00111110",15678 => "00110101",15679 => "10101100",15680 => "10001110",15681 => "01100000",15682 => "01101011",15683 => "11001001",15684 => "11100111",15685 => "11110000",15686 => "10011000",15687 => "11110100",15688 => "11110001",15689 => "00010101",15690 => "01001001",15691 => "11110110",15692 => "01111101",15693 => "00110111",15694 => "11000010",15695 => "01110101",15696 => "01011010",15697 => "00010110",15698 => "00000101",15699 => "00100010",15700 => "01101000",15701 => "10001110",15702 => "10100001",15703 => "01000101",15704 => "01111110",15705 => "00001111",15706 => "00110001",15707 => "11111011",15708 => "00111001",15709 => "10101100",15710 => "01110010",15711 => "01110001",15712 => "00110100",15713 => "11100010",15714 => "10111101",15715 => "10110111",15716 => "11001110",15717 => "10100110",15718 => "11001111",15719 => "00110100",15720 => "11010001",15721 => "00100111",15722 => "11001010",15723 => "11000011",15724 => "00100110",15725 => "10011001",15726 => "10100011",15727 => "10111110",15728 => "01010001",15729 => "01011000",15730 => "10101011",15731 => "00001101",15732 => "11110101",15733 => "10101101",15734 => "00001111",15735 => "00111001",15736 => "10010010",15737 => "11110100",15738 => "10101111",15739 => "10000010",15740 => "10011100",15741 => "01010011",15742 => "10011000",15743 => "11101000",15744 => "10100100",15745 => "11011100",15746 => "00011100",15747 => "01001110",15748 => "00111110",15749 => "01110010",15750 => "00011111",15751 => "11101001",15752 => "01100101",15753 => "00100101",15754 => "00000010",15755 => "01000010",15756 => "10101011",15757 => "10011100",15758 => "00100010",15759 => "11101000",15760 => "10000010",15761 => "11111110",15762 => "01111101",15763 => "00010011",15764 => "11110110",15765 => "10001011",15766 => "01000001",15767 => "10001011",15768 => "11110100",15769 => "01111001",15770 => "01000111",15771 => "00100100",15772 => "11001110",15773 => "00100110",15774 => "01011011",15775 => "10010111",15776 => "10101000",15777 => "01100111",15778 => "00100001",15779 => "10001110",15780 => "01111110",15781 => "10111010",15782 => "00101011",15783 => "00101100",15784 => "11000001",15785 => "01110011",15786 => "11101010",15787 => "00110011",15788 => "10011011",15789 => "00010111",15790 => "01100111",15791 => "11010010",15792 => "00100010",15793 => "00001111",15794 => "01000010",15795 => "10101011",15796 => "01001001",15797 => "10101000",15798 => "00111111",15799 => "01100010",15800 => "00101100",15801 => "00011111",15802 => "01110001",15803 => "11111011",15804 => "11010010",15805 => "00101101",15806 => "11111110",15807 => "11011010",15808 => "01111110",15809 => "01001010",15810 => "01111100",15811 => "10000111",15812 => "01011111",15813 => "01111101",15814 => "00100011",15815 => "00000000",15816 => "11111011",15817 => "11100000",15818 => "01010011",15819 => "11011001",15820 => "10100011",15821 => "10001001",15822 => "11000100",15823 => "10101101",15824 => "11010010",15825 => "11100001",15826 => "01100011",15827 => "10000001",15828 => "01000110",15829 => "10111100",15830 => "11011000",15831 => "10000110",15832 => "10110111",15833 => "10111100",15834 => "10000110",15835 => "11000011",15836 => "10001000",15837 => "00010100",15838 => "11000011",15839 => "01110101",15840 => "01110001",15841 => "11001101",15842 => "01001110",15843 => "10001011",15844 => "10101001",15845 => "10110100",15846 => "11011010",15847 => "11010101",15848 => "00000001",15849 => "11011001",15850 => "10110111",15851 => "01000111",15852 => "10110100",15853 => "11001101",15854 => "11101001",15855 => "10111110",15856 => "10011100",15857 => "00100011",15858 => "01100000",15859 => "01011111",15860 => "10010111",15861 => "10001100",15862 => "01010110",15863 => "11101110",15864 => "01000100",15865 => "01011001",15866 => "01101111",15867 => "11101110",15868 => "10010111",15869 => "11100101",15870 => "10000010",15871 => "00010000",15872 => "00010111",15873 => "11101100",15874 => "01010111",15875 => "00000101",15876 => "10001010",15877 => "10100111",15878 => "00101001",15879 => "11100111",15880 => "01100001",15881 => "10101011",15882 => "01100100",15883 => "10110111",15884 => "10100110",15885 => "11011100",15886 => "11011110",15887 => "00100000",15888 => "11110011",15889 => "10100101",15890 => "00001100",15891 => "10111010",15892 => "00010011",15893 => "00110101",15894 => "10001000",15895 => "10101110",15896 => "11101001",15897 => "11001000",15898 => "10101010",15899 => "10010010",15900 => "11011100",15901 => "01101011",15902 => "01000000",15903 => "00000001",15904 => "10000110",15905 => "10100000",15906 => "11101011",15907 => "00011101",15908 => "11101110",15909 => "01001110",15910 => "00010010",15911 => "00011111",15912 => "01000010",15913 => "10110001",15914 => "11111000",15915 => "11110101",15916 => "11000001",15917 => "01101011",15918 => "10001011",15919 => "11101001",15920 => "11111001",15921 => "01010110",15922 => "10010101",15923 => "10010101",15924 => "11000000",15925 => "00000001",15926 => "01110100",15927 => "00110001",15928 => "10011101",15929 => "10111010",15930 => "10001011",15931 => "00000001",15932 => "11010000",15933 => "00110101",15934 => "11001111",15935 => "01001010",15936 => "01011101",15937 => "10010000",15938 => "11101110",15939 => "00000011",15940 => "10010011",15941 => "11000101",15942 => "11110101",15943 => "00111001",15944 => "10010000",15945 => "00100110",15946 => "10010100",15947 => "11001110",15948 => "11100110",15949 => "10100010",15950 => "10000111",15951 => "01010110",15952 => "00000110",15953 => "11000100",15954 => "11101101",15955 => "01010011",15956 => "01010010",15957 => "01011000",15958 => "11111000",15959 => "11110010",15960 => "11101101",15961 => "01011010",15962 => "11000111",15963 => "10010100",15964 => "11111100",15965 => "11001101",15966 => "01101101",15967 => "00100110",15968 => "01000011",15969 => "11111110",15970 => "01000001",15971 => "01010011",15972 => "00010101",15973 => "01001010",15974 => "00110010",15975 => "10001100",15976 => "00111010",15977 => "10101111",15978 => "10000010",15979 => "00000111",15980 => "11000001",15981 => "11001010",15982 => "01111011",15983 => "11100111",15984 => "00001011",15985 => "11010111",15986 => "11001001",15987 => "11011110",15988 => "01000010",15989 => "10001110",15990 => "10001101",15991 => "00100010",15992 => "00010010",15993 => "11010111",15994 => "01010110",15995 => "01100111",15996 => "00010101",15997 => "11100010",15998 => "10110101",15999 => "00110010",16000 => "01000100",16001 => "00000011",16002 => "10110010",16003 => "10000101",16004 => "01111100",16005 => "10011101",16006 => "10001111",16007 => "10010110",16008 => "11110000",16009 => "11101010",16010 => "11001101",16011 => "00101101",16012 => "01001000",16013 => "10111010",16014 => "10000001",16015 => "11110101",16016 => "10010111",16017 => "00101101",16018 => "00101110",16019 => "01010000",16020 => "00111000",16021 => "11000011",16022 => "10110011",16023 => "10100111",16024 => "01100111",16025 => "01100010",16026 => "11011110",16027 => "11110101",16028 => "00111100",16029 => "10101100",16030 => "00010000",16031 => "00100010",16032 => "10000100",16033 => "10111110",16034 => "01011010",16035 => "10100010",16036 => "10101111",16037 => "01100010",16038 => "01111110",16039 => "01011011",16040 => "11111011",16041 => "01101101",16042 => "00010110",16043 => "01111111",16044 => "00110001",16045 => "00011110",16046 => "11010011",16047 => "00101000",16048 => "11011000",16049 => "01010011",16050 => "00010010",16051 => "01111111",16052 => "10010000",16053 => "10001010",16054 => "10100000",16055 => "01110101",16056 => "10000110",16057 => "10100110",16058 => "11000011",16059 => "11000110",16060 => "01100111",16061 => "00000001",16062 => "01001100",16063 => "10011101",16064 => "10110111",16065 => "01100000",16066 => "01011101",16067 => "11100000",16068 => "11100011",16069 => "10111010",16070 => "00101000",16071 => "10011100",16072 => "11110001",16073 => "11001111",16074 => "01111100",16075 => "01111100",16076 => "01111111",16077 => "01011100",16078 => "00001011",16079 => "00110010",16080 => "11111100",16081 => "10001110",16082 => "11010010",16083 => "00000011",16084 => "10110100",16085 => "11010001",16086 => "00101100",16087 => "01101011",16088 => "00110100",16089 => "11010101",16090 => "01100111",16091 => "10000010",16092 => "10110110",16093 => "11000000",16094 => "01110110",16095 => "11100100",16096 => "00111000",16097 => "10101001",16098 => "00010101",16099 => "11000110",16100 => "10010011",16101 => "00010101",16102 => "00110100",16103 => "00010110",16104 => "10110010",16105 => "10011110",16106 => "11100011",16107 => "01001101",16108 => "11011110",16109 => "11101001",16110 => "11000001",16111 => "00101010",16112 => "10000001",16113 => "00010010",16114 => "10011101",16115 => "00101100",16116 => "00111111",16117 => "01110011",16118 => "11011110",16119 => "10001100",16120 => "11010100",16121 => "01011011",16122 => "11100001",16123 => "11011100",16124 => "11101000",16125 => "00100000",16126 => "00010010",16127 => "10111000",16128 => "10100101",16129 => "01100010",16130 => "11000011",16131 => "10111010",16132 => "10010111",16133 => "11011000",16134 => "10110001",16135 => "01100010",16136 => "10010011",16137 => "00101100",16138 => "11010100",16139 => "10101001",16140 => "01101111",16141 => "01010010",16142 => "00110111",16143 => "00101111",16144 => "11110100",16145 => "10101101",16146 => "10001101",16147 => "00110110",16148 => "10111100",16149 => "00011111",16150 => "10111111",16151 => "00000000",16152 => "01111000",16153 => "01000011",16154 => "01011100",16155 => "11000100",16156 => "11001111",16157 => "11000101",16158 => "01111000",16159 => "01010001",16160 => "01100001",16161 => "01000101",16162 => "00110001",16163 => "10000011",16164 => "11010100",16165 => "01011011",16166 => "10011011",16167 => "01001100",16168 => "00010001",16169 => "00101001",16170 => "01100101",16171 => "01010101",16172 => "01100000",16173 => "11010011",16174 => "10011110",16175 => "01100110",16176 => "00100010",16177 => "11110000",16178 => "10111010",16179 => "11010101",16180 => "10010001",16181 => "01111111",16182 => "11010000",16183 => "01100010",16184 => "10011100",16185 => "00010101",16186 => "00001001",16187 => "01101110",16188 => "10100011",16189 => "11000111",16190 => "11001111",16191 => "00110110",16192 => "00011001",16193 => "01111100",16194 => "01100010",16195 => "11111011",16196 => "01111011",16197 => "10101110",16198 => "01001010",16199 => "01000010",16200 => "10110101",16201 => "00110100",16202 => "01001000",16203 => "11010000",16204 => "11111111",16205 => "01111001",16206 => "01111000",16207 => "10010001",16208 => "00101000",16209 => "10011111",16210 => "10000010",16211 => "00110100",16212 => "11010010",16213 => "00000011",16214 => "00111000",16215 => "10101010",16216 => "11010010",16217 => "11110100",16218 => "10110010",16219 => "10001110",16220 => "11101001",16221 => "00111111",16222 => "00001011",16223 => "11000010",16224 => "11100011",16225 => "10110011",16226 => "00011010",16227 => "10000100",16228 => "01011101",16229 => "11011001",16230 => "11000000",16231 => "00101010",16232 => "11011001",16233 => "11100111",16234 => "11000110",16235 => "00110110",16236 => "11111101",16237 => "11011001",16238 => "11011000",16239 => "00011010",16240 => "01101101",16241 => "01110011",16242 => "01000000",16243 => "00111010",16244 => "11000111",16245 => "01111100",16246 => "01111100",16247 => "11000111",16248 => "10011111",16249 => "11101001",16250 => "01101001",16251 => "00101101",16252 => "01010010",16253 => "00110000",16254 => "10000000",16255 => "11011111",16256 => "01100101",16257 => "01001011",16258 => "00000111",16259 => "10111001",16260 => "00000111",16261 => "01110110",16262 => "00011001",16263 => "10100101",16264 => "10010011",16265 => "10100110",16266 => "00101101",16267 => "10111011",16268 => "01001100",16269 => "10000011",16270 => "10001000",16271 => "11001100",16272 => "01011111",16273 => "00101101",16274 => "00110000",16275 => "10111101",16276 => "10100100",16277 => "10011000",16278 => "01011111",16279 => "11101000",16280 => "01101100",16281 => "11001101",16282 => "00101111",16283 => "10100010",16284 => "00000001",16285 => "10000100",16286 => "00001100",16287 => "00010111",16288 => "10100000",16289 => "01111101",16290 => "10110111",16291 => "11001000",16292 => "00010110",16293 => "11110100",16294 => "10111110",16295 => "10110100",16296 => "00000110",16297 => "00001101",16298 => "10100000",16299 => "10000010",16300 => "11000111",16301 => "10011001",16302 => "10110001",16303 => "10101101",16304 => "11111110",16305 => "01011011",16306 => "01100000",16307 => "01001011",16308 => "01000001",16309 => "01010000",16310 => "01111010",16311 => "10011110",16312 => "10101101",16313 => "10000010",16314 => "01001101",16315 => "00101010",16316 => "10010110",16317 => "01110100",16318 => "11111010",16319 => "00011001",16320 => "01011001",16321 => "10000011",16322 => "01101100",16323 => "00111100",16324 => "01111011",16325 => "01110100",16326 => "10110100",16327 => "10110011",16328 => "00011000",16329 => "10001110",16330 => "10010001",16331 => "01110010",16332 => "11001101",16333 => "11100101",16334 => "10100111",16335 => "10101011",16336 => "01000110",16337 => "11101101",16338 => "01110010",16339 => "00010111",16340 => "11010101",16341 => "01110000",16342 => "10001011",16343 => "00100100",16344 => "10101010",16345 => "01111101",16346 => "01001100",16347 => "11111110",16348 => "01011011",16349 => "01100110",16350 => "11011000",16351 => "10001000",16352 => "01100000",16353 => "01100001",16354 => "01110010",16355 => "00110011",16356 => "01010011",16357 => "00110101",16358 => "10001110",16359 => "11010010",16360 => "11100110",16361 => "11010100",16362 => "11101110",16363 => "11100111",16364 => "00000110",16365 => "10000100",16366 => "10110000",16367 => "10000010",16368 => "00011011",16369 => "11111111",16370 => "11101111",16371 => "11011101",16372 => "00001011",16373 => "01010111",16374 => "11111100",16375 => "10001111",16376 => "01110010",16377 => "11111001",16378 => "00000111",16379 => "01111100",16380 => "01011011",16381 => "10110111",16382 => "10001101",16383 => "01111010",16384 => "11001100",16385 => "00111100",16386 => "11111011",16387 => "01010100",16388 => "01100110",16389 => "00001111",16390 => "01110011",16391 => "11000101",16392 => "00010111",16393 => "01110011",16394 => "11101101",16395 => "10000011",16396 => "10101011",16397 => "00111011",16398 => "11101101",16399 => "01111000",16400 => "00001000",16401 => "01110101",16402 => "01100101",16403 => "10111110",16404 => "01011110",16405 => "11011101",16406 => "11000011",16407 => "10010001",16408 => "11101111",16409 => "11001000",16410 => "11100100",16411 => "00011010",16412 => "01100111",16413 => "00111010",16414 => "11001011",16415 => "11011000",16416 => "00011100",16417 => "11111000",16418 => "00111011",16419 => "00010110",16420 => "11011011",16421 => "11000110",16422 => "01000001",16423 => "01011110",16424 => "11101000",16425 => "10011000",16426 => "10111100",16427 => "10100111",16428 => "01000010",16429 => "01001101",16430 => "00010101",16431 => "00001011",16432 => "01110000",16433 => "00010010",16434 => "01010110",16435 => "00001111",16436 => "00010110",16437 => "11110101",16438 => "10010100",16439 => "10111000",16440 => "10111000",16441 => "00000000",16442 => "10001011",16443 => "01000100",16444 => "11110000",16445 => "11110011",16446 => "00100000",16447 => "00100110",16448 => "00111101",16449 => "11011101",16450 => "10000000",16451 => "11000110",16452 => "11001100",16453 => "10000011",16454 => "11110100",16455 => "11100000",16456 => "11010001",16457 => "11000001",16458 => "00011110",16459 => "01110100",16460 => "11011001",16461 => "01000010",16462 => "11100010",16463 => "00100100",16464 => "00111001",16465 => "10100001",16466 => "01000110",16467 => "01010011",16468 => "10010010",16469 => "01111100",16470 => "11011101",16471 => "00100111",16472 => "11101010",16473 => "00010010",16474 => "01101001",16475 => "01001110",16476 => "11001011",16477 => "00011000",16478 => "01110100",16479 => "10001111",16480 => "01010110",16481 => "01111011",16482 => "01100100",16483 => "11010000",16484 => "01111111",16485 => "01111000",16486 => "11110111",16487 => "01101110",16488 => "00001111",16489 => "00110010",16490 => "11110101",16491 => "01110111",16492 => "10100100",16493 => "00001011",16494 => "10000011",16495 => "01110010",16496 => "10101101",16497 => "01010111",16498 => "01100100",16499 => "01111101",16500 => "00011100",16501 => "10110011",16502 => "10000111",16503 => "10110011",16504 => "00000111",16505 => "01101010",16506 => "01001111",16507 => "10001111",16508 => "10111001",16509 => "11101000",16510 => "01110001",16511 => "01101110",16512 => "10101001",16513 => "01110000",16514 => "01000011",16515 => "01100010",16516 => "01111100",16517 => "11011000",16518 => "01010001",16519 => "01110111",16520 => "10001011",16521 => "10100111",16522 => "11011001",16523 => "01000011",16524 => "11111111",16525 => "01011100",16526 => "00110110",16527 => "01101001",16528 => "10001001",16529 => "10110011",16530 => "11001111",16531 => "11101011",16532 => "00010001",16533 => "10111111",16534 => "10111000",16535 => "01010110",16536 => "11100110",16537 => "11100110",16538 => "00110110",16539 => "01110111",16540 => "10011101",16541 => "01010010",16542 => "00101111",16543 => "11001000",16544 => "01011000",16545 => "10001000",16546 => "01100101",16547 => "11110011",16548 => "11101111",16549 => "11001001",16550 => "10110001",16551 => "00111001",16552 => "01001110",16553 => "11011011",16554 => "01101101",16555 => "01100001",16556 => "00010010",16557 => "00011010",16558 => "00000010",16559 => "11011101",16560 => "00001010",16561 => "00100011",16562 => "00011101",16563 => "00001100",16564 => "10000110",16565 => "00010001",16566 => "01011010",16567 => "11000110",16568 => "00100010",16569 => "11000101",16570 => "01111111",16571 => "00010001",16572 => "11000000",16573 => "10111001",16574 => "10000001",16575 => "10001001",16576 => "10100111",16577 => "10001110",16578 => "10101010",16579 => "11100110",16580 => "10101110",16581 => "01001011",16582 => "11000101",16583 => "10011011",16584 => "11011010",16585 => "00000101",16586 => "00001010",16587 => "00101111",16588 => "11110011",16589 => "10100100",16590 => "11010001",16591 => "10000100",16592 => "00111101",16593 => "00010101",16594 => "10011010",16595 => "11000011",16596 => "10110110",16597 => "01011010",16598 => "10110010",16599 => "00100100",16600 => "11001111",16601 => "10101000",16602 => "11101111",16603 => "10001010",16604 => "10010001",16605 => "10101001",16606 => "11110110",16607 => "00110000",16608 => "11011011",16609 => "01010000",16610 => "01011001",16611 => "10011010",16612 => "10001100",16613 => "00001111",16614 => "00110000",16615 => "01110100",16616 => "01101011",16617 => "11100010",16618 => "00001110",16619 => "11001111",16620 => "10101011",16621 => "01101001",16622 => "11011111",16623 => "01000001",16624 => "01100000",16625 => "10100111",16626 => "00010001",16627 => "01101001",16628 => "00111110",16629 => "01110000",16630 => "00001110",16631 => "10100010",16632 => "11110110",16633 => "11000010",16634 => "11110110",16635 => "01000100",16636 => "00011001",16637 => "10101001",16638 => "00101101",16639 => "11001100",16640 => "11111010",16641 => "00101101",16642 => "00110011",16643 => "01101101",16644 => "01111011",16645 => "00101001",16646 => "00001011",16647 => "10101111",16648 => "01111111",16649 => "10111110",16650 => "01010100",16651 => "01110010",16652 => "00110101",16653 => "10100101",16654 => "11011000",16655 => "11100100",16656 => "01001100",16657 => "01001010",16658 => "11001011",16659 => "11011111",16660 => "11001101",16661 => "01011101",16662 => "11010011",16663 => "00101101",16664 => "11001100",16665 => "10010100",16666 => "10011101",16667 => "11011001",16668 => "01011011",16669 => "11001010",16670 => "11011010",16671 => "00110011",16672 => "00101010",16673 => "00101000",16674 => "00000100",16675 => "00000010",16676 => "11110011",16677 => "10100001",16678 => "10011101",16679 => "10001010",16680 => "10100100",16681 => "01100001",16682 => "11011111",16683 => "11001100",16684 => "01011001",16685 => "11111111",16686 => "11011010",16687 => "11101010",16688 => "10101110",16689 => "00111101",16690 => "11110001",16691 => "00001001",16692 => "10101010",16693 => "11010000",16694 => "11110001",16695 => "10101111",16696 => "10101001",16697 => "10100000",16698 => "11001010",16699 => "11101100",16700 => "01001101",16701 => "01001101",16702 => "11001100",16703 => "10110100",16704 => "00100011",16705 => "00111111",16706 => "10010001",16707 => "11111000",16708 => "00000101",16709 => "11001000",16710 => "01011010",16711 => "11100100",16712 => "10100111",16713 => "00111101",16714 => "01100101",16715 => "00101110",16716 => "01110011",16717 => "00101000",16718 => "00111101",16719 => "00001111",16720 => "01010000",16721 => "01010010",16722 => "10011111",16723 => "10110010",16724 => "10100000",16725 => "01000010",16726 => "01111101",16727 => "01110001",16728 => "11100111",16729 => "00011001",16730 => "01000000",16731 => "00111101",16732 => "11101000",16733 => "10010111",16734 => "01001111",16735 => "01000000",16736 => "01110010",16737 => "10110110",16738 => "00101110",16739 => "01110110",16740 => "10011011",16741 => "01001100",16742 => "01001111",16743 => "10110100",16744 => "00010001",16745 => "00101111",16746 => "01101110",16747 => "01101110",16748 => "00101110",16749 => "01100001",16750 => "00001000",16751 => "10110111",16752 => "11100011",16753 => "00011000",16754 => "10011110",16755 => "10101101",16756 => "01011010",16757 => "00011100",16758 => "11101011",16759 => "10111111",16760 => "00011101",16761 => "11011011",16762 => "01101010",16763 => "00010100",16764 => "11110010",16765 => "00010111",16766 => "01110010",16767 => "00010111",16768 => "00101010",16769 => "00111011",16770 => "00100010",16771 => "01000100",16772 => "11111111",16773 => "11110110",16774 => "01101101",16775 => "00111110",16776 => "11100010",16777 => "10110100",16778 => "01001010",16779 => "01111000",16780 => "11110110",16781 => "00101000",16782 => "11110100",16783 => "10001010",16784 => "01001110",16785 => "00011111",16786 => "11100010",16787 => "11101010",16788 => "01001100",16789 => "11111100",16790 => "01011100",16791 => "00111000",16792 => "10001011",16793 => "00001010",16794 => "11110101",16795 => "01110001",16796 => "10100010",16797 => "01010000",16798 => "01011000",16799 => "01011001",16800 => "00010001",16801 => "10001000",16802 => "10001001",16803 => "10111100",16804 => "01001000",16805 => "01101101",16806 => "01110110",16807 => "00010110",16808 => "10101000",16809 => "10101110",16810 => "11111001",16811 => "01101110",16812 => "11101010",16813 => "10111000",16814 => "01001101",16815 => "01011011",16816 => "10011100",16817 => "01010101",16818 => "00101011",16819 => "10100001",16820 => "01100101",16821 => "01000110",16822 => "00001101",16823 => "01111111",16824 => "01011100",16825 => "10001000",16826 => "11010000",16827 => "11101100",16828 => "00111110",16829 => "01000010",16830 => "01100000",16831 => "10101001",16832 => "10011101",16833 => "10000000",16834 => "11101101",16835 => "11011110",16836 => "01011101",16837 => "00001010",16838 => "01111100",16839 => "00001100",16840 => "00100101",16841 => "01101111",16842 => "01010111",16843 => "11111111",16844 => "01100011",16845 => "01110110",16846 => "01110111",16847 => "01110100",16848 => "00011110",16849 => "00010000",16850 => "01110110",16851 => "10000010",16852 => "10100001",16853 => "10111011",16854 => "10101110",16855 => "01001110",16856 => "10100101",16857 => "01100101",16858 => "00001101",16859 => "10011111",16860 => "01010010",16861 => "10010001",16862 => "11111010",16863 => "11110001",16864 => "00001100",16865 => "11010100",16866 => "00010111",16867 => "10010100",16868 => "11100101",16869 => "00011101",16870 => "00110100",16871 => "10100100",16872 => "11111110",16873 => "10000001",16874 => "10010110",16875 => "10010010",16876 => "10010001",16877 => "10110100",16878 => "11000011",16879 => "01011000",16880 => "01101010",16881 => "00111111",16882 => "01111110",16883 => "11000101",16884 => "00100110",16885 => "00101101",16886 => "01100011",16887 => "10011001",16888 => "10010001",16889 => "10011010",16890 => "00111110",16891 => "11001101",16892 => "01100111",16893 => "00000000",16894 => "10010100",16895 => "01100010",16896 => "01111110",16897 => "10110010",16898 => "10010100",16899 => "11010000",16900 => "00000001",16901 => "10100000",16902 => "11100111",16903 => "11010110",16904 => "10111101",16905 => "00100011",16906 => "10110001",16907 => "01110000",16908 => "00010001",16909 => "10010011",16910 => "10101001",16911 => "01010010",16912 => "01000111",16913 => "11100000",16914 => "01111100",16915 => "10110010",16916 => "00100011",16917 => "01101000",16918 => "01100001",16919 => "01100010",16920 => "10011101",16921 => "00000100",16922 => "10001000",16923 => "10010110",16924 => "11010011",16925 => "11000101",16926 => "01110100",16927 => "10001000",16928 => "10010000",16929 => "01000000",16930 => "01111001",16931 => "10000101",16932 => "00001010",16933 => "10001010",16934 => "10000011",16935 => "10011111",16936 => "00001011",16937 => "10010011",16938 => "00111111",16939 => "10110011",16940 => "10001010",16941 => "01001000",16942 => "00111111",16943 => "01100011",16944 => "10100011",16945 => "00001010",16946 => "01001101",16947 => "01001011",16948 => "00100111",16949 => "10100111",16950 => "11100011",16951 => "00011100",16952 => "10101011",16953 => "10111001",16954 => "11110111",16955 => "00110101",16956 => "11011001",16957 => "01100011",16958 => "01011010",16959 => "01001001",16960 => "01111011",16961 => "10000100",16962 => "00001001",16963 => "10100010",16964 => "10101111",16965 => "10100000",16966 => "11100101",16967 => "01011111",16968 => "01110101",16969 => "00111101",16970 => "10101110",16971 => "11001010",16972 => "10101101",16973 => "00011111",16974 => "01011111",16975 => "10100001",16976 => "10011010",16977 => "11001110",16978 => "01111100",16979 => "11000100",16980 => "01010001",16981 => "00110100",16982 => "01000101",16983 => "11111010",16984 => "11111010",16985 => "00110010",16986 => "11011011",16987 => "11110000",16988 => "11100010",16989 => "01100001",16990 => "00100111",16991 => "11000011",16992 => "01001111",16993 => "00111110",16994 => "01101111",16995 => "01010111",16996 => "00111110",16997 => "01011111",16998 => "00011100",16999 => "00001000",17000 => "01111101",17001 => "00110001",17002 => "01110111",17003 => "10000011",17004 => "01101110",17005 => "11010011",17006 => "00111000",17007 => "10001110",17008 => "10011000",17009 => "01011010",17010 => "01010001",17011 => "01100101",17012 => "11000110",17013 => "01001111",17014 => "11011000",17015 => "11011110",17016 => "01001011",17017 => "10111100",17018 => "00010110",17019 => "11000011",17020 => "10000010",17021 => "11101100",17022 => "11101101",17023 => "11100101",17024 => "10000100",17025 => "11110111",17026 => "11001011",17027 => "10111011",17028 => "11100100",17029 => "10100000",17030 => "10101100",17031 => "00000000",17032 => "00100111",17033 => "01000011",17034 => "00100011",17035 => "10010110",17036 => "10100111",17037 => "00010010",17038 => "10011101",17039 => "00101110",17040 => "01011100",17041 => "10111111",17042 => "00000011",17043 => "01011111",17044 => "10100001",17045 => "01001011",17046 => "01001110",17047 => "10111011",17048 => "01111010",17049 => "01000011",17050 => "11100010",17051 => "01000000",17052 => "10100111",17053 => "10011111",17054 => "01001001",17055 => "00011000",17056 => "01100011",17057 => "01011010",17058 => "00110010",17059 => "11001100",17060 => "10111101",17061 => "11001101",17062 => "10111000",17063 => "10101111",17064 => "00101101",17065 => "11100011",17066 => "01111111",17067 => "01011010",17068 => "11000110",17069 => "11110101",17070 => "11110000",17071 => "01101110",17072 => "10000101",17073 => "11111110",17074 => "11101101",17075 => "11100010",17076 => "10110110",17077 => "11000001",17078 => "01100000",17079 => "00001101",17080 => "00000010",17081 => "01000001",17082 => "01010010",17083 => "01110111",17084 => "11101000",17085 => "00110000",17086 => "01010010",17087 => "11101010",17088 => "00000000",17089 => "10101000",17090 => "01111010",17091 => "01110010",17092 => "11111010",17093 => "10110010",17094 => "11100010",17095 => "00001110",17096 => "01010000",17097 => "10111000",17098 => "00000110",17099 => "11100011",17100 => "00001101",17101 => "00000010",17102 => "11100001",17103 => "10011111",17104 => "11010000",17105 => "11011000",17106 => "00111000",17107 => "00011000",17108 => "10110000",17109 => "01101111",17110 => "01011110",17111 => "00000110",17112 => "10110001",17113 => "00010010",17114 => "10101010",17115 => "01001111",17116 => "10001011",17117 => "01011000",17118 => "01010100",17119 => "00110101",17120 => "10101000",17121 => "00100011",17122 => "00000111",17123 => "11010110",17124 => "01001010",17125 => "01101110",17126 => "10011001",17127 => "10100011",17128 => "10000001",17129 => "00111100",17130 => "11101001",17131 => "00111110",17132 => "11011111",17133 => "00000101",17134 => "01011011",17135 => "10010010",17136 => "00001100",17137 => "10000001",17138 => "01111010",17139 => "11101000",17140 => "10100110",17141 => "00010001",17142 => "00000001",17143 => "11000001",17144 => "01100110",17145 => "10101001",17146 => "00011011",17147 => "11000001",17148 => "10111011",17149 => "11000101",17150 => "11100001",17151 => "11110110",17152 => "11000111",17153 => "10001111",17154 => "10100111",17155 => "00110100",17156 => "10111000",17157 => "11011000",17158 => "01101001",17159 => "11111010",17160 => "11100001",17161 => "01101100",17162 => "01111001",17163 => "10011010",17164 => "11110100",17165 => "01000101",17166 => "01101010",17167 => "00000101",17168 => "11111011",17169 => "01100110",17170 => "00001111",17171 => "01001101",17172 => "10011111",17173 => "11110001",17174 => "10010101",17175 => "10010100",17176 => "01100100",17177 => "01111100",17178 => "11110111",17179 => "01011101",17180 => "11001100",17181 => "11100011",17182 => "11100001",17183 => "00100011",17184 => "01010100",17185 => "10100000",17186 => "01100001",17187 => "11001101",17188 => "11111001",17189 => "10100010",17190 => "10101110",17191 => "01101100",17192 => "00001011",17193 => "00010000",17194 => "10110110",17195 => "01101011",17196 => "00011111",17197 => "10001000",17198 => "01001100",17199 => "11101101",17200 => "01101010",17201 => "00000010",17202 => "10001111",17203 => "00010100",17204 => "01100100",17205 => "10101010",17206 => "00010010",17207 => "00011101",17208 => "00101110",17209 => "10001011",17210 => "01011111",17211 => "10110100",17212 => "10101000",17213 => "01100000",17214 => "10010101",17215 => "11101101",17216 => "10111101",17217 => "00010001",17218 => "00100111",17219 => "10111110",17220 => "00111111",17221 => "01010000",17222 => "11010011",17223 => "01101011",17224 => "10101100",17225 => "01111001",17226 => "01011111",17227 => "10000100",17228 => "00001101",17229 => "00111111",17230 => "00101101",17231 => "01100110",17232 => "01010010",17233 => "10001101",17234 => "01110101",17235 => "11100011",17236 => "11000111",17237 => "10101010",17238 => "01111010",17239 => "00100001",17240 => "10011100",17241 => "10011001",17242 => "01110100",17243 => "10100110",17244 => "01001100",17245 => "00110010",17246 => "01000100",17247 => "00100111",17248 => "00100011",17249 => "11101101",17250 => "01100110",17251 => "11111111",17252 => "01000101",17253 => "00101100",17254 => "00100000",17255 => "11111011",17256 => "11000100",17257 => "10001111",17258 => "10010001",17259 => "01111000",17260 => "10100001",17261 => "11010110",17262 => "10001100",17263 => "00110100",17264 => "10001110",17265 => "00101110",17266 => "11010000",17267 => "00100001",17268 => "01001101",17269 => "00100101",17270 => "11010001",17271 => "01000101",17272 => "10011110",17273 => "11100101",17274 => "11000001",17275 => "10011101",17276 => "10000000",17277 => "00000011",17278 => "11100000",17279 => "00000010",17280 => "01110101",17281 => "11110001",17282 => "00110101",17283 => "00111010",17284 => "00000100",17285 => "11111111",17286 => "01011001",17287 => "01010111",17288 => "00010011",17289 => "10000110",17290 => "01110000",17291 => "10110100",17292 => "10100100",17293 => "10110111",17294 => "11111000",17295 => "00100000",17296 => "11011111",17297 => "10011110",17298 => "10001101",17299 => "01101001",17300 => "10111000",17301 => "01100111",17302 => "00001111",17303 => "00101110",17304 => "11100001",17305 => "11110111",17306 => "01011110",17307 => "01001100",17308 => "10011110",17309 => "01010010",17310 => "01000010",17311 => "11011101",17312 => "01010100",17313 => "00111010",17314 => "10110100",17315 => "11100011",17316 => "10111100",17317 => "00010000",17318 => "11010001",17319 => "10011000",17320 => "11111010",17321 => "11111100",17322 => "10110011",17323 => "10100101",17324 => "00100100",17325 => "01110100",17326 => "00011101",17327 => "10110000",17328 => "00100010",17329 => "01001101",17330 => "11011010",17331 => "00110011",17332 => "00110010",17333 => "00100001",17334 => "00000101",17335 => "11100100",17336 => "01010011",17337 => "00010001",17338 => "11001011",17339 => "00011110",17340 => "01101100",17341 => "11011001",17342 => "01110011",17343 => "11111111",17344 => "01100001",17345 => "01001111",17346 => "00000001",17347 => "00001111",17348 => "01110111",17349 => "10100110",17350 => "10000110",17351 => "10001111",17352 => "01011010",17353 => "00001000",17354 => "11001000",17355 => "00001111",17356 => "01000110",17357 => "11101100",17358 => "10000101",17359 => "11011010",17360 => "01001100",17361 => "00100010",17362 => "00001001",17363 => "10111110",17364 => "11101000",17365 => "10110111",17366 => "11011000",17367 => "10010101",17368 => "11001111",17369 => "10110111",17370 => "00100110",17371 => "10110110",17372 => "10011110",17373 => "00010110",17374 => "01000001",17375 => "11100111",17376 => "01001000",17377 => "01111011",17378 => "10111011",17379 => "11111100",17380 => "01000110",17381 => "01111100",17382 => "00100010",17383 => "01100101",17384 => "01100100",17385 => "01100101",17386 => "00101010",17387 => "10001110",17388 => "00101110",17389 => "11001101",17390 => "01100000",17391 => "00111101",17392 => "10011111",17393 => "10011100",17394 => "00101011",17395 => "01111010",17396 => "01000000",17397 => "00001000",17398 => "01000101",17399 => "10001011",17400 => "11011001",17401 => "10000001",17402 => "11110001",17403 => "10011100",17404 => "00000001",17405 => "01110001",17406 => "10011011",17407 => "10001001",17408 => "00110111",17409 => "11100011",17410 => "00011111",17411 => "10001010",17412 => "11001000",17413 => "00011111",17414 => "00111110",17415 => "00100100",17416 => "11001111",17417 => "00010101",17418 => "01110101",17419 => "10010110",17420 => "10011010",17421 => "11000101",17422 => "01001101",17423 => "11111010",17424 => "11111010",17425 => "00101101",17426 => "10011100",17427 => "00101110",17428 => "01010100",17429 => "00111110",17430 => "10010110",17431 => "10001101",17432 => "01010011",17433 => "00101010",17434 => "01000000",17435 => "10000010",17436 => "00101010",17437 => "10101001",17438 => "01100100",17439 => "00001011",17440 => "10001010",17441 => "10100100",17442 => "00100000",17443 => "01100111",17444 => "01100000",17445 => "01101010",17446 => "01000110",17447 => "00110110",17448 => "11100011",17449 => "00101110",17450 => "10001010",17451 => "11110001",17452 => "10110101",17453 => "11111010",17454 => "00101101",17455 => "11001011",17456 => "11110010",17457 => "00010111",17458 => "00010110",17459 => "01010110",17460 => "11000000",17461 => "11011100",17462 => "01010101",17463 => "11111101",17464 => "11111110",17465 => "01010001",17466 => "00111011",17467 => "01111010",17468 => "11110011",17469 => "00100100",17470 => "00000100",17471 => "10100001",17472 => "01110001",17473 => "01010000",17474 => "10111101",17475 => "00011110",17476 => "00001000",17477 => "01001000",17478 => "00000111",17479 => "01001011",17480 => "00010010",17481 => "11100001",17482 => "01101110",17483 => "01111000",17484 => "11101010",17485 => "11100111",17486 => "01000000",17487 => "10000010",17488 => "11101100",17489 => "10010110",17490 => "01011110",17491 => "01001101",17492 => "01001010",17493 => "01110000",17494 => "10000011",17495 => "10010000",17496 => "11011001",17497 => "00110100",17498 => "11111011",17499 => "01001100",17500 => "00111001",17501 => "01101100",17502 => "01001100",17503 => "00101101",17504 => "10011101",17505 => "01001101",17506 => "00111000",17507 => "01011010",17508 => "10011111",17509 => "01001100",17510 => "11111001",17511 => "11110011",17512 => "10000100",17513 => "01001100",17514 => "11001000",17515 => "11100011",17516 => "11100010",17517 => "01110101",17518 => "10110001",17519 => "11001001",17520 => "01110001",17521 => "00110110",17522 => "00110011",17523 => "00111111",17524 => "10010100",17525 => "00010000",17526 => "01000010",17527 => "10111100",17528 => "01010000",17529 => "11000010",17530 => "11110010",17531 => "10111010",17532 => "01010111",17533 => "00110100",17534 => "10011110",17535 => "00110011",17536 => "00011110",17537 => "01110100",17538 => "01000101",17539 => "10011101",17540 => "00110101",17541 => "10110001",17542 => "01101010",17543 => "01000001",17544 => "11010000",17545 => "00101111",17546 => "11011011",17547 => "00100011",17548 => "11110011",17549 => "10010001",17550 => "11110001",17551 => "01010101",17552 => "01000001",17553 => "01010101",17554 => "11001011",17555 => "01010111",17556 => "00001000",17557 => "01110001",17558 => "10111011",17559 => "10110100",17560 => "10110000",17561 => "11010111",17562 => "01010100",17563 => "01111011",17564 => "11000110",17565 => "10011001",17566 => "10010000",17567 => "01111110",17568 => "00011010",17569 => "10011011",17570 => "01000101",17571 => "10111110",17572 => "10101010",17573 => "00110100",17574 => "11010001",17575 => "01000011",17576 => "01111100",17577 => "00010011",17578 => "10011101",17579 => "00100100",17580 => "11100011",17581 => "00111100",17582 => "00001101",17583 => "11011001",17584 => "00010110",17585 => "11011100",17586 => "11111110",17587 => "01011000",17588 => "01001010",17589 => "10010111",17590 => "00111010",17591 => "00110000",17592 => "10100110",17593 => "01000000",17594 => "10100010",17595 => "10000000",17596 => "01010000",17597 => "10101101",17598 => "00110101",17599 => "00101100",17600 => "01111110",17601 => "11001011",17602 => "10100100",17603 => "00001100",17604 => "00110110",17605 => "00010100",17606 => "00100110",17607 => "01101001",17608 => "10001110",17609 => "10000101",17610 => "11011011",17611 => "01101100",17612 => "00000111",17613 => "10011010",17614 => "00000010",17615 => "11000100",17616 => "01100000",17617 => "01001011",17618 => "11100100",17619 => "01010100",17620 => "10001110",17621 => "00111010",17622 => "01100000",17623 => "11101011",17624 => "01111101",17625 => "00001111",17626 => "10011100",17627 => "11100101",17628 => "00000000",17629 => "01010000",17630 => "11101110",17631 => "10000001",17632 => "10100111",17633 => "10111101",17634 => "10101001",17635 => "10100101",17636 => "11000101",17637 => "00110111",17638 => "01010010",17639 => "11111101",17640 => "00011101",17641 => "01010101",17642 => "10011011",17643 => "00011001",17644 => "11101001",17645 => "01001101",17646 => "11011001",17647 => "00111001",17648 => "11100100",17649 => "11101010",17650 => "00110111",17651 => "11010111",17652 => "10010001",17653 => "00101111",17654 => "00100101",17655 => "11100110",17656 => "00000110",17657 => "00011100",17658 => "10100000",17659 => "00000001",17660 => "00100100",17661 => "11110010",17662 => "01101010",17663 => "00011000",17664 => "10010110",17665 => "10000001",17666 => "00010110",17667 => "01111101",17668 => "00001001",17669 => "11000000",17670 => "11101000",17671 => "11110101",17672 => "10010010",17673 => "00011010",17674 => "10100100",17675 => "01000110",17676 => "10010111",17677 => "10000011",17678 => "00110011",17679 => "00011001",17680 => "11011110",17681 => "10101100",17682 => "01111111",17683 => "10001111",17684 => "11100000",17685 => "10110010",17686 => "01011100",17687 => "10011001",17688 => "10001011",17689 => "00010101",17690 => "01000110",17691 => "10100111",17692 => "01001000",17693 => "01011111",17694 => "00000000",17695 => "11001110",17696 => "11001010",17697 => "11010001",17698 => "01000101",17699 => "10010101",17700 => "11000001",17701 => "01100010",17702 => "10000000",17703 => "00010010",17704 => "01011001",17705 => "10000100",17706 => "11100001",17707 => "00101110",17708 => "01010000",17709 => "00110100",17710 => "00100010",17711 => "01101111",17712 => "11110110",17713 => "10101111",17714 => "00101100",17715 => "10101010",17716 => "00011011",17717 => "10100111",17718 => "00010110",17719 => "01111000",17720 => "11000111",17721 => "00111011",17722 => "00100110",17723 => "01111111",17724 => "11111100",17725 => "10100010",17726 => "11110100",17727 => "11101111",17728 => "01110110",17729 => "01011001",17730 => "01100101",17731 => "01101000",17732 => "10111011",17733 => "00101001",17734 => "00100011",17735 => "00111010",17736 => "01011111",17737 => "00101010",17738 => "10110101",17739 => "01111000",17740 => "01111011",17741 => "10011110",17742 => "01100010",17743 => "10101110",17744 => "01011000",17745 => "01111011",17746 => "01000111",17747 => "11010100",17748 => "11011010",17749 => "10000111",17750 => "11010000",17751 => "00010001",17752 => "00000110",17753 => "01001011",17754 => "10101100",17755 => "11100111",17756 => "10111101",17757 => "00100111",17758 => "11000010",17759 => "01101010",17760 => "10000000",17761 => "10101100",17762 => "11110111",17763 => "11000111",17764 => "00000010",17765 => "00000110",17766 => "01011011",17767 => "10100001",17768 => "10110100",17769 => "11101010",17770 => "10011001",17771 => "11000000",17772 => "11110000",17773 => "11100101",17774 => "11110011",17775 => "11100100",17776 => "01011101",17777 => "00111011",17778 => "10110010",17779 => "00010101",17780 => "11101000",17781 => "10001000",17782 => "10111010",17783 => "11110101",17784 => "01110000",17785 => "10101111",17786 => "11100011",17787 => "01000111",17788 => "11010001",17789 => "00111110",17790 => "00101101",17791 => "10001101",17792 => "11110101",17793 => "00101110",17794 => "01110011",17795 => "00000100",17796 => "00110101",17797 => "11010011",17798 => "00101111",17799 => "01000010",17800 => "10101100",17801 => "00011111",17802 => "01111101",17803 => "11100010",17804 => "11110100",17805 => "10100110",17806 => "11010110",17807 => "11101100",17808 => "11100001",17809 => "01101011",17810 => "01100101",17811 => "00010000",17812 => "00010100",17813 => "11011011",17814 => "11110000",17815 => "11111000",17816 => "00101101",17817 => "11101011",17818 => "00010110",17819 => "11100000",17820 => "00111111",17821 => "00110111",17822 => "01000110",17823 => "11101100",17824 => "00111111",17825 => "01111100",17826 => "11000001",17827 => "11001000",17828 => "10010010",17829 => "01011100",17830 => "00000000",17831 => "00000100",17832 => "00001000",17833 => "10010001",17834 => "00000001",17835 => "00001111",17836 => "11001010",17837 => "01110001",17838 => "01111011",17839 => "10101101",17840 => "00110101",17841 => "01001101",17842 => "10001000",17843 => "10011010",17844 => "00101011",17845 => "01000111",17846 => "00000010",17847 => "10111111",17848 => "00001110",17849 => "00000111",17850 => "00001101",17851 => "11011010",17852 => "00000111",17853 => "01010000",17854 => "10101110",17855 => "10010111",17856 => "11001101",17857 => "01101111",17858 => "10010111",17859 => "01110110",17860 => "10001111",17861 => "10111011",17862 => "10100101",17863 => "11110010",17864 => "00001000",17865 => "11110100",17866 => "01010101",17867 => "10010110",17868 => "11000000",17869 => "00001010",17870 => "10011000",17871 => "01110101",17872 => "11111111",17873 => "10110111",17874 => "10101101",17875 => "00110101",17876 => "10100110",17877 => "10001010",17878 => "00100001",17879 => "10010110",17880 => "10101101",17881 => "10100100",17882 => "01010000",17883 => "11110100",17884 => "10001000",17885 => "00010110",17886 => "00001111",17887 => "10100000",17888 => "10111110",17889 => "01010010",17890 => "01000001",17891 => "11101111",17892 => "00100010",17893 => "01111101",17894 => "01001111",17895 => "01000111",17896 => "10001010",17897 => "11100101",17898 => "01111100",17899 => "10111110",17900 => "10101010",17901 => "11100110",17902 => "00100100",17903 => "01000010",17904 => "00111111",17905 => "11100111",17906 => "10111111",17907 => "10001111",17908 => "10110010",17909 => "00110000",17910 => "00100101",17911 => "11011111",17912 => "10011010",17913 => "10010100",17914 => "00111100",17915 => "10010010",17916 => "11000100",17917 => "11000101",17918 => "00101101",17919 => "11010001",17920 => "11010010",17921 => "10010000",17922 => "11101000",17923 => "10110011",17924 => "01010010",17925 => "01101010",17926 => "00000101",17927 => "11011011",17928 => "10000111",17929 => "00100010",17930 => "10100010",17931 => "10001110",17932 => "00000010",17933 => "11110010",17934 => "11110110",17935 => "01001010",17936 => "11001110",17937 => "00101001",17938 => "00000000",17939 => "10010001",17940 => "00001000",17941 => "00111110",17942 => "10110011",17943 => "01011000",17944 => "00001110",17945 => "00010010",17946 => "00010010",17947 => "10101101",17948 => "00010100",17949 => "01010011",17950 => "10110000",17951 => "01010011",17952 => "01011100",17953 => "11011011",17954 => "00001010",17955 => "11110010",17956 => "01100000",17957 => "00001101",17958 => "00100010",17959 => "11100100",17960 => "11001011",17961 => "01110111",17962 => "00101101",17963 => "11010000",17964 => "01010111",17965 => "00001011",17966 => "01100110",17967 => "10010000",17968 => "10100110",17969 => "00010000",17970 => "00100001",17971 => "11110010",17972 => "00000010",17973 => "00000110",17974 => "10100111",17975 => "01111011",17976 => "10001100",17977 => "11011010",17978 => "11111111",17979 => "10110101",17980 => "11010001",17981 => "00101110",17982 => "00000010",17983 => "01010101",17984 => "10001110",17985 => "00111110",17986 => "10000110",17987 => "01000111",17988 => "10111101",17989 => "01010001",17990 => "01011111",17991 => "10110011",17992 => "10100000",17993 => "01011110",17994 => "11100111",17995 => "11000111",17996 => "01100011",17997 => "10011111",17998 => "10000111",17999 => "10011100",18000 => "10110110",18001 => "01010010",18002 => "00001101",18003 => "00011111",18004 => "11100111",18005 => "10010110",18006 => "11111000",18007 => "10111101",18008 => "00010111",18009 => "00001110",18010 => "01010101",18011 => "01011111",18012 => "01101001",18013 => "01111000",18014 => "10101010",18015 => "11110010",18016 => "01101100",18017 => "11000011",18018 => "01110110",18019 => "10110110",18020 => "01110010",18021 => "11000101",18022 => "01110101",18023 => "10100101",18024 => "10010101",18025 => "10101111",18026 => "11001100",18027 => "01010000",18028 => "10100001",18029 => "01001011",18030 => "00011001",18031 => "10100110",18032 => "11110101",18033 => "00111111",18034 => "01011110",18035 => "10110010",18036 => "00001101",18037 => "11011101",18038 => "10000101",18039 => "01011000",18040 => "11011011",18041 => "00011110",18042 => "01111100",18043 => "00101100",18044 => "00101101",18045 => "01111000",18046 => "11100000",18047 => "00010110",18048 => "10010101",18049 => "00110111",18050 => "01100100",18051 => "01011101",18052 => "01111111",18053 => "01000010",18054 => "10100100",18055 => "11000100",18056 => "00010000",18057 => "00111000",18058 => "00010000",18059 => "11000110",18060 => "00100100",18061 => "11001011",18062 => "10101000",18063 => "01111001",18064 => "11101111",18065 => "10001110",18066 => "00111101",18067 => "00011001",18068 => "11110010",18069 => "11000111",18070 => "10000101",18071 => "01100100",18072 => "01101111",18073 => "11001000",18074 => "00101010",18075 => "00000011",18076 => "01000010",18077 => "10100111",18078 => "11100110",18079 => "01011001",18080 => "01000110",18081 => "10110110",18082 => "00100110",18083 => "01110101",18084 => "11100101",18085 => "10110111",18086 => "11001010",18087 => "10000101",18088 => "10110100",18089 => "11001101",18090 => "10010011",18091 => "00001101",18092 => "01101011",18093 => "01101100",18094 => "01000011",18095 => "11100011",18096 => "01001100",18097 => "01100011",18098 => "01001010",18099 => "01001010",18100 => "01011000",18101 => "01111111",18102 => "01101111",18103 => "01010101",18104 => "00110010",18105 => "00011010",18106 => "11100110",18107 => "01111100",18108 => "10101100",18109 => "11111010",18110 => "10011110",18111 => "10110011",18112 => "00010110",18113 => "10011101",18114 => "00000101",18115 => "10001110",18116 => "11000010",18117 => "01111100",18118 => "10100001",18119 => "01110101",18120 => "11110110",18121 => "11001111",18122 => "10010001",18123 => "11000110",18124 => "01010010",18125 => "10101111",18126 => "10110000",18127 => "10101000",18128 => "10100101",18129 => "00101110",18130 => "11111111",18131 => "01111000",18132 => "10011001",18133 => "10000111",18134 => "00001000",18135 => "10011011",18136 => "01110111",18137 => "00010111",18138 => "10010101",18139 => "01010100",18140 => "10001000",18141 => "10101000",18142 => "10000100",18143 => "11000110",18144 => "00011011",18145 => "11110001",18146 => "00010100",18147 => "10000010",18148 => "10110111",18149 => "11000001",18150 => "01100111",18151 => "00110100",18152 => "11101111",18153 => "01011000",18154 => "10101011",18155 => "01011001",18156 => "10111001",18157 => "11010111",18158 => "01011010",18159 => "10100011",18160 => "10010100",18161 => "11011110",18162 => "10001011",18163 => "11001111",18164 => "01000100",18165 => "00111100",18166 => "11100001",18167 => "00101010",18168 => "00010001",18169 => "00101100",18170 => "01110011",18171 => "01010111",18172 => "10100010",18173 => "00101010",18174 => "01100000",18175 => "11111001",18176 => "01110101",18177 => "10000000",18178 => "10000000",18179 => "01110010",18180 => "10100000",18181 => "01000001",18182 => "11110101",18183 => "10100100",18184 => "01101111",18185 => "11101111",18186 => "01001101",18187 => "00100000",18188 => "11110101",18189 => "11001000",18190 => "01100010",18191 => "11100111",18192 => "11110110",18193 => "10011100",18194 => "00010100",18195 => "00001110",18196 => "11010110",18197 => "10100110",18198 => "00010001",18199 => "10001010",18200 => "01001101",18201 => "10001101",18202 => "11001101",18203 => "10011010",18204 => "00110010",18205 => "00001011",18206 => "01000010",18207 => "00000101",18208 => "10011010",18209 => "10000110",18210 => "00000101",18211 => "01111100",18212 => "00110000",18213 => "10111111",18214 => "00110010",18215 => "11000111",18216 => "10011110",18217 => "10111001",18218 => "01011000",18219 => "10001001",18220 => "01010110",18221 => "00110111",18222 => "01001000",18223 => "01110111",18224 => "11111110",18225 => "00011000",18226 => "00101010",18227 => "11011000",18228 => "01001000",18229 => "10100101",18230 => "11010011",18231 => "10011010",18232 => "11101001",18233 => "11111101",18234 => "11010011",18235 => "10100001",18236 => "00001111",18237 => "11011110",18238 => "00101010",18239 => "01101101",18240 => "01001110",18241 => "10100110",18242 => "00010111",18243 => "00000101",18244 => "01111110",18245 => "00000101",18246 => "10010110",18247 => "01001110",18248 => "11101000",18249 => "11010111",18250 => "11111100",18251 => "00110011",18252 => "10011101",18253 => "11011001",18254 => "10011111",18255 => "00011100",18256 => "10101000",18257 => "10111000",18258 => "10101010",18259 => "10110011",18260 => "00000011",18261 => "11011000",18262 => "11011000",18263 => "10101011",18264 => "00000011",18265 => "11111001",18266 => "01101010",18267 => "00001010",18268 => "11010010",18269 => "10100111",18270 => "01010101",18271 => "00101011",18272 => "00000010",18273 => "11001100",18274 => "00011011",18275 => "00100001",18276 => "10110101",18277 => "00101101",18278 => "00011111",18279 => "11100110",18280 => "10110111",18281 => "00100000",18282 => "10111101",18283 => "01010011",18284 => "10001000",18285 => "11000101",18286 => "10001010",18287 => "01000010",18288 => "00111100",18289 => "11010110",18290 => "00011010",18291 => "10111000",18292 => "10011110",18293 => "00001001",18294 => "10101101",18295 => "01111111",18296 => "00001000",18297 => "10100000",18298 => "11001100",18299 => "10001010",18300 => "00101101",18301 => "01111001",18302 => "01000000",18303 => "01000100",18304 => "01111010",18305 => "01001010",18306 => "01100011",18307 => "11000100",18308 => "11001111",18309 => "10010101",18310 => "00010100",18311 => "00000000",18312 => "11100110",18313 => "00100111",18314 => "10010000",18315 => "00111000",18316 => "00100010",18317 => "11010001",18318 => "11110111",18319 => "11011101",18320 => "10011000",18321 => "10000110",18322 => "00101101",18323 => "10110111",18324 => "00010111",18325 => "11011100",18326 => "11001110",18327 => "01000010",18328 => "01011110",18329 => "10010100",18330 => "10010100",18331 => "00010101",18332 => "10110000",18333 => "01010101",18334 => "11100101",18335 => "00111110",18336 => "00000111",18337 => "00010011",18338 => "10000111",18339 => "10010010",18340 => "10000111",18341 => "01000110",18342 => "01001001",18343 => "00000101",18344 => "01110110",18345 => "10110110",18346 => "01100110",18347 => "00111100",18348 => "11000001",18349 => "11010011",18350 => "01110100",18351 => "01011010",18352 => "11011011",18353 => "11110110",18354 => "11101111",18355 => "10100110",18356 => "01011100",18357 => "10100111",18358 => "11111100",18359 => "00101111",18360 => "00111111",18361 => "10101110",18362 => "11101111",18363 => "11000000",18364 => "01010011",18365 => "11001011",18366 => "00011011",18367 => "10010000",18368 => "10100011",18369 => "00000110",18370 => "11101011",18371 => "11010001",18372 => "00001100",18373 => "10010100",18374 => "01000101",18375 => "00110111",18376 => "10111010",18377 => "01101101",18378 => "01100101",18379 => "01010100",18380 => "10000110",18381 => "11111110",18382 => "10101010",18383 => "11001111",18384 => "01100111",18385 => "00110100",18386 => "00111010",18387 => "00001011",18388 => "01000110",18389 => "01000101",18390 => "00010110",18391 => "10100010",18392 => "10101011",18393 => "00010101",18394 => "11101011",18395 => "10100110",18396 => "00010000",18397 => "00101100",18398 => "11001010",18399 => "10011110",18400 => "00101001",18401 => "10001011",18402 => "01100011",18403 => "00111110",18404 => "01101101",18405 => "11100001",18406 => "10011011",18407 => "10110110",18408 => "00001101",18409 => "10001110",18410 => "01101111",18411 => "11011111",18412 => "10101001",18413 => "10010110",18414 => "10101100",18415 => "00100011",18416 => "11101010",18417 => "11111001",18418 => "11100011",18419 => "10101110",18420 => "10101110",18421 => "00011110",18422 => "00111010",18423 => "00100110",18424 => "00111011",18425 => "00100010",18426 => "00000100",18427 => "01011010",18428 => "01110010",18429 => "01100010",18430 => "11011100",18431 => "01011010",18432 => "11011100",18433 => "10010010",18434 => "01110110",18435 => "00010000",18436 => "00101101",18437 => "00000101",18438 => "01111110",18439 => "00011100",18440 => "00110100",18441 => "11111010",18442 => "11110000",18443 => "01111111",18444 => "00010010",18445 => "01001100",18446 => "01010010",18447 => "01001000",18448 => "00001010",18449 => "01011010",18450 => "00001111",18451 => "11010010",18452 => "10011010",18453 => "01100100",18454 => "00001010",18455 => "00101001",18456 => "11111000",18457 => "11110000",18458 => "00011000",18459 => "10010100",18460 => "11001010",18461 => "01000101",18462 => "11000101",18463 => "10000100",18464 => "01101011",18465 => "01100010",18466 => "11101101",18467 => "01101011",18468 => "01010001",18469 => "10011001",18470 => "11001100",18471 => "00010100",18472 => "00111110",18473 => "10010010",18474 => "01001011",18475 => "00000000",18476 => "00001010",18477 => "00111011",18478 => "10011111",18479 => "01101110",18480 => "00000011",18481 => "00000011",18482 => "11110101",18483 => "10110000",18484 => "01001100",18485 => "11000011",18486 => "11000000",18487 => "00101000",18488 => "10100101",18489 => "00010101",18490 => "00011110",18491 => "00100011",18492 => "00101001",18493 => "01011011",18494 => "00110101",18495 => "10000110",18496 => "01110010",18497 => "10011010",18498 => "01010000",18499 => "00011110",18500 => "11101100",18501 => "11111101",18502 => "01000100",18503 => "10110111",18504 => "00101001",18505 => "11101011",18506 => "01001111",18507 => "01111101",18508 => "00000000",18509 => "10000011",18510 => "00010101",18511 => "00100001",18512 => "10111011",18513 => "11100110",18514 => "11000111",18515 => "00100110",18516 => "11101111",18517 => "11010110",18518 => "10000010",18519 => "10011110",18520 => "01101010",18521 => "01010100",18522 => "01011010",18523 => "01101101",18524 => "11110011",18525 => "00001001",18526 => "00001001",18527 => "01000000",18528 => "01111110",18529 => "01011111",18530 => "00000110",18531 => "11001111",18532 => "01011110",18533 => "11100010",18534 => "01010111",18535 => "10111011",18536 => "10000011",18537 => "00011100",18538 => "10101011",18539 => "01000100",18540 => "00101111",18541 => "10100001",18542 => "11001100",18543 => "01000111",18544 => "00111101",18545 => "11100110",18546 => "10001100",18547 => "11100100",18548 => "01010010",18549 => "00011110",18550 => "01110011",18551 => "11111011",18552 => "00010000",18553 => "01001011",18554 => "01000001",18555 => "10101110",18556 => "11101011",18557 => "11011000",18558 => "00001101",18559 => "01010101",18560 => "01000110",18561 => "11101010",18562 => "11110011",18563 => "01001010",18564 => "10000110",18565 => "00001110",18566 => "01000000",18567 => "10101010",18568 => "10011110",18569 => "01100111",18570 => "00010110",18571 => "10011100",18572 => "00111101",18573 => "01001110",18574 => "11111010",18575 => "01110001",18576 => "11000101",18577 => "10000111",18578 => "10010010",18579 => "11010101",18580 => "11011000",18581 => "01000110",18582 => "01010001",18583 => "11110000",18584 => "00110100",18585 => "01101010",18586 => "01101000",18587 => "01000111",18588 => "11011000",18589 => "10100110",18590 => "00100110",18591 => "01100000",18592 => "01000000",18593 => "10100100",18594 => "10001100",18595 => "11010111",18596 => "00000111",18597 => "00110111",18598 => "10001011",18599 => "10110010",18600 => "11000000",18601 => "10101010",18602 => "10110100",18603 => "01110101",18604 => "10100111",18605 => "10010011",18606 => "10000011",18607 => "11110110",18608 => "10101100",18609 => "01010111",18610 => "01101100",18611 => "10011010",18612 => "11100000",18613 => "00100010",18614 => "10000110",18615 => "00111100",18616 => "10010111",18617 => "00110111",18618 => "01001000",18619 => "01110101",18620 => "11011100",18621 => "00100000",18622 => "11101011",18623 => "01100111",18624 => "11100010",18625 => "00001011",18626 => "11110101",18627 => "11101100",18628 => "11100101",18629 => "10111100",18630 => "00101010",18631 => "01000011",18632 => "10111101",18633 => "11010010",18634 => "00100111",18635 => "11100000",18636 => "11001010",18637 => "10011011",18638 => "11010000",18639 => "01010010",18640 => "10011111",18641 => "00011010",18642 => "10011111",18643 => "10010000",18644 => "10010100",18645 => "10111010",18646 => "11010110",18647 => "10001011",18648 => "00011000",18649 => "10101100",18650 => "11111001",18651 => "10000001",18652 => "00111111",18653 => "11111011",18654 => "11010011",18655 => "10111100",18656 => "01011000",18657 => "01001001",18658 => "10000001",18659 => "10101110",18660 => "11111010",18661 => "10011010",18662 => "10000011",18663 => "11111100",18664 => "10000100",18665 => "00101011",18666 => "01010101",18667 => "10010000",18668 => "01010110",18669 => "01110101",18670 => "11010101",18671 => "11001000",18672 => "10100100",18673 => "10111010",18674 => "00001011",18675 => "10010100",18676 => "00010010",18677 => "10110101",18678 => "10001101",18679 => "10100111",18680 => "01011001",18681 => "00111110",18682 => "11111001",18683 => "01111111",18684 => "01101010",18685 => "01010011",18686 => "10100100",18687 => "11111000",18688 => "00011101",18689 => "11111111",18690 => "00000110",18691 => "00101001",18692 => "10010011",18693 => "01111111",18694 => "00100110",18695 => "11100110",18696 => "01010000",18697 => "01000011",18698 => "00100101",18699 => "01001100",18700 => "11101101",18701 => "01000101",18702 => "01100010",18703 => "10001001",18704 => "10100110",18705 => "10110101",18706 => "00001000",18707 => "11000011",18708 => "01110110",18709 => "10100011",18710 => "01001101",18711 => "11101100",18712 => "00100010",18713 => "10101000",18714 => "00001100",18715 => "01110000",18716 => "11101111",18717 => "01011101",18718 => "00101010",18719 => "01000010",18720 => "00010001",18721 => "01111000",18722 => "00011010",18723 => "11111100",18724 => "10110111",18725 => "10101000",18726 => "00101110",18727 => "10010001",18728 => "00010000",18729 => "01100101",18730 => "10010000",18731 => "11101111",18732 => "11010101",18733 => "01110010",18734 => "10110100",18735 => "10110011",18736 => "01011011",18737 => "10010000",18738 => "10111101",18739 => "01001010",18740 => "10000111",18741 => "10011010",18742 => "00101010",18743 => "01111100",18744 => "01000111",18745 => "01110110",18746 => "00011000",18747 => "00000010",18748 => "11110010",18749 => "00101000",18750 => "10010111",18751 => "01110010",18752 => "01101010",18753 => "10010010",18754 => "00101111",18755 => "11010111",18756 => "00001101",18757 => "10101111",18758 => "00000100",18759 => "11110000",18760 => "01100101",18761 => "10100001",18762 => "10000110",18763 => "11110011",18764 => "10001001",18765 => "01011000",18766 => "10111001",18767 => "11111010",18768 => "10011101",18769 => "01100010",18770 => "00011101",18771 => "10011101",18772 => "01010011",18773 => "10010010",18774 => "10100110",18775 => "01001011",18776 => "10011101",18777 => "01100100",18778 => "01000011",18779 => "00011111",18780 => "01000110",18781 => "01011001",18782 => "00111000",18783 => "11111011",18784 => "01001100",18785 => "00101101",18786 => "00111101",18787 => "00100101",18788 => "11010110",18789 => "00010100",18790 => "01001000",18791 => "00001111",18792 => "00111111",18793 => "10010001",18794 => "00100110",18795 => "01101001",18796 => "11101001",18797 => "00111001",18798 => "10000000",18799 => "10111011",18800 => "00000001",18801 => "00000000",18802 => "01110101",18803 => "01000110",18804 => "10000101",18805 => "00111100",18806 => "01100110",18807 => "00111101",18808 => "01010000",18809 => "01100110",18810 => "11111010",18811 => "00101110",18812 => "10010101",18813 => "10110101",18814 => "11110011",18815 => "10011110",18816 => "01101111",18817 => "11100111",18818 => "01110101",18819 => "11001001",18820 => "11000011",18821 => "01100101",18822 => "11111100",18823 => "11001010",18824 => "00111001",18825 => "10001110",18826 => "10111000",18827 => "10101111",18828 => "10100110",18829 => "01101010",18830 => "00100111",18831 => "10000010",18832 => "00011110",18833 => "00101001",18834 => "00001111",18835 => "00001000",18836 => "10010100",18837 => "00000010",18838 => "01111011",18839 => "00111010",18840 => "10101100",18841 => "00111000",18842 => "11100010",18843 => "10010100",18844 => "00011011",18845 => "00001010",18846 => "01100000",18847 => "00010110",18848 => "01011001",18849 => "00110110",18850 => "01000000",18851 => "10111111",18852 => "00110101",18853 => "10111101",18854 => "01111111",18855 => "11001111",18856 => "10111010",18857 => "10101110",18858 => "10011110",18859 => "10011101",18860 => "00001101",18861 => "00100010",18862 => "10010100",18863 => "01010000",18864 => "00001000",18865 => "10100100",18866 => "11111000",18867 => "11010100",18868 => "01101001",18869 => "01000011",18870 => "10010111",18871 => "01000100",18872 => "00001101",18873 => "11100101",18874 => "00110111",18875 => "11111100",18876 => "11010110",18877 => "00100001",18878 => "10111001",18879 => "00110100",18880 => "00011011",18881 => "10010001",18882 => "01110010",18883 => "11010100",18884 => "00000000",18885 => "00000000",18886 => "00010110",18887 => "11000000",18888 => "01000111",18889 => "11000111",18890 => "00010001",18891 => "10101000",18892 => "11000111",18893 => "10010100",18894 => "10000101",18895 => "00111110",18896 => "00000010",18897 => "11111011",18898 => "00110001",18899 => "10111110",18900 => "01110001",18901 => "10001011",18902 => "00000011",18903 => "01101110",18904 => "01101010",18905 => "11110010",18906 => "11111100",18907 => "11011101",18908 => "10111010",18909 => "01011011",18910 => "11111010",18911 => "00101101",18912 => "01010111",18913 => "10111100",18914 => "00010101",18915 => "01010000",18916 => "11001011",18917 => "11111101",18918 => "11000110",18919 => "01110100",18920 => "10000000",18921 => "00010101",18922 => "11110101",18923 => "00011100",18924 => "00111001",18925 => "01000001",18926 => "00011100",18927 => "11001010",18928 => "00001010",18929 => "11110011",18930 => "10010001",18931 => "11110111",18932 => "00010101",18933 => "10011001",18934 => "11001000",18935 => "11110010",18936 => "01001111",18937 => "10100010",18938 => "10100010",18939 => "11011100",18940 => "01100111",18941 => "01000100",18942 => "01100111",18943 => "01101001",18944 => "00000110",18945 => "11011111",18946 => "00010110",18947 => "11101001",18948 => "00111001",18949 => "11010110",18950 => "01110100",18951 => "00111011",18952 => "10011101",18953 => "10110111",18954 => "00100101",18955 => "01010100",18956 => "00100110",18957 => "11010101",18958 => "01111000",18959 => "10100011",18960 => "00010010",18961 => "01101011",18962 => "00100010",18963 => "10000110",18964 => "11111000",18965 => "10110111",18966 => "11100010",18967 => "11001011",18968 => "10100101",18969 => "10010000",18970 => "01101011",18971 => "01001101",18972 => "10010100",18973 => "01001001",18974 => "10100011",18975 => "11101110",18976 => "01010011",18977 => "01111001",18978 => "10000100",18979 => "01000110",18980 => "01101101",18981 => "10110110",18982 => "01000010",18983 => "00110101",18984 => "10010010",18985 => "00001100",18986 => "00111100",18987 => "00100101",18988 => "11111110",18989 => "11100011",18990 => "11110001",18991 => "11100001",18992 => "11100001",18993 => "10101101",18994 => "10110100",18995 => "10111111",18996 => "11001101",18997 => "01111100",18998 => "00101111",18999 => "10000111",19000 => "00101111",19001 => "10110101",19002 => "11010110",19003 => "10000100",19004 => "01011011",19005 => "01100100",19006 => "10000111",19007 => "11010000",19008 => "11110110",19009 => "10010010",19010 => "10110100",19011 => "01001000",19012 => "01011011",19013 => "10100110",19014 => "01101110",19015 => "00110010",19016 => "11001100",19017 => "11000011",19018 => "01011010",19019 => "11111100",19020 => "00110111",19021 => "00010101",19022 => "00000001",19023 => "00111100",19024 => "00110101",19025 => "01010100",19026 => "00001110",19027 => "01101000",19028 => "11010010",19029 => "11001110",19030 => "11110000",19031 => "00111101",19032 => "10111000",19033 => "11110001",19034 => "11010010",19035 => "11111110",19036 => "11011111",19037 => "11100010",19038 => "01101110",19039 => "01100101",19040 => "10101101",19041 => "00111100",19042 => "11000101",19043 => "00011000",19044 => "01110110",19045 => "11110100",19046 => "10001101",19047 => "01110011",19048 => "10000000",19049 => "01011100",19050 => "10101010",19051 => "10111110",19052 => "01111100",19053 => "00011110",19054 => "00110001",19055 => "00001000",19056 => "10011011",19057 => "00110001",19058 => "01010111",19059 => "10111000",19060 => "01010000",19061 => "11100011",19062 => "10110011",19063 => "00001101",19064 => "01001101",19065 => "01100111",19066 => "11010111",19067 => "11000100",19068 => "11001001",19069 => "10010111",19070 => "10001100",19071 => "00110000",19072 => "10001010",19073 => "01011011",19074 => "10010101",19075 => "10000101",19076 => "00110010",19077 => "00010000",19078 => "11110101",19079 => "00100100",19080 => "01100010",19081 => "00011011",19082 => "01001011",19083 => "00100000",19084 => "10111111",19085 => "10110000",19086 => "01010111",19087 => "10011110",19088 => "11000110",19089 => "00101101",19090 => "00110000",19091 => "10001010",19092 => "11111101",19093 => "11010011",19094 => "01011111",19095 => "00001001",19096 => "10000101",19097 => "01100100",19098 => "00010110",19099 => "11010110",19100 => "00101110",19101 => "01001001",19102 => "11100010",19103 => "11001000",19104 => "01110100",19105 => "10000010",19106 => "10011011",19107 => "10010110",19108 => "10001110",19109 => "00110010",19110 => "11100010",19111 => "11010100",19112 => "00010111",19113 => "11101011",19114 => "11110011",19115 => "01000011",19116 => "10110101",19117 => "10101000",19118 => "11101100",19119 => "01000001",19120 => "00000110",19121 => "00111000",19122 => "00001110",19123 => "10000100",19124 => "00110110",19125 => "01000001",19126 => "00001010",19127 => "01101010",19128 => "00111001",19129 => "11010101",19130 => "01111011",19131 => "01101101",19132 => "01001010",19133 => "10010101",19134 => "10110111",19135 => "00101101",19136 => "11111100",19137 => "00110100",19138 => "11101000",19139 => "00100101",19140 => "11110110",19141 => "11100111",19142 => "00101011",19143 => "11011101",19144 => "01000010",19145 => "00100000",19146 => "11110010",19147 => "01101010",19148 => "10101110",19149 => "00010000",19150 => "00110010",19151 => "11101110",19152 => "01111100",19153 => "00101110",19154 => "11011011",19155 => "01111000",19156 => "10101000",19157 => "11111110",19158 => "11100110",19159 => "01011111",19160 => "10011101",19161 => "01011011",19162 => "10111101",19163 => "10111011",19164 => "01011110",19165 => "01111011",19166 => "10111001",19167 => "00100000",19168 => "01000001",19169 => "00110110",19170 => "01101101",19171 => "01111000",19172 => "11110011",19173 => "00001010",19174 => "00111000",19175 => "00100101",19176 => "00110001",19177 => "10011101",19178 => "11000100",19179 => "00011100",19180 => "10000111",19181 => "01001110",19182 => "11100100",19183 => "10000010",19184 => "10000011",19185 => "00010000",19186 => "10010000",19187 => "00000110",19188 => "11011101",19189 => "00111010",19190 => "11111100",19191 => "10111100",19192 => "00010010",19193 => "10100100",19194 => "10111001",19195 => "11001001",19196 => "00100000",19197 => "01001000",19198 => "10010001",19199 => "01010010",19200 => "01000101",19201 => "10100101",19202 => "00101011",19203 => "00111011",19204 => "10101100",19205 => "01100110",19206 => "11000001",19207 => "01001111",19208 => "01101011",19209 => "01100101",19210 => "10011010",19211 => "01110111",19212 => "00001001",19213 => "10000001",19214 => "10010100",19215 => "00011100",19216 => "10110110",19217 => "11100100",19218 => "11001110",19219 => "10011011",19220 => "01011101",19221 => "01110010",19222 => "10010101",19223 => "11000001",19224 => "01111101",19225 => "00101110",19226 => "01100011",19227 => "01101101",19228 => "10100110",19229 => "11110011",19230 => "00101111",19231 => "10001000",19232 => "10101001",19233 => "10011011",19234 => "00010111",19235 => "00110010",19236 => "01011110",19237 => "11100110",19238 => "01011111",19239 => "10010111",19240 => "11101110",19241 => "10011100",19242 => "10000000",19243 => "01011110",19244 => "00111100",19245 => "10010011",19246 => "11010100",19247 => "11010001",19248 => "11001111",19249 => "10110010",19250 => "11010001",19251 => "00011010",19252 => "10100011",19253 => "11001010",19254 => "01101010",19255 => "01010101",19256 => "11110101",19257 => "11001010",19258 => "01000100",19259 => "10110110",19260 => "01011011",19261 => "11001111",19262 => "11010101",19263 => "11011010",19264 => "11101001",19265 => "11000110",19266 => "11101101",19267 => "00101011",19268 => "01011100",19269 => "00011110",19270 => "10100111",19271 => "11101001",19272 => "00000101",19273 => "01000110",19274 => "00101011",19275 => "10111011",19276 => "11111011",19277 => "00100000",19278 => "01110000",19279 => "01100100",19280 => "00110110",19281 => "00101001",19282 => "11011100",19283 => "01100101",19284 => "01101110",19285 => "10100010",19286 => "00101110",19287 => "10000100",19288 => "11111110",19289 => "10100011",19290 => "11001011",19291 => "10000111",19292 => "00000110",19293 => "11001100",19294 => "00000100",19295 => "11110110",19296 => "11110010",19297 => "00100111",19298 => "01101010",19299 => "00001101",19300 => "00111010",19301 => "01010101",19302 => "00111010",19303 => "00011011",19304 => "10101001",19305 => "01111110",19306 => "00110000",19307 => "00101010",19308 => "00100000",19309 => "10100000",19310 => "11110111",19311 => "10100011",19312 => "11110110",19313 => "11100000",19314 => "00111011",19315 => "00001100",19316 => "00000100",19317 => "00001111",19318 => "01111001",19319 => "11001101",19320 => "10110100",19321 => "11010001",19322 => "01100110",19323 => "00100011",19324 => "10011011",19325 => "10101001",19326 => "11110001",19327 => "11001010",19328 => "10011101",19329 => "01111101",19330 => "11111000",19331 => "00101101",19332 => "00000100",19333 => "01111100",19334 => "11100000",19335 => "11100000",19336 => "00010111",19337 => "00000101",19338 => "01000111",19339 => "01000100",19340 => "01011001",19341 => "11101101",19342 => "11010010",19343 => "10000110",19344 => "11010010",19345 => "01101100",19346 => "01110010",19347 => "01110101",19348 => "10010101",19349 => "10110001",19350 => "10010100",19351 => "01110010",19352 => "10010011",19353 => "00010000",19354 => "00010100",19355 => "00101001",19356 => "00110111",19357 => "00001111",19358 => "10110111",19359 => "01011101",19360 => "00101001",19361 => "00001001",19362 => "10110001",19363 => "01010100",19364 => "10101100",19365 => "11111010",19366 => "01110001",19367 => "11000101",19368 => "00101011",19369 => "11001111",19370 => "01110011",19371 => "00010000",19372 => "00000001",19373 => "00001100",19374 => "11101010",19375 => "00001010",19376 => "00110110",19377 => "00011100",19378 => "00100100",19379 => "10101100",19380 => "01101100",19381 => "00111001",19382 => "10000011",19383 => "10010000",19384 => "11101100",19385 => "11011100",19386 => "01110000",19387 => "01010011",19388 => "00110011",19389 => "10110110",19390 => "01110110",19391 => "00000101",19392 => "01001110",19393 => "00101010",19394 => "00011001",19395 => "11010101",19396 => "11010010",19397 => "11000101",19398 => "10000010",19399 => "10101011",19400 => "00010011",19401 => "11001011",19402 => "00101101",19403 => "01010101",19404 => "00111000",19405 => "10011110",19406 => "00111100",19407 => "01001000",19408 => "01000100",19409 => "10101101",19410 => "00111101",19411 => "00101111",19412 => "00110000",19413 => "01100101",19414 => "10010100",19415 => "11111001",19416 => "01110001",19417 => "10011001",19418 => "10111010",19419 => "10111011",19420 => "10011110",19421 => "10111001",19422 => "01110011",19423 => "11000100",19424 => "11000101",19425 => "10111110",19426 => "01111001",19427 => "00011000",19428 => "10101010",19429 => "00111110",19430 => "10111000",19431 => "11110010",19432 => "10010101",19433 => "10110101",19434 => "01100100",19435 => "01000010",19436 => "00101111",19437 => "10111001",19438 => "00101001",19439 => "00000000",19440 => "10111100",19441 => "01000000",19442 => "01111001",19443 => "00101000",19444 => "10010110",19445 => "01001100",19446 => "10100010",19447 => "00101000",19448 => "11111110",19449 => "00010111",19450 => "11110100",19451 => "01000100",19452 => "00111110",19453 => "11001111",19454 => "11001010",19455 => "01101000",19456 => "01100101",19457 => "01101000",19458 => "01101000",19459 => "11101001",19460 => "01111100",19461 => "11111010",19462 => "00011000",19463 => "10101100",19464 => "00101110",19465 => "11000010",19466 => "10000001",19467 => "00100001",19468 => "10111010",19469 => "10010000",19470 => "00101011",19471 => "00001000",19472 => "00100010",19473 => "01010000",19474 => "00111011",19475 => "01110011",19476 => "00010100",19477 => "10000111",19478 => "01010011",19479 => "10111000",19480 => "11110101",19481 => "00001100",19482 => "10100110",19483 => "00001011",19484 => "01101111",19485 => "01111010",19486 => "00010101",19487 => "11100000",19488 => "00001011",19489 => "00001100",19490 => "11000100",19491 => "11011001",19492 => "01101001",19493 => "00011010",19494 => "10111110",19495 => "10101000",19496 => "10011100",19497 => "00101010",19498 => "00101111",19499 => "01010011",19500 => "00011000",19501 => "00011011",19502 => "11111101",19503 => "01011001",19504 => "00111100",19505 => "00000010",19506 => "01000100",19507 => "00011000",19508 => "01011110",19509 => "00000011",19510 => "11011001",19511 => "11111101",19512 => "11001110",19513 => "00011001",19514 => "01001010",19515 => "10101011",19516 => "01001100",19517 => "00000100",19518 => "01011001",19519 => "00110011",19520 => "01110111",19521 => "01101010",19522 => "01001110",19523 => "00101100",19524 => "00101010",19525 => "11111011",19526 => "11111010",19527 => "11110110",19528 => "11010011",19529 => "11001010",19530 => "01110000",19531 => "10011011",19532 => "10010111",19533 => "01011001",19534 => "11100110",19535 => "00001011",19536 => "10110101",19537 => "01101101",19538 => "11101001",19539 => "01111011",19540 => "01010100",19541 => "10001101",19542 => "11111010",19543 => "10010000",19544 => "10111110",19545 => "01101011",19546 => "10010010",19547 => "10010000",19548 => "10111101",19549 => "10011100",19550 => "10011100",19551 => "01101111",19552 => "01111010",19553 => "11000010",19554 => "10011101",19555 => "11101111",19556 => "00111010",19557 => "01101011",19558 => "00111000",19559 => "10010101",19560 => "01010001",19561 => "10001000",19562 => "11011101",19563 => "01001010",19564 => "11001010",19565 => "00001011",19566 => "00010001",19567 => "10110010",19568 => "01010100",19569 => "10011010",19570 => "00011010",19571 => "00101111",19572 => "11000000",19573 => "10110100",19574 => "10101001",19575 => "10110001",19576 => "01000011",19577 => "00110011",19578 => "01111000",19579 => "01111101",19580 => "00010001",19581 => "01110111",19582 => "00100010",19583 => "00011101",19584 => "10010101",19585 => "01001111",19586 => "11110010",19587 => "01011001",19588 => "00011001",19589 => "00010111",19590 => "01101000",19591 => "11001111",19592 => "00111110",19593 => "00100101",19594 => "11110100",19595 => "00100010",19596 => "01111001",19597 => "00001001",19598 => "01000100",19599 => "00011101",19600 => "10000111",19601 => "01100111",19602 => "00111000",19603 => "11101101",19604 => "00110010",19605 => "01010100",19606 => "01010001",19607 => "00011101",19608 => "11011110",19609 => "11111100",19610 => "10101000",19611 => "10111101",19612 => "00111001",19613 => "11110110",19614 => "10110100",19615 => "11011111",19616 => "11100000",19617 => "11100001",19618 => "00101001",19619 => "01101111",19620 => "01011110",19621 => "01000011",19622 => "01001010",19623 => "11011100",19624 => "10111010",19625 => "11000110",19626 => "01000001",19627 => "00011011",19628 => "01001001",19629 => "00001000",19630 => "11101110",19631 => "01101110",19632 => "00001001",19633 => "11001111",19634 => "10010001",19635 => "00101100",19636 => "10000001",19637 => "11110001",19638 => "00001100",19639 => "10001001",19640 => "00110011",19641 => "11111010",19642 => "11110111",19643 => "00001111",19644 => "01100111",19645 => "10010111",19646 => "01001011",19647 => "01010101",19648 => "10000111",19649 => "00001011",19650 => "11000101",19651 => "01000101",19652 => "01101010",19653 => "01001001",19654 => "10001111",19655 => "10011101",19656 => "01011011",19657 => "10001010",19658 => "10100000",19659 => "00010001",19660 => "00100000",19661 => "11011000",19662 => "00110011",19663 => "01001101",19664 => "10101010",19665 => "00101010",19666 => "01111011",19667 => "10101010",19668 => "00010010",19669 => "01011010",19670 => "01011001",19671 => "10111011",19672 => "01011111",19673 => "00001101",19674 => "00111010",19675 => "11111000",19676 => "10010110",19677 => "01101111",19678 => "01011110",19679 => "11010100",19680 => "10101010",19681 => "01001100",19682 => "01011000",19683 => "01110011",19684 => "10010100",19685 => "01011011",19686 => "11011110",19687 => "01100101",19688 => "10000110",19689 => "11011111",19690 => "10101001",19691 => "10100001",19692 => "01001101",19693 => "00011000",19694 => "01001111",19695 => "01001000",19696 => "10010011",19697 => "11011010",19698 => "01000010",19699 => "01111011",19700 => "10100100",19701 => "11011100",19702 => "01111101",19703 => "01000111",19704 => "10101101",19705 => "00111111",19706 => "11010111",19707 => "10011100",19708 => "01101011",19709 => "11010100",19710 => "10111110",19711 => "11010011",19712 => "10010110",19713 => "10100001",19714 => "10000000",19715 => "00110100",19716 => "00011111",19717 => "00100110",19718 => "11000011",19719 => "00010010",19720 => "10111101",19721 => "10001011",19722 => "00110011",19723 => "10111100",19724 => "11100011",19725 => "10110110",19726 => "11011111",19727 => "01101101",19728 => "00001001",19729 => "00110010",19730 => "11000000",19731 => "01000101",19732 => "00000100",19733 => "01000011",19734 => "00111100",19735 => "01110000",19736 => "00010001",19737 => "10101111",19738 => "11000111",19739 => "00011100",19740 => "11000011",19741 => "00011001",19742 => "00011011",19743 => "10001111",19744 => "01111011",19745 => "00100010",19746 => "11101101",19747 => "01010000",19748 => "01010111",19749 => "11001111",19750 => "11100001",19751 => "01011011",19752 => "10001111",19753 => "01010000",19754 => "11111100",19755 => "11000010",19756 => "01000101",19757 => "11101001",19758 => "01011111",19759 => "00111101",19760 => "01011001",19761 => "10010110",19762 => "10101010",19763 => "10100001",19764 => "10011011",19765 => "11100110",19766 => "00011011",19767 => "11000000",19768 => "11001010",19769 => "10100110",19770 => "11010100",19771 => "01101001",19772 => "11110101",19773 => "11111010",19774 => "11011110",19775 => "11111110",19776 => "00000111",19777 => "00111100",19778 => "01001011",19779 => "10000110",19780 => "01111001",19781 => "01101010",19782 => "10001110",19783 => "00010000",19784 => "01000100",19785 => "10101100",19786 => "01001001",19787 => "11010101",19788 => "10111111",19789 => "11000101",19790 => "01000000",19791 => "01111011",19792 => "11000100",19793 => "11100011",19794 => "11001010",19795 => "10110101",19796 => "00101011",19797 => "00001001",19798 => "01100011",19799 => "11111000",19800 => "11001100",19801 => "01011100",19802 => "00101111",19803 => "01011011",19804 => "11010101",19805 => "10001111",19806 => "10001111",19807 => "10110100",19808 => "10101000",19809 => "01001001",19810 => "11100011",19811 => "01101011",19812 => "01111001",19813 => "00100000",19814 => "01110010",19815 => "11100011",19816 => "01001011",19817 => "11010101",19818 => "00110101",19819 => "00011100",19820 => "10001110",19821 => "00111101",19822 => "01001010",19823 => "00001111",19824 => "10001010",19825 => "10000001",19826 => "11111000",19827 => "00100110",19828 => "01010011",19829 => "11000001",19830 => "01101101",19831 => "11110001",19832 => "11110000",19833 => "11010100",19834 => "00011010",19835 => "10000100",19836 => "01110110",19837 => "10110101",19838 => "10000001",19839 => "01111011",19840 => "11010001",19841 => "00110000",19842 => "10001000",19843 => "01010110",19844 => "00110011",19845 => "00111111",19846 => "01010000",19847 => "10010010",19848 => "00101011",19849 => "01010010",19850 => "11000011",19851 => "10101010",19852 => "10101000",19853 => "10111000",19854 => "10111110",19855 => "00011101",19856 => "10111000",19857 => "00110000",19858 => "10011011",19859 => "01000100",19860 => "00011001",19861 => "00110101",19862 => "11001011",19863 => "10111110",19864 => "00011001",19865 => "00100010",19866 => "11110000",19867 => "11100010",19868 => "00111111",19869 => "00100000",19870 => "00001101",19871 => "11100001",19872 => "01111001",19873 => "00110011",19874 => "00000010",19875 => "11101011",19876 => "10000010",19877 => "00010101",19878 => "10110111",19879 => "11011011",19880 => "01101011",19881 => "11000110",19882 => "11011100",19883 => "10001011",19884 => "00001011",19885 => "11001111",19886 => "11110111",19887 => "01010111",19888 => "11101001",19889 => "10110000",19890 => "01000111",19891 => "11010100",19892 => "11011000",19893 => "01110011",19894 => "10011011",19895 => "00011011",19896 => "01110011",19897 => "00000010",19898 => "10001111",19899 => "00001000",19900 => "00100010",19901 => "11101100",19902 => "11110001",19903 => "00001110",19904 => "01111100",19905 => "01011011",19906 => "10011000",19907 => "11110110",19908 => "11010100",19909 => "01101011",19910 => "11100010",19911 => "11100100",19912 => "00001100",19913 => "00110000",19914 => "11000100",19915 => "10100011",19916 => "00100111",19917 => "10111010",19918 => "00011001",19919 => "01111000",19920 => "00110011",19921 => "00000110",19922 => "01001010",19923 => "11110000",19924 => "00110111",19925 => "11111101",19926 => "10111000",19927 => "10011011",19928 => "00010011",19929 => "00000001",19930 => "10000110",19931 => "10100010",19932 => "00100011",19933 => "10100110",19934 => "00000111",19935 => "01011001",19936 => "01001010",19937 => "00001011",19938 => "10111100",19939 => "00101010",19940 => "10110010",19941 => "00101110",19942 => "01111011",19943 => "11101110",19944 => "10010000",19945 => "10111000",19946 => "01110011",19947 => "01011100",19948 => "01111010",19949 => "11110111",19950 => "11001011",19951 => "10110000",19952 => "01100000",19953 => "10101000",19954 => "00001000",19955 => "00001001",19956 => "10011100",19957 => "00101011",19958 => "11001101",19959 => "01101100",19960 => "10010000",19961 => "11100010",19962 => "11000110",19963 => "11110100",19964 => "11101011",19965 => "00011001",19966 => "10101011",19967 => "11011101",19968 => "11100111",19969 => "00000010",19970 => "00010101",19971 => "00000010",19972 => "11101011",19973 => "00111110",19974 => "01100011",19975 => "11111100",19976 => "01100101",19977 => "10011010",19978 => "11100110",19979 => "01111111",19980 => "01110001",19981 => "11100101",19982 => "00011111",19983 => "01100010",19984 => "11001101",19985 => "11111101",19986 => "01011111",19987 => "10111000",19988 => "11010011",19989 => "10000001",19990 => "01101100",19991 => "01000000",19992 => "10011100",19993 => "01100111",19994 => "01101100",19995 => "10110001",19996 => "01000001",19997 => "10100011",19998 => "11001000",19999 => "00111010",20000 => "10001000",20001 => "10100101",20002 => "10101000",20003 => "01111010",20004 => "01101111",20005 => "00101011",20006 => "11000100",20007 => "10001101",20008 => "10001100",20009 => "01011000",20010 => "11110011",20011 => "11000100",20012 => "00011011",20013 => "01111100",20014 => "10111100",20015 => "11010110",20016 => "01101100",20017 => "00000011",20018 => "10101001",20019 => "11011100",20020 => "01001110",20021 => "00011011",20022 => "00010111",20023 => "01000111",20024 => "01000010",20025 => "10110011",20026 => "01010011",20027 => "00111100",20028 => "10000110",20029 => "01110011",20030 => "10010101",20031 => "01100001",20032 => "00010001",20033 => "01111000",20034 => "00110010",20035 => "00111001",20036 => "01110001",20037 => "11100110",20038 => "00000101",20039 => "01000011",20040 => "00111101",20041 => "11100110",20042 => "11100100",20043 => "01111010",20044 => "01100001",20045 => "10010001",20046 => "01111110",20047 => "10010111",20048 => "00000100",20049 => "00010000",20050 => "00000001",20051 => "01010010",20052 => "00111110",20053 => "10110110",20054 => "01000010",20055 => "11111011",20056 => "11001111",20057 => "11010110",20058 => "11001011",20059 => "10001000",20060 => "10000110",20061 => "01110101",20062 => "11011010",20063 => "10011011",20064 => "00001001",20065 => "01101001",20066 => "10111110",20067 => "10011111",20068 => "10101110",20069 => "11100111",20070 => "01000000",20071 => "10100011",20072 => "00010011",20073 => "00011011",20074 => "11010100",20075 => "01001011",20076 => "11111010",20077 => "11111111",20078 => "10011110",20079 => "00101110",20080 => "11111110",20081 => "00010010",20082 => "11111011",20083 => "11111000",20084 => "01010101",20085 => "01011011",20086 => "01000001",20087 => "00101111",20088 => "01111001",20089 => "00110011",20090 => "01101110",20091 => "11001010",20092 => "00011110",20093 => "10011011",20094 => "00000001",20095 => "01011001",20096 => "11001001",20097 => "11010001",20098 => "11001111",20099 => "01100010",20100 => "11100110",20101 => "01101111",20102 => "01100000",20103 => "11100111",20104 => "00100110",20105 => "11001100",20106 => "01011100",20107 => "01010000",20108 => "11001101",20109 => "01010010",20110 => "01010110",20111 => "11111111",20112 => "10110111",20113 => "11001111",20114 => "01101100",20115 => "00000010",20116 => "10011001",20117 => "10111010",20118 => "01111111",20119 => "11100101",20120 => "11101010",20121 => "10011010",20122 => "01001011",20123 => "01110101",20124 => "11101000",20125 => "11000000",20126 => "11001101",20127 => "00001101",20128 => "11110100",20129 => "10111100",20130 => "10111100",20131 => "01111101",20132 => "11101111",20133 => "10101110",20134 => "10101111",20135 => "11001100",20136 => "00101101",20137 => "01010001",20138 => "00110101",20139 => "00101110",20140 => "10011111",20141 => "11101011",20142 => "11001010",20143 => "00000100",20144 => "01011011",20145 => "01110101",20146 => "10010101",20147 => "00101111",20148 => "01101100",20149 => "10101011",20150 => "00101001",20151 => "10110011",20152 => "01100011",20153 => "11101011",20154 => "01101010",20155 => "11011011",20156 => "11010110",20157 => "00000000",20158 => "11100010",20159 => "11110000",20160 => "10100010",20161 => "11101000",20162 => "10001000",20163 => "10111101",20164 => "10001101",20165 => "11000001",20166 => "00001111",20167 => "01100001",20168 => "10010000",20169 => "11110001",20170 => "11000011",20171 => "00101010",20172 => "00110001",20173 => "11000001",20174 => "10101010",20175 => "10110100",20176 => "00101000",20177 => "11100011",20178 => "10000100",20179 => "11010010",20180 => "10011110",20181 => "01010100",20182 => "10010000",20183 => "00010111",20184 => "01000000",20185 => "11110000",20186 => "01001011",20187 => "00000100",20188 => "00100110",20189 => "10110011",20190 => "10111101",20191 => "11010010",20192 => "01111000",20193 => "10001001",20194 => "01011001",20195 => "11111011",20196 => "10111101",20197 => "01011001",20198 => "00000100",20199 => "11000110",20200 => "01111011",20201 => "11001101",20202 => "00101101",20203 => "00110100",20204 => "01110011",20205 => "00110101",20206 => "10100110",20207 => "11101000",20208 => "01110011",20209 => "10011011",20210 => "00100100",20211 => "00011101",20212 => "00110000",20213 => "11101000",20214 => "00011101",20215 => "11001011",20216 => "11011110",20217 => "01010011",20218 => "00100111",20219 => "11010010",20220 => "11101101",20221 => "01001010",20222 => "11001100",20223 => "00010100",20224 => "01000000",20225 => "00101010",20226 => "00101011",20227 => "11100100",20228 => "01011110",20229 => "10010011",20230 => "00011001",20231 => "11110000",20232 => "00000000",20233 => "11001001",20234 => "01000010",20235 => "00000110",20236 => "01111010",20237 => "10101011",20238 => "10100101",20239 => "11000111",20240 => "00101010",20241 => "01101100",20242 => "01000010",20243 => "01001100",20244 => "01001000",20245 => "00111100",20246 => "01010010",20247 => "00111001",20248 => "10001101",20249 => "10100001",20250 => "11111111",20251 => "11101000",20252 => "00010111",20253 => "11111101",20254 => "10101101",20255 => "10101111",20256 => "00001001",20257 => "11010010",20258 => "01011000",20259 => "11000111",20260 => "10001011",20261 => "01001001",20262 => "11111100",20263 => "00111000",20264 => "10001000",20265 => "11101100",20266 => "11101101",20267 => "01101011",20268 => "11100011",20269 => "11010000",20270 => "10100011",20271 => "11011100",20272 => "10010100",20273 => "01101010",20274 => "00000111",20275 => "01010100",20276 => "01111001",20277 => "10000000",20278 => "10101000",20279 => "11000110",20280 => "10011101",20281 => "00110010",20282 => "00110110",20283 => "10111000",20284 => "00001001",20285 => "00010110",20286 => "10100010",20287 => "11000011",20288 => "00100010",20289 => "10010100",20290 => "11100111",20291 => "10110000",20292 => "11101100",20293 => "10100001",20294 => "10101111",20295 => "00111001",20296 => "01110001",20297 => "10001100",20298 => "00100011",20299 => "10000111",20300 => "01000101",20301 => "00000101",20302 => "01001110",20303 => "01010110",20304 => "10011000",20305 => "10110100",20306 => "10000111",20307 => "11111001",20308 => "10000111",20309 => "01000101",20310 => "01000110",20311 => "00110101",20312 => "00010100",20313 => "00001001",20314 => "10001001",20315 => "01000001",20316 => "01110110",20317 => "00010110",20318 => "10011010",20319 => "01100010",20320 => "11111110",20321 => "01110000",20322 => "00000010",20323 => "01110100",20324 => "00010011",20325 => "11011001",20326 => "01000011",20327 => "10110000",20328 => "01100111",20329 => "11011111",20330 => "10010001",20331 => "01110101",20332 => "11010011",20333 => "10101001",20334 => "01111011",20335 => "01011100",20336 => "10111100",20337 => "10100001",20338 => "01111100",20339 => "00110000",20340 => "10110010",20341 => "01100111",20342 => "10000100",20343 => "10100010",20344 => "10000110",20345 => "00100110",20346 => "10011010",20347 => "10101001",20348 => "01101110",20349 => "00010001",20350 => "00111110",20351 => "00001100",20352 => "00001000",20353 => "01010110",20354 => "01011000",20355 => "10110111",20356 => "11111110",20357 => "01111111",20358 => "01111110",20359 => "10001000",20360 => "10100100",20361 => "10000010",20362 => "10101011",20363 => "10100101",20364 => "11011110",20365 => "00011100",20366 => "10010010",20367 => "00101010",20368 => "11010010",20369 => "00001101",20370 => "01011111",20371 => "10111001",20372 => "01101111",20373 => "01011000",20374 => "10001000",20375 => "10110000",20376 => "00011010",20377 => "11100101",20378 => "00000001",20379 => "00101001",20380 => "00010101",20381 => "11011100",20382 => "10111010",20383 => "00001101",20384 => "10110100",20385 => "11010100",20386 => "00010011",20387 => "10101101",20388 => "01000001",20389 => "11000100",20390 => "10110010",20391 => "00011101",20392 => "01101011",20393 => "11010110",20394 => "11100000",20395 => "01101001",20396 => "11101100",20397 => "10000010",20398 => "00111010",20399 => "00111011",20400 => "01011001",20401 => "11100110",20402 => "01001101",20403 => "00001110",20404 => "00101101",20405 => "00010101",20406 => "00000111",20407 => "10001010",20408 => "01111111",20409 => "00010011",20410 => "11101101",20411 => "00110001",20412 => "11110001",20413 => "01111001",20414 => "01111101",20415 => "11100100",20416 => "01001000",20417 => "00101001",20418 => "01110111",20419 => "01101010",20420 => "00111110",20421 => "01101100",20422 => "10010011",20423 => "00000001",20424 => "11110011",20425 => "10010010",20426 => "11111001",20427 => "11110000",20428 => "01111000",20429 => "11000001",20430 => "00111100",20431 => "01100000",20432 => "00111010",20433 => "10110001",20434 => "10101010",20435 => "10001001",20436 => "10001110",20437 => "00101111",20438 => "00001010",20439 => "11010101",20440 => "10010001",20441 => "01001001",20442 => "10101111",20443 => "10010010",20444 => "01100110",20445 => "01011101",20446 => "00010111",20447 => "11011010",20448 => "11010100",20449 => "00100101",20450 => "01001110",20451 => "01011010",20452 => "00111001",20453 => "10011111",20454 => "01010110",20455 => "11101111",20456 => "10101011",20457 => "11011101",20458 => "10010101",20459 => "01001111",20460 => "11011110",20461 => "00011010",20462 => "11111110",20463 => "01011101",20464 => "10011101",20465 => "11111000",20466 => "11100101",20467 => "11010000",20468 => "11101100",20469 => "10010100",20470 => "10110011",20471 => "10010000",20472 => "11010111",20473 => "00111010",20474 => "01001111",20475 => "10111100",20476 => "10001101",20477 => "11111011",20478 => "10000111",20479 => "10010110",20480 => "10010010",20481 => "00000001",20482 => "11011010",20483 => "10110000",20484 => "10000011",20485 => "10101110",20486 => "00110011",20487 => "01010101",20488 => "00100001",20489 => "11011001",20490 => "11001100",20491 => "00100011",20492 => "01000110",20493 => "10000101",20494 => "00111100",20495 => "10011101",20496 => "01100101",20497 => "01111111",20498 => "01100110",20499 => "10101101",20500 => "11110001",20501 => "11010001",20502 => "10001011",20503 => "01010010",20504 => "00000000",20505 => "01101010",20506 => "00001100",20507 => "00101010",20508 => "01011000",20509 => "10101000",20510 => "11101001",20511 => "00011011",20512 => "11100111",20513 => "10000110",20514 => "01100011",20515 => "11111001",20516 => "10011110",20517 => "01111011",20518 => "11001000",20519 => "01110100",20520 => "00110010",20521 => "11011111",20522 => "00101010",20523 => "00100010",20524 => "01110110",20525 => "01010010",20526 => "11010100",20527 => "11110001",20528 => "11011010",20529 => "00010010",20530 => "01011101",20531 => "01111001",20532 => "01000000",20533 => "11111010",20534 => "11010010",20535 => "11011100",20536 => "01001001",20537 => "11111000",20538 => "01010001",20539 => "00010100",20540 => "11101000",20541 => "11001111",20542 => "11110011",20543 => "11110111",20544 => "10010011",20545 => "11010110",20546 => "10101001",20547 => "00110100",20548 => "11100011",20549 => "11000111",20550 => "11100010",20551 => "10011001",20552 => "11010000",20553 => "00001111",20554 => "00001100",20555 => "00000101",20556 => "11110100",20557 => "01000101",20558 => "10100100",20559 => "10010000",20560 => "00010110",20561 => "00000100",20562 => "01101000",20563 => "11010101",20564 => "00110100",20565 => "10101101",20566 => "00101001",20567 => "10001100",20568 => "10101011",20569 => "10000100",20570 => "10100111",20571 => "10110001",20572 => "00000101",20573 => "11011100",20574 => "10010011",20575 => "01110001",20576 => "00100101",20577 => "10111001",20578 => "10011000",20579 => "00100101",20580 => "00111011",20581 => "01110011",20582 => "11011101",20583 => "11100000",20584 => "00101001",20585 => "01111110",20586 => "11001010",20587 => "01000110",20588 => "01000110",20589 => "10111001",20590 => "01001110",20591 => "01111101",20592 => "10001010",20593 => "01101000",20594 => "01101101",20595 => "11011001",20596 => "00011011",20597 => "00110100",20598 => "00011110",20599 => "00101001",20600 => "10010011",20601 => "11111011",20602 => "01001000",20603 => "00100011",20604 => "00101110",20605 => "11111000",20606 => "01001101",20607 => "01011111",20608 => "10010110",20609 => "00000110",20610 => "00001011",20611 => "10011101",20612 => "10111010",20613 => "10111100",20614 => "00001100",20615 => "00010001",20616 => "10000011",20617 => "10100001",20618 => "11110100",20619 => "00010010",20620 => "01001100",20621 => "00011111",20622 => "01010100",20623 => "11110101",20624 => "01110101",20625 => "11101011",20626 => "00100011",20627 => "01110100",20628 => "00100100",20629 => "01010001",20630 => "01100000",20631 => "01010111",20632 => "11010111",20633 => "01001111",20634 => "01100101",20635 => "00001100",20636 => "11001001",20637 => "00010101",20638 => "10010000",20639 => "00101111",20640 => "10110110",20641 => "01010111",20642 => "00100011",20643 => "10001010",20644 => "01001111",20645 => "00010110",20646 => "00110101",20647 => "01001001",20648 => "01110101",20649 => "00110100",20650 => "00001111",20651 => "11100001",20652 => "00111000",20653 => "10010101",20654 => "00000010",20655 => "01011000",20656 => "00011011",20657 => "11110100",20658 => "01110001",20659 => "00000100",20660 => "01111011",20661 => "01010111",20662 => "11110101",20663 => "01000001",20664 => "11001111",20665 => "10010001",20666 => "00001100",20667 => "00101101",20668 => "11111110",20669 => "01100001",20670 => "10000100",20671 => "11010100",20672 => "10010010",20673 => "00110010",20674 => "00101111",20675 => "10010100",20676 => "11000001",20677 => "00111000",20678 => "01000011",20679 => "01011010",20680 => "00110010",20681 => "11100110",20682 => "10111000",20683 => "00100000",20684 => "10101111",20685 => "11110111",20686 => "11011011",20687 => "11110100",20688 => "00100011",20689 => "10111000",20690 => "10000101",20691 => "10010011",20692 => "00101011",20693 => "00001001",20694 => "11011110",20695 => "10011110",20696 => "01001000",20697 => "00000101",20698 => "10100100",20699 => "01101110",20700 => "01001111",20701 => "11111110",20702 => "11001100",20703 => "11000101",20704 => "11011110",20705 => "11000001",20706 => "01011011",20707 => "10100010",20708 => "11011010",20709 => "10110111",20710 => "01011001",20711 => "00110101",20712 => "11110000",20713 => "00101010",20714 => "11000011",20715 => "11011101",20716 => "01110000",20717 => "01101100",20718 => "00011010",20719 => "11011001",20720 => "10010001",20721 => "00101111",20722 => "00000100",20723 => "10110101",20724 => "00110000",20725 => "00111101",20726 => "01010111",20727 => "11001110",20728 => "11011001",20729 => "01111000",20730 => "11010010",20731 => "00001111",20732 => "01011001",20733 => "01000011",20734 => "10101100",20735 => "11111100",20736 => "01001000",20737 => "01011001",20738 => "01001100",20739 => "00001011",20740 => "11000010",20741 => "00110110",20742 => "00000011",20743 => "11110101",20744 => "00101100",20745 => "01010010",20746 => "11001100",20747 => "00001000",20748 => "00101001",20749 => "10000110",20750 => "01100000",20751 => "00000111",20752 => "01101010",20753 => "10001101",20754 => "10100001",20755 => "01111000",20756 => "00110111",20757 => "11101111",20758 => "00101101",20759 => "00000010",20760 => "01100101",20761 => "11001100",20762 => "11010001",20763 => "10110100",20764 => "11111001",20765 => "10000100",20766 => "10100001",20767 => "01001101",20768 => "11010111",20769 => "00010011",20770 => "11110111",20771 => "00000011",20772 => "01101100",20773 => "10110000",20774 => "01000101",20775 => "11000000",20776 => "10010010",20777 => "11111100",20778 => "11100000",20779 => "11011100",20780 => "11101010",20781 => "00101010",20782 => "11110101",20783 => "10000101",20784 => "01110000",20785 => "11010110",20786 => "00000001",20787 => "00110100",20788 => "00101101",20789 => "10111100",20790 => "00011100",20791 => "00110101",20792 => "00000101",20793 => "11111001",20794 => "01000110",20795 => "10010011",20796 => "00110111",20797 => "00001000",20798 => "00101110",20799 => "10011111",20800 => "11000111",20801 => "11111111",20802 => "10111110",20803 => "00101000",20804 => "10010110",20805 => "10100110",20806 => "11010000",20807 => "11000001",20808 => "10011111",20809 => "01010001",20810 => "00101001",20811 => "00000110",20812 => "11100101",20813 => "10111101",20814 => "00010111",20815 => "01101110",20816 => "00001101",20817 => "10101110",20818 => "11000110",20819 => "11001001",20820 => "10011110",20821 => "11011110",20822 => "11101101",20823 => "00000001",20824 => "01011110",20825 => "01100111",20826 => "00110010",20827 => "01001110",20828 => "01101011",20829 => "01010101",20830 => "10110100",20831 => "11001001",20832 => "11000010",20833 => "10000000",20834 => "01111000",20835 => "00000100",20836 => "11001010",20837 => "10100000",20838 => "01010000",20839 => "00000001",20840 => "11101101",20841 => "01111111",20842 => "10011000",20843 => "11010110",20844 => "01100100",20845 => "10111010",20846 => "10010110",20847 => "11100100",20848 => "11111011",20849 => "00000110",20850 => "00101101",20851 => "11111011",20852 => "00111001",20853 => "10111000",20854 => "01111000",20855 => "01111101",20856 => "00100001",20857 => "11011001",20858 => "11111111",20859 => "10100110",20860 => "00110011",20861 => "11111110",20862 => "10010001",20863 => "10011000",20864 => "11110101",20865 => "00101111",20866 => "10001000",20867 => "11011110",20868 => "10010101",20869 => "10111100",20870 => "10000111",20871 => "11011110",20872 => "10111011",20873 => "11000001",20874 => "10111110",20875 => "00110110",20876 => "01100010",20877 => "00111101",20878 => "10000100",20879 => "11111011",20880 => "10111000",20881 => "00010100",20882 => "01011100",20883 => "10100011",20884 => "01100001",20885 => "00101010",20886 => "01101111",20887 => "10111000",20888 => "11100011",20889 => "10010010",20890 => "00010010",20891 => "00011110",20892 => "10100001",20893 => "00101010",20894 => "00010000",20895 => "10110010",20896 => "11100010",20897 => "11110010",20898 => "01000100",20899 => "10110011",20900 => "00111110",20901 => "11110000",20902 => "11100101",20903 => "10010011",20904 => "00110100",20905 => "10000100",20906 => "11101001",20907 => "10100110",20908 => "10010110",20909 => "01100101",20910 => "00000110",20911 => "01100001",20912 => "11110100",20913 => "00000001",20914 => "10111111",20915 => "11111101",20916 => "00001111",20917 => "00011001",20918 => "00010000",20919 => "10100000",20920 => "11000100",20921 => "01101010",20922 => "01010100",20923 => "11001110",20924 => "11001101",20925 => "10101110",20926 => "10111011",20927 => "10110000",20928 => "00011110",20929 => "10100000",20930 => "10101110",20931 => "10011000",20932 => "01110100",20933 => "00110001",20934 => "00000111",20935 => "00011111",20936 => "00011110",20937 => "01001100",20938 => "10010001",20939 => "01111101",20940 => "01111111",20941 => "01001001",20942 => "11110110",20943 => "10100011",20944 => "00100111",20945 => "00001001",20946 => "00101100",20947 => "10101011",20948 => "10001100",20949 => "11111011",20950 => "01110110",20951 => "11110110",20952 => "00001010",20953 => "11001111",20954 => "10110100",20955 => "00000011",20956 => "10010011",20957 => "01100101",20958 => "01010001",20959 => "10000110",20960 => "01011001",20961 => "11000000",20962 => "10000011",20963 => "00011110",20964 => "10101011",20965 => "11101101",20966 => "11100101",20967 => "11110110",20968 => "00111100",20969 => "00011011",20970 => "10101101",20971 => "00010011",20972 => "01011001",20973 => "11000011",20974 => "10100000",20975 => "10001010",20976 => "00010100",20977 => "01000001",20978 => "01000111",20979 => "10111101",20980 => "00000110",20981 => "10010110",20982 => "11011011",20983 => "00111010",20984 => "10011101",20985 => "10001110",20986 => "10001000",20987 => "00111111",20988 => "00000110",20989 => "00110001",20990 => "00001011",20991 => "11101001",20992 => "11100011",20993 => "10010110",20994 => "00011000",20995 => "00100000",20996 => "01000010",20997 => "10110110",20998 => "10001010",20999 => "01110010",21000 => "00001101",21001 => "00100101",21002 => "00101000",21003 => "10010111",21004 => "11010010",21005 => "11101110",21006 => "11111011",21007 => "10110100",21008 => "11101011",21009 => "00010000",21010 => "00001111",21011 => "00100111",21012 => "10001011",21013 => "01011000",21014 => "10001100",21015 => "00111100",21016 => "01110011",21017 => "11100011",21018 => "10110010",21019 => "10111010",21020 => "11100001",21021 => "01100000",21022 => "01010101",21023 => "01001101",21024 => "10101110",21025 => "01011010",21026 => "11001111",21027 => "10011111",21028 => "00110000",21029 => "10101111",21030 => "10101111",21031 => "10111110",21032 => "11111110",21033 => "00000111",21034 => "11110110",21035 => "00011101",21036 => "01111100",21037 => "01000111",21038 => "01110100",21039 => "11000011",21040 => "10001011",21041 => "10000110",21042 => "11010001",21043 => "00010110",21044 => "01110000",21045 => "11111011",21046 => "10001001",21047 => "00010100",21048 => "11111000",21049 => "00110000",21050 => "01011011",21051 => "01101110",21052 => "01001101",21053 => "11101011",21054 => "01101100",21055 => "10101100",21056 => "01100110",21057 => "11000000",21058 => "00000011",21059 => "11010101",21060 => "01011011",21061 => "10110010",21062 => "11011000",21063 => "00101011",21064 => "01001001",21065 => "11011010",21066 => "00110101",21067 => "01111100",21068 => "10110010",21069 => "00110111",21070 => "00100010",21071 => "01101001",21072 => "00101011",21073 => "00011001",21074 => "00101000",21075 => "10000000",21076 => "11110110",21077 => "01010111",21078 => "10111001",21079 => "10000111",21080 => "01010000",21081 => "10000000",21082 => "11011010",21083 => "10011101",21084 => "00111110",21085 => "00110110",21086 => "00100101",21087 => "10001110",21088 => "00110000",21089 => "11110101",21090 => "01111111",21091 => "11100001",21092 => "10101001",21093 => "01000011",21094 => "10001011",21095 => "11110000",21096 => "11111100",21097 => "00111000",21098 => "10101111",21099 => "11011010",21100 => "10111011",21101 => "10111000",21102 => "01100001",21103 => "01010101",21104 => "11101111",21105 => "01011100",21106 => "11101001",21107 => "11000111",21108 => "11000101",21109 => "01100110",21110 => "01111101",21111 => "00111011",21112 => "10010101",21113 => "11011101",21114 => "01110011",21115 => "00000100",21116 => "11010100",21117 => "01101011",21118 => "01001010",21119 => "11000010",21120 => "01001000",21121 => "01100100",21122 => "01001111",21123 => "01101110",21124 => "01001000",21125 => "00001110",21126 => "00000110",21127 => "00100010",21128 => "11001010",21129 => "00111111",21130 => "10000101",21131 => "00000111",21132 => "10010110",21133 => "00100000",21134 => "10000110",21135 => "10111001",21136 => "10010110",21137 => "10100011",21138 => "10000000",21139 => "10110110",21140 => "10101111",21141 => "11011001",21142 => "11000010",21143 => "11011101",21144 => "00001001",21145 => "00001001",21146 => "00110110",21147 => "01011001",21148 => "10011011",21149 => "00001100",21150 => "10000011",21151 => "01111000",21152 => "11101001",21153 => "10000010",21154 => "11100100",21155 => "11000101",21156 => "10111111",21157 => "10101111",21158 => "00110001",21159 => "00001000",21160 => "00101110",21161 => "11111011",21162 => "01000011",21163 => "11110101",21164 => "01001010",21165 => "00101110",21166 => "10111110",21167 => "11100111",21168 => "01010010",21169 => "00101011",21170 => "00110000",21171 => "01001001",21172 => "01101011",21173 => "00001011",21174 => "11101111",21175 => "01101100",21176 => "11100110",21177 => "10101100",21178 => "00100001",21179 => "11111110",21180 => "11110000",21181 => "11010101",21182 => "01011000",21183 => "00000101",21184 => "01011000",21185 => "01100000",21186 => "10010111",21187 => "01100110",21188 => "01111011",21189 => "01100101",21190 => "11111100",21191 => "10001110",21192 => "11010011",21193 => "01100001",21194 => "10111111",21195 => "00011100",21196 => "10001011",21197 => "11111011",21198 => "01101001",21199 => "11000010",21200 => "01010100",21201 => "01000000",21202 => "01101000",21203 => "10011011",21204 => "10100000",21205 => "10000110",21206 => "01110000",21207 => "01100101",21208 => "01100100",21209 => "01010000",21210 => "01110110",21211 => "00101111",21212 => "01000101",21213 => "10110100",21214 => "11011000",21215 => "10110100",21216 => "00010010",21217 => "00111001",21218 => "01101111",21219 => "00110110",21220 => "10010100",21221 => "00000000",21222 => "01001101",21223 => "10101110",21224 => "01111010",21225 => "10101010",21226 => "01011101",21227 => "11110001",21228 => "10100001",21229 => "01000011",21230 => "11111101",21231 => "01110000",21232 => "10010111",21233 => "00011010",21234 => "11100011",21235 => "10110101",21236 => "01010011",21237 => "11101010",21238 => "10111111",21239 => "11111111",21240 => "11011111",21241 => "10100101",21242 => "01100000",21243 => "10110100",21244 => "00101010",21245 => "11101000",21246 => "10110001",21247 => "10111110",21248 => "11100010",21249 => "10001010",21250 => "11111111",21251 => "11011100",21252 => "00000001",21253 => "10001001",21254 => "01100110",21255 => "10110010",21256 => "01000111",21257 => "11001000",21258 => "11110111",21259 => "11110000",21260 => "10010010",21261 => "11101110",21262 => "00110011",21263 => "00010011",21264 => "00001011",21265 => "01000100",21266 => "11101111",21267 => "01110100",21268 => "00000001",21269 => "11011110",21270 => "01100011",21271 => "00111000",21272 => "10001101",21273 => "00000010",21274 => "01101110",21275 => "11010110",21276 => "00110101",21277 => "11001111",21278 => "11110010",21279 => "00101110",21280 => "01101010",21281 => "11010111",21282 => "01000111",21283 => "11100011",21284 => "11110001",21285 => "00100110",21286 => "00001101",21287 => "00001001",21288 => "00011000",21289 => "10111010",21290 => "00000100",21291 => "01101010",21292 => "00111101",21293 => "00010010",21294 => "11100001",21295 => "11110000",21296 => "10000000",21297 => "01110111",21298 => "10100011",21299 => "01100100",21300 => "11011111",21301 => "01001101",21302 => "11110111",21303 => "11100010",21304 => "00100110",21305 => "11011111",21306 => "00001101",21307 => "10100111",21308 => "01100001",21309 => "10011010",21310 => "01001000",21311 => "10001110",21312 => "00011100",21313 => "11001011",21314 => "11010111",21315 => "11110111",21316 => "00111100",21317 => "00111111",21318 => "00010011",21319 => "10010101",21320 => "01001001",21321 => "00101011",21322 => "10001111",21323 => "01100010",21324 => "00001100",21325 => "11001110",21326 => "01101100",21327 => "01010111",21328 => "10110110",21329 => "11110110",21330 => "10010111",21331 => "00101111",21332 => "01100011",21333 => "11111100",21334 => "00101100",21335 => "11100010",21336 => "11100100",21337 => "01111011",21338 => "00011100",21339 => "01101101",21340 => "10011010",21341 => "10011001",21342 => "01000000",21343 => "10110000",21344 => "11111110",21345 => "11010100",21346 => "00001100",21347 => "00101010",21348 => "00101101",21349 => "01110110",21350 => "00001111",21351 => "00001110",21352 => "01010001",21353 => "00001111",21354 => "10110100",21355 => "11110000",21356 => "11100010",21357 => "10111010",21358 => "10111010",21359 => "10010110",21360 => "00000001",21361 => "11100000",21362 => "00001101",21363 => "01101011",21364 => "00111011",21365 => "11110100",21366 => "11101010",21367 => "00111010",21368 => "00101010",21369 => "10111100",21370 => "10110010",21371 => "11001011",21372 => "00000100",21373 => "00110111",21374 => "10100010",21375 => "00100010",21376 => "00110010",21377 => "10000111",21378 => "11000001",21379 => "01101100",21380 => "01000011",21381 => "00011000",21382 => "11101111",21383 => "01000111",21384 => "00010111",21385 => "00011100",21386 => "10001011",21387 => "00001001",21388 => "11110100",21389 => "00011111",21390 => "00011101",21391 => "01110101",21392 => "10011001",21393 => "10111100",21394 => "11111001",21395 => "11100011",21396 => "11011000",21397 => "01101110",21398 => "01000101",21399 => "01100110",21400 => "10001000",21401 => "00110001",21402 => "11110011",21403 => "01001100",21404 => "10010100",21405 => "11101011",21406 => "00101001",21407 => "00111000",21408 => "01011001",21409 => "10110111",21410 => "01001101",21411 => "10000100",21412 => "10101011",21413 => "00010011",21414 => "11110101",21415 => "10111100",21416 => "00111110",21417 => "01000000",21418 => "01001011",21419 => "10001000",21420 => "10111101",21421 => "00111000",21422 => "11111100",21423 => "01110111",21424 => "01001111",21425 => "11000000",21426 => "10010001",21427 => "01011110",21428 => "00010101",21429 => "10101111",21430 => "00100111",21431 => "10100000",21432 => "01100010",21433 => "11110010",21434 => "01010110",21435 => "01011100",21436 => "00000001",21437 => "10110111",21438 => "01010101",21439 => "00111101",21440 => "11011100",21441 => "10001100",21442 => "10011100",21443 => "10001111",21444 => "11011100",21445 => "00011010",21446 => "10110111",21447 => "00000101",21448 => "00101010",21449 => "10000011",21450 => "01100001",21451 => "10010100",21452 => "01100011",21453 => "01000111",21454 => "01000111",21455 => "11010001",21456 => "11101010",21457 => "11001010",21458 => "10101000",21459 => "10001110",21460 => "01101110",21461 => "01011001",21462 => "01100010",21463 => "00111001",21464 => "00001011",21465 => "10010000",21466 => "11110001",21467 => "10011110",21468 => "01000000",21469 => "10101101",21470 => "01100000",21471 => "01000100",21472 => "01001111",21473 => "11001000",21474 => "01101100",21475 => "00001101",21476 => "01000100",21477 => "00111010",21478 => "00101110",21479 => "01010000",21480 => "01000100",21481 => "01100001",21482 => "00100100",21483 => "00000100",21484 => "00111011",21485 => "00011100",21486 => "10011000",21487 => "11010001",21488 => "11110101",21489 => "10001000",21490 => "11000111",21491 => "00001011",21492 => "00001110",21493 => "11001100",21494 => "10011100",21495 => "00101000",21496 => "10100010",21497 => "11010000",21498 => "10001111",21499 => "00010001",21500 => "11011100",21501 => "10001110",21502 => "11110001",21503 => "11100010",21504 => "00100110",21505 => "01100110",21506 => "01110111",21507 => "11000101",21508 => "01011011",21509 => "01111000",21510 => "11101110",21511 => "11011111",21512 => "01100110",21513 => "01101001",21514 => "00101100",21515 => "00000100",21516 => "11011011",21517 => "00100010",21518 => "00010101",21519 => "00000110",21520 => "11011000",21521 => "00111010",21522 => "00111001",21523 => "00011110",21524 => "10111001",21525 => "10000001",21526 => "10101001",21527 => "10111110",21528 => "11100100",21529 => "00111100",21530 => "00100001",21531 => "01100111",21532 => "11010010",21533 => "00011110",21534 => "00111011",21535 => "11100101",21536 => "10110010",21537 => "01000101",21538 => "00000101",21539 => "10011010",21540 => "10011110",21541 => "00110111",21542 => "00111111",21543 => "11111001",21544 => "01011000",21545 => "10111100",21546 => "11110000",21547 => "00000000",21548 => "10101010",21549 => "10011011",21550 => "00100011",21551 => "01000011",21552 => "11110001",21553 => "00110011",21554 => "11111100",21555 => "00111110",21556 => "01001010",21557 => "10000101",21558 => "11111000",21559 => "00101001",21560 => "11011101",21561 => "00110100",21562 => "11100001",21563 => "01110000",21564 => "01101111",21565 => "10111111",21566 => "10100000",21567 => "00101011",21568 => "01111101",21569 => "01110001",21570 => "11101111",21571 => "10100110",21572 => "01101111",21573 => "01001101",21574 => "11110100",21575 => "11000011",21576 => "11000100",21577 => "11100000",21578 => "01100011",21579 => "10001101",21580 => "10010001",21581 => "01001001",21582 => "10101101",21583 => "00101111",21584 => "01011100",21585 => "10111101",21586 => "00111000",21587 => "10010100",21588 => "00111101",21589 => "11011110",21590 => "01111110",21591 => "00101011",21592 => "10100011",21593 => "00000011",21594 => "11010001",21595 => "00100001",21596 => "01010000",21597 => "00001011",21598 => "00001000",21599 => "11100100",21600 => "01100110",21601 => "10000010",21602 => "11100101",21603 => "00101111",21604 => "10011100",21605 => "01011110",21606 => "10001101",21607 => "11001101",21608 => "10100101",21609 => "01011110",21610 => "11001010",21611 => "01101001",21612 => "00111011",21613 => "01100011",21614 => "10100011",21615 => "10011001",21616 => "01101110",21617 => "11001101",21618 => "01000011",21619 => "10111110",21620 => "01010100",21621 => "10010110",21622 => "11011100",21623 => "11011011",21624 => "11011111",21625 => "10101011",21626 => "01000000",21627 => "10010101",21628 => "01101111",21629 => "00110010",21630 => "00001010",21631 => "10001111",21632 => "01101011",21633 => "01100111",21634 => "00000110",21635 => "00101001",21636 => "01110111",21637 => "11010000",21638 => "01100101",21639 => "01010001",21640 => "01011010",21641 => "01011011",21642 => "00000111",21643 => "01100111",21644 => "01111010",21645 => "11001000",21646 => "10001101",21647 => "11111101",21648 => "11000111",21649 => "01101000",21650 => "00000101",21651 => "11010000",21652 => "10000110",21653 => "10010100",21654 => "00110000",21655 => "10110001",21656 => "01011001",21657 => "00101000",21658 => "11101111",21659 => "10111110",21660 => "01111000",21661 => "00000100",21662 => "10001111",21663 => "01011011",21664 => "11010111",21665 => "01010100",21666 => "10110000",21667 => "00010110",21668 => "01000001",21669 => "00101011",21670 => "10010000",21671 => "01111100",21672 => "11001001",21673 => "00111101",21674 => "01100110",21675 => "00010001",21676 => "10011001",21677 => "00101011",21678 => "00001010",21679 => "00100110",21680 => "00110101",21681 => "00010100",21682 => "00011100",21683 => "10010010",21684 => "11010110",21685 => "00001000",21686 => "00000101",21687 => "11010011",21688 => "11000001",21689 => "11010110",21690 => "11100111",21691 => "00100011",21692 => "01001000",21693 => "00111010",21694 => "10101010",21695 => "00010101",21696 => "00010000",21697 => "10001101",21698 => "00010010",21699 => "11001101",21700 => "00011101",21701 => "10010101",21702 => "11011011",21703 => "01110100",21704 => "01010111",21705 => "01000001",21706 => "01100000",21707 => "11001010",21708 => "11101010",21709 => "00000101",21710 => "11111110",21711 => "00111111",21712 => "00001011",21713 => "10011111",21714 => "00101100",21715 => "01011010",21716 => "00010100",21717 => "00010000",21718 => "11001001",21719 => "10011111",21720 => "11101101",21721 => "00101101",21722 => "10000010",21723 => "11010000",21724 => "00111011",21725 => "11011110",21726 => "11011110",21727 => "10000110",21728 => "01000010",21729 => "00011110",21730 => "10011111",21731 => "00000111",21732 => "01101101",21733 => "01110000",21734 => "10010100",21735 => "11111001",21736 => "01001000",21737 => "10111111",21738 => "11101111",21739 => "11111011",21740 => "11100010",21741 => "00010011",21742 => "01100101",21743 => "00111110",21744 => "01110110",21745 => "00110011",21746 => "01000010",21747 => "01010100",21748 => "10000001",21749 => "01110001",21750 => "01010111",21751 => "10100011",21752 => "11101010",21753 => "00101100",21754 => "00100001",21755 => "01101011",21756 => "00100001",21757 => "01000011",21758 => "01101001",21759 => "01110100",21760 => "00100111",21761 => "11101101",21762 => "00000001",21763 => "01011110",21764 => "10110110",21765 => "01111010",21766 => "10101011",21767 => "11010010",21768 => "00000101",21769 => "01110010",21770 => "01111011",21771 => "00111001",21772 => "01100100",21773 => "10111000",21774 => "11100011",21775 => "11010111",21776 => "10011100",21777 => "00001111",21778 => "00001000",21779 => "11010101",21780 => "01100100",21781 => "11000111",21782 => "01101110",21783 => "10011101",21784 => "01010010",21785 => "11111110",21786 => "11110111",21787 => "10001010",21788 => "00001100",21789 => "00101010",21790 => "10010010",21791 => "10011111",21792 => "00111110",21793 => "01001000",21794 => "01001010",21795 => "11111100",21796 => "10111001",21797 => "00010111",21798 => "00001000",21799 => "11001000",21800 => "10000110",21801 => "01111001",21802 => "01110010",21803 => "01100111",21804 => "11111101",21805 => "10010011",21806 => "10011011",21807 => "01100100",21808 => "11101111",21809 => "10000100",21810 => "01000100",21811 => "11110100",21812 => "01010011",21813 => "01101010",21814 => "01000010",21815 => "01010000",21816 => "00011000",21817 => "01101011",21818 => "00001111",21819 => "00010110",21820 => "00110011",21821 => "01001000",21822 => "11000000",21823 => "11010100",21824 => "00000110",21825 => "01111100",21826 => "11110110",21827 => "00011101",21828 => "10010010",21829 => "11011000",21830 => "10001100",21831 => "01000010",21832 => "00010110",21833 => "10110001",21834 => "01100111",21835 => "01010000",21836 => "11000011",21837 => "00101011",21838 => "10100000",21839 => "11101100",21840 => "00011000",21841 => "11010101",21842 => "11100011",21843 => "11001001",21844 => "00010111",21845 => "00011000",21846 => "00000011",21847 => "11011101",21848 => "11011101",21849 => "01101011",21850 => "01111001",21851 => "00100010",21852 => "11101000",21853 => "10000001",21854 => "01110010",21855 => "10100111",21856 => "11010010",21857 => "00011011",21858 => "00100100",21859 => "00110101",21860 => "01100000",21861 => "11101000",21862 => "01101101",21863 => "00110100",21864 => "00110111",21865 => "10100100",21866 => "10100100",21867 => "01001101",21868 => "01100101",21869 => "00110001",21870 => "11100110",21871 => "00000000",21872 => "00101100",21873 => "11110110",21874 => "11011011",21875 => "00111001",21876 => "00100010",21877 => "01011010",21878 => "00010110",21879 => "00101001",21880 => "01101000",21881 => "10000110",21882 => "11101000",21883 => "11110100",21884 => "11001000",21885 => "00111101",21886 => "11010011",21887 => "11100100",21888 => "10101100",21889 => "11001100",21890 => "00001110",21891 => "11001110",21892 => "01111010",21893 => "10011111",21894 => "01101111",21895 => "00011001",21896 => "10100010",21897 => "00010011",21898 => "00111000",21899 => "11110010",21900 => "10001110",21901 => "10100110",21902 => "00000010",21903 => "11011011",21904 => "00010111",21905 => "00001001",21906 => "10110111",21907 => "10001011",21908 => "11000110",21909 => "00111000",21910 => "10111111",21911 => "00101010",21912 => "00000110",21913 => "00010000",21914 => "10100001",21915 => "00011100",21916 => "00101010",21917 => "10001100",21918 => "10010001",21919 => "00100111",21920 => "10111010",21921 => "01101001",21922 => "10111010",21923 => "10101001",21924 => "01011011",21925 => "11100110",21926 => "11001110",21927 => "00000101",21928 => "00001110",21929 => "00010001",21930 => "11011101",21931 => "01111110",21932 => "10001001",21933 => "10111111",21934 => "10101110",21935 => "01001001",21936 => "10010111",21937 => "10110010",21938 => "00111111",21939 => "01010101",21940 => "11110100",21941 => "00101011",21942 => "10111100",21943 => "10011111",21944 => "10110100",21945 => "01110100",21946 => "01110010",21947 => "11111101",21948 => "00110111",21949 => "10111000",21950 => "00001101",21951 => "10111100",21952 => "00100000",21953 => "10100110",21954 => "11101010",21955 => "11100011",21956 => "10111011",21957 => "10110000",21958 => "11111000",21959 => "10011000",21960 => "10110010",21961 => "01100101",21962 => "11001010",21963 => "11100100",21964 => "10011100",21965 => "00110000",21966 => "11010100",21967 => "10100011",21968 => "11011010",21969 => "01100100",21970 => "01001011",21971 => "01000001",21972 => "01001001",21973 => "11010101",21974 => "01000111",21975 => "11101000",21976 => "00100001",21977 => "11011111",21978 => "11101000",21979 => "10001011",21980 => "11111110",21981 => "01010100",21982 => "10010100",21983 => "10111001",21984 => "11000110",21985 => "11100110",21986 => "10010011",21987 => "11000101",21988 => "00000101",21989 => "10101100",21990 => "00010011",21991 => "01000010",21992 => "01000101",21993 => "01010011",21994 => "10111111",21995 => "11011111",21996 => "10110011",21997 => "11000111",21998 => "01000111",21999 => "11101010",22000 => "11001111",22001 => "00101110",22002 => "00000000",22003 => "00010011",22004 => "01010111",22005 => "01101010",22006 => "01010010",22007 => "01100100",22008 => "01010111",22009 => "00010000",22010 => "10110111",22011 => "10011100",22012 => "00001100",22013 => "11011110",22014 => "00010011",22015 => "01010010",22016 => "10100011",22017 => "11110111",22018 => "00010011",22019 => "11001001",22020 => "01100000",22021 => "00001101",22022 => "10000101",22023 => "11010001",22024 => "11011011",22025 => "10100010",22026 => "00001110",22027 => "01100111",22028 => "11001111",22029 => "01101011",22030 => "00001001",22031 => "10111100",22032 => "00010110",22033 => "10101010",22034 => "10001101",22035 => "10001111",22036 => "00100010",22037 => "01101101",22038 => "00100001",22039 => "10001011",22040 => "10100011",22041 => "01010000",22042 => "11011100",22043 => "00000010",22044 => "11111111",22045 => "10111010",22046 => "11101100",22047 => "00000001",22048 => "11001010",22049 => "01001101",22050 => "11010100",22051 => "00110110",22052 => "11111110",22053 => "11100000",22054 => "01010001",22055 => "10010011",22056 => "01111101",22057 => "01111000",22058 => "01011101",22059 => "01001111",22060 => "00101110",22061 => "10101100",22062 => "11010000",22063 => "00001010",22064 => "01110000",22065 => "10100011",22066 => "10100010",22067 => "01010100",22068 => "11100101",22069 => "10011100",22070 => "00110000",22071 => "11001011",22072 => "01100110",22073 => "11110101",22074 => "01010110",22075 => "10101111",22076 => "10000010",22077 => "11001001",22078 => "10110011",22079 => "11111100",22080 => "11110110",22081 => "00001101",22082 => "10010110",22083 => "01111001",22084 => "10101101",22085 => "10111100",22086 => "01101000",22087 => "10010000",22088 => "10100111",22089 => "00000110",22090 => "01101101",22091 => "00100000",22092 => "00000010",22093 => "10010001",22094 => "11110100",22095 => "01110111",22096 => "10111101",22097 => "00111010",22098 => "00000101",22099 => "11010000",22100 => "01000011",22101 => "01101111",22102 => "00110101",22103 => "00110101",22104 => "11100011",22105 => "00111110",22106 => "00111000",22107 => "00000101",22108 => "01111010",22109 => "01010101",22110 => "10111010",22111 => "11000000",22112 => "11010011",22113 => "00110011",22114 => "10000100",22115 => "10010101",22116 => "10011110",22117 => "00010100",22118 => "11101101",22119 => "00101000",22120 => "00001110",22121 => "00010111",22122 => "11001110",22123 => "10101001",22124 => "10001101",22125 => "00000100",22126 => "00000100",22127 => "00010011",22128 => "01100111",22129 => "00101001",22130 => "01000011",22131 => "10111001",22132 => "01110010",22133 => "01100110",22134 => "11011111",22135 => "00110110",22136 => "10100110",22137 => "11111111",22138 => "00101101",22139 => "10001101",22140 => "00000001",22141 => "11110001",22142 => "10111110",22143 => "11100001",22144 => "10101010",22145 => "00110101",22146 => "01001010",22147 => "10010111",22148 => "01001101",22149 => "11011111",22150 => "01000100",22151 => "00111000",22152 => "10110100",22153 => "10010101",22154 => "00101001",22155 => "11011100",22156 => "11110101",22157 => "10111110",22158 => "10011111",22159 => "11101101",22160 => "11000110",22161 => "11011011",22162 => "01010010",22163 => "01000111",22164 => "01100101",22165 => "00000011",22166 => "00101000",22167 => "01101100",22168 => "01001010",22169 => "01111001",22170 => "00011101",22171 => "10111111",22172 => "01110110",22173 => "01011010",22174 => "00101001",22175 => "11001110",22176 => "10001011",22177 => "00011010",22178 => "00011011",22179 => "01111100",22180 => "00110110",22181 => "01001000",22182 => "10101011",22183 => "11011111",22184 => "11010010",22185 => "01000000",22186 => "00011100",22187 => "11100101",22188 => "11110100",22189 => "10001011",22190 => "00000110",22191 => "10110010",22192 => "01111110",22193 => "01101100",22194 => "11001110",22195 => "01111111",22196 => "00101001",22197 => "00010111",22198 => "00110111",22199 => "00011100",22200 => "10110100",22201 => "00110010",22202 => "00101011",22203 => "10010001",22204 => "11101011",22205 => "10101100",22206 => "10110011",22207 => "01100000",22208 => "01010011",22209 => "11111001",22210 => "11101110",22211 => "01100001",22212 => "00101001",22213 => "10110100",22214 => "10010011",22215 => "00001010",22216 => "11101011",22217 => "11110100",22218 => "10101110",22219 => "00110001",22220 => "00100010",22221 => "01100010",22222 => "00001001",22223 => "10001000",22224 => "01110110",22225 => "10011110",22226 => "11011100",22227 => "11000000",22228 => "11000110",22229 => "01100100",22230 => "10011010",22231 => "11000000",22232 => "01111011",22233 => "11001000",22234 => "10111010",22235 => "00110011",22236 => "11011110",22237 => "00101100",22238 => "01100001",22239 => "10000100",22240 => "00101011",22241 => "01101001",22242 => "11000010",22243 => "01011100",22244 => "01101011",22245 => "01010101",22246 => "01101110",22247 => "00011000",22248 => "11100101",22249 => "10011100",22250 => "00010011",22251 => "10010100",22252 => "00111010",22253 => "11001100",22254 => "10111101",22255 => "01101110",22256 => "11111111",22257 => "11110001",22258 => "10101001",22259 => "11000000",22260 => "10101000",22261 => "00011101",22262 => "11110111",22263 => "00100000",22264 => "01110010",22265 => "11010111",22266 => "01010010",22267 => "01000001",22268 => "01011010",22269 => "11001010",22270 => "01010111",22271 => "11000111",22272 => "11001011",22273 => "11011111",22274 => "10001111",22275 => "01110110",22276 => "01000101",22277 => "00101111",22278 => "10001100",22279 => "11110110",22280 => "10010111",22281 => "11111111",22282 => "10110010",22283 => "11010011",22284 => "11011100",22285 => "00110100",22286 => "11100111",22287 => "11110010",22288 => "00100000",22289 => "11011110",22290 => "11010011",22291 => "00000111",22292 => "11110100",22293 => "11101001",22294 => "11001111",22295 => "10111000",22296 => "10110111",22297 => "11000110",22298 => "10101010",22299 => "01011100",22300 => "00011001",22301 => "10101110",22302 => "01010011",22303 => "11011101",22304 => "01011100",22305 => "00100000",22306 => "10100101",22307 => "10110001",22308 => "11100110",22309 => "11111101",22310 => "11100110",22311 => "00101111",22312 => "00100001",22313 => "01000100",22314 => "00100000",22315 => "10101001",22316 => "01110010",22317 => "10000010",22318 => "10010110",22319 => "11100001",22320 => "11100100",22321 => "01000001",22322 => "00001101",22323 => "01101000",22324 => "10011110",22325 => "01011100",22326 => "10010000",22327 => "10010100",22328 => "11111101",22329 => "10010010",22330 => "11000100",22331 => "00000111",22332 => "10001111",22333 => "01111011",22334 => "10111100",22335 => "00111000",22336 => "11110100",22337 => "00010110",22338 => "11110110",22339 => "11011101",22340 => "10101000",22341 => "01110011",22342 => "11001011",22343 => "00100101",22344 => "01110101",22345 => "00101101",22346 => "01100011",22347 => "11001100",22348 => "10001001",22349 => "11001110",22350 => "00111100",22351 => "10110010",22352 => "10011101",22353 => "10110111",22354 => "01100111",22355 => "11000000",22356 => "01101000",22357 => "00010101",22358 => "01101001",22359 => "01100100",22360 => "11000100",22361 => "01111011",22362 => "00110010",22363 => "11011001",22364 => "00100111",22365 => "10000010",22366 => "01111111",22367 => "10100101",22368 => "00111010",22369 => "01101111",22370 => "00010011",22371 => "01000000",22372 => "11111111",22373 => "10011000",22374 => "00100000",22375 => "00000110",22376 => "10011011",22377 => "11110000",22378 => "10010101",22379 => "00000010",22380 => "10011100",22381 => "00111100",22382 => "10011010",22383 => "00101100",22384 => "01110011",22385 => "01111001",22386 => "10111010",22387 => "01000100",22388 => "01011111",22389 => "11111011",22390 => "11001011",22391 => "00011101",22392 => "01001000",22393 => "10000111",22394 => "01111111",22395 => "10001001",22396 => "11010000",22397 => "10010111",22398 => "11000011",22399 => "01111000",22400 => "01111010",22401 => "00101011",22402 => "00110001",22403 => "11010011",22404 => "11111111",22405 => "00100011",22406 => "01011101",22407 => "10100100",22408 => "00011000",22409 => "11001100",22410 => "01010111",22411 => "00100110",22412 => "11101100",22413 => "11111101",22414 => "01000100",22415 => "00111101",22416 => "01000111",22417 => "01011111",22418 => "00000000",22419 => "00011110",22420 => "11010111",22421 => "01110111",22422 => "10000100",22423 => "00011001",22424 => "00001100",22425 => "11010101",22426 => "10100010",22427 => "10110001",22428 => "01010000",22429 => "00001001",22430 => "00001010",22431 => "00011011",22432 => "10010111",22433 => "00101011",22434 => "10011011",22435 => "11010111",22436 => "11101100",22437 => "11110000",22438 => "10100001",22439 => "00111000",22440 => "10100101",22441 => "00001010",22442 => "11111011",22443 => "10100011",22444 => "11011001",22445 => "00100011",22446 => "10111100",22447 => "10100000",22448 => "00100111",22449 => "01110001",22450 => "11000110",22451 => "11111111",22452 => "11011001",22453 => "11100111",22454 => "11111110",22455 => "00100101",22456 => "00111111",22457 => "00101001",22458 => "10101101",22459 => "00010011",22460 => "10110110",22461 => "01010011",22462 => "10100110",22463 => "10110000",22464 => "00001011",22465 => "10101111",22466 => "00011010",22467 => "00011000",22468 => "00100101",22469 => "00100101",22470 => "11100000",22471 => "10101101",22472 => "00000001",22473 => "10110110",22474 => "01001101",22475 => "11001101",22476 => "00110011",22477 => "10001011",22478 => "01011000",22479 => "10111000",22480 => "10010001",22481 => "11101101",22482 => "01001100",22483 => "11100100",22484 => "11000011",22485 => "11101011",22486 => "00110110",22487 => "11010110",22488 => "00010110",22489 => "00111001",22490 => "11111101",22491 => "01000100",22492 => "10010101",22493 => "01111101",22494 => "10111100",22495 => "10010011",22496 => "10100101",22497 => "01001010",22498 => "00001111",22499 => "10110001",22500 => "00100000",22501 => "11111011",22502 => "00110110",22503 => "01000001",22504 => "10100100",22505 => "10000001",22506 => "10010111",22507 => "11100110",22508 => "10110001",22509 => "01111111",22510 => "10100100",22511 => "11111011",22512 => "10000111",22513 => "11101001",22514 => "00010010",22515 => "11001010",22516 => "01101111",22517 => "10110111",22518 => "10100111",22519 => "00101001",22520 => "00000100",22521 => "01001111",22522 => "00011000",22523 => "00010111",22524 => "11000001",22525 => "00110110",22526 => "10000010",22527 => "00101101",22528 => "11010100",22529 => "10001111",22530 => "01010100",22531 => "10010010",22532 => "10010010",22533 => "01111111",22534 => "00010111",22535 => "00010100",22536 => "01110011",22537 => "00101110",22538 => "01001000",22539 => "10011011",22540 => "01101111",22541 => "00001110",22542 => "00011100",22543 => "00010100",22544 => "10011000",22545 => "11100010",22546 => "00010001",22547 => "10011111",22548 => "00010011",22549 => "11110110",22550 => "11101101",22551 => "11101001",22552 => "10101011",22553 => "01011001",22554 => "00100111",22555 => "11011100",22556 => "11111100",22557 => "00000101",22558 => "01010010",22559 => "01100010",22560 => "01110101",22561 => "10010100",22562 => "00010111",22563 => "10010111",22564 => "01100101",22565 => "01000001",22566 => "01111100",22567 => "11100011",22568 => "10101010",22569 => "01010010",22570 => "11000110",22571 => "00101000",22572 => "11000010",22573 => "11010111",22574 => "00100000",22575 => "01001011",22576 => "01011000",22577 => "10111001",22578 => "10111111",22579 => "00111100",22580 => "11011001",22581 => "10010001",22582 => "10110001",22583 => "00111011",22584 => "10110011",22585 => "00100100",22586 => "10011100",22587 => "01000011",22588 => "10110001",22589 => "11110001",22590 => "10101100",22591 => "11000110",22592 => "00111010",22593 => "00011111",22594 => "11011100",22595 => "01000000",22596 => "11011001",22597 => "10110101",22598 => "01110110",22599 => "01100100",22600 => "11011100",22601 => "01000110",22602 => "11101000",22603 => "01100100",22604 => "11110001",22605 => "00101011",22606 => "00011111",22607 => "01000000",22608 => "00101110",22609 => "11110010",22610 => "01101011",22611 => "11000110",22612 => "11011001",22613 => "01000110",22614 => "01101011",22615 => "10011101",22616 => "11001001",22617 => "11111000",22618 => "11110111",22619 => "01100011",22620 => "01111010",22621 => "10011101",22622 => "10111111",22623 => "00000010",22624 => "00101110",22625 => "10111010",22626 => "10001111",22627 => "11111111",22628 => "11100111",22629 => "10110110",22630 => "10101011",22631 => "01111010",22632 => "10000110",22633 => "10010011",22634 => "00111110",22635 => "11101111",22636 => "10101100",22637 => "10110011",22638 => "10100101",22639 => "00101101",22640 => "01001111",22641 => "00110001",22642 => "10010111",22643 => "11001110",22644 => "11111100",22645 => "10101100",22646 => "10100010",22647 => "01000101",22648 => "01101101",22649 => "11000001",22650 => "11100101",22651 => "00101001",22652 => "00100110",22653 => "10110011",22654 => "11111011",22655 => "10111101",22656 => "00101000",22657 => "11110000",22658 => "00011111",22659 => "10011011",22660 => "01011010",22661 => "00100010",22662 => "01000000",22663 => "00101110",22664 => "00101010",22665 => "00100000",22666 => "01111100",22667 => "10010000",22668 => "10110101",22669 => "00111110",22670 => "10011111",22671 => "10100111",22672 => "10010101",22673 => "01001011",22674 => "11011100",22675 => "11000110",22676 => "11001010",22677 => "10100001",22678 => "00000010",22679 => "10110011",22680 => "11101011",22681 => "01010111",22682 => "00101101",22683 => "11101000",22684 => "01011011",22685 => "01110100",22686 => "10010100",22687 => "01110110",22688 => "11111001",22689 => "00000011",22690 => "10011110",22691 => "11100011",22692 => "11101101",22693 => "00110010",22694 => "00101111",22695 => "10011001",22696 => "10000100",22697 => "01100110",22698 => "11101100",22699 => "10110110",22700 => "11101110",22701 => "10010110",22702 => "11100011",22703 => "11110011",22704 => "11101100",22705 => "01110111",22706 => "10000001",22707 => "01101100",22708 => "00111101",22709 => "01111100",22710 => "00101110",22711 => "11100011",22712 => "11111001",22713 => "00011100",22714 => "10001010",22715 => "10111101",22716 => "10001100",22717 => "00010000",22718 => "11001001",22719 => "00101000",22720 => "00101101",22721 => "01100110",22722 => "00001100",22723 => "01000001",22724 => "01000111",22725 => "01001010",22726 => "00101110",22727 => "00010111",22728 => "00100001",22729 => "10010111",22730 => "01010000",22731 => "11110101",22732 => "10011111",22733 => "11100000",22734 => "00110111",22735 => "01001101",22736 => "11100111",22737 => "10011001",22738 => "00000011",22739 => "11000001",22740 => "00001011",22741 => "00100110",22742 => "00111001",22743 => "01011011",22744 => "01110101",22745 => "00110001",22746 => "10010101",22747 => "10010010",22748 => "11010000",22749 => "00101001",22750 => "10010110",22751 => "10001001",22752 => "10101110",22753 => "10100100",22754 => "11110110",22755 => "01011010",22756 => "00011110",22757 => "00001001",22758 => "10111011",22759 => "01011111",22760 => "10011001",22761 => "00011100",22762 => "10010110",22763 => "10110100",22764 => "11110000",22765 => "01011011",22766 => "11111010",22767 => "01000010",22768 => "10000011",22769 => "00000000",22770 => "11110110",22771 => "11000110",22772 => "00001111",22773 => "10010100",22774 => "01111110",22775 => "11100111",22776 => "11001000",22777 => "10010010",22778 => "01111111",22779 => "11011110",22780 => "00001100",22781 => "01100000",22782 => "11101010",22783 => "11001000",22784 => "10011001",22785 => "01110010",22786 => "11010101",22787 => "11010001",22788 => "00001010",22789 => "11101100",22790 => "11101110",22791 => "11110011",22792 => "11011111",22793 => "01001101",22794 => "00110110",22795 => "10101100",22796 => "11100110",22797 => "10110100",22798 => "10001100",22799 => "11001001",22800 => "00111001",22801 => "00010000",22802 => "00111101",22803 => "00000100",22804 => "01001110",22805 => "01010110",22806 => "01001110",22807 => "01100101",22808 => "00011101",22809 => "10110000",22810 => "00111011",22811 => "00010100",22812 => "00010000",22813 => "11100110",22814 => "10010000",22815 => "00001001",22816 => "10101010",22817 => "01111010",22818 => "00011101",22819 => "00111101",22820 => "11010110",22821 => "11011001",22822 => "11000001",22823 => "11000011",22824 => "11101110",22825 => "11110101",22826 => "10001101",22827 => "00011011",22828 => "01101101",22829 => "11010001",22830 => "00100011",22831 => "11111111",22832 => "01110110",22833 => "10000110",22834 => "11110100",22835 => "00000111",22836 => "10001111",22837 => "01101010",22838 => "01111011",22839 => "10010110",22840 => "10101100",22841 => "00000111",22842 => "11101000",22843 => "00000000",22844 => "10010111",22845 => "11100111",22846 => "00011011",22847 => "01100001",22848 => "01101001",22849 => "10100000",22850 => "00010010",22851 => "11000101",22852 => "00001010",22853 => "01111000",22854 => "01011110",22855 => "00110100",22856 => "11000000",22857 => "01110111",22858 => "01101111",22859 => "01110001",22860 => "10111100",22861 => "11111100",22862 => "01110001",22863 => "01010110",22864 => "11011101",22865 => "11101111",22866 => "00111000",22867 => "00010100",22868 => "10101011",22869 => "11110101",22870 => "01101110",22871 => "01100100",22872 => "11110110",22873 => "11111001",22874 => "01011101",22875 => "00010111",22876 => "10000001",22877 => "10011001",22878 => "01111111",22879 => "00110010",22880 => "10100101",22881 => "01110010",22882 => "00110110",22883 => "10000101",22884 => "10001110",22885 => "01100001",22886 => "00101111",22887 => "01100011",22888 => "10110110",22889 => "11001010",22890 => "10011001",22891 => "00101101",22892 => "00101010",22893 => "11011010",22894 => "00100011",22895 => "01101111",22896 => "11111010",22897 => "01010110",22898 => "11010000",22899 => "01111111",22900 => "01000101",22901 => "10001001",22902 => "10110000",22903 => "10001111",22904 => "10111010",22905 => "10011110",22906 => "01010011",22907 => "11100101",22908 => "01101111",22909 => "00101001",22910 => "01110010",22911 => "10000101",22912 => "10000111",22913 => "01110111",22914 => "01100110",22915 => "10101110",22916 => "11000100",22917 => "01100110",22918 => "01011010",22919 => "01100110",22920 => "10101001",22921 => "10000101",22922 => "11010001",22923 => "10011110",22924 => "10011100",22925 => "10011000",22926 => "10010000",22927 => "00101011",22928 => "10011001",22929 => "01110001",22930 => "11100101",22931 => "00100110",22932 => "01101011",22933 => "00001011",22934 => "00010001",22935 => "01110111",22936 => "01111011",22937 => "00001111",22938 => "00111100",22939 => "01111110",22940 => "10001000",22941 => "00111011",22942 => "01111101",22943 => "11110011",22944 => "01000001",22945 => "11000001",22946 => "10110000",22947 => "00101110",22948 => "00011100",22949 => "01100001",22950 => "00111011",22951 => "10010000",22952 => "00100010",22953 => "01010001",22954 => "10100110",22955 => "10100110",22956 => "10111100",22957 => "00001100",22958 => "01001100",22959 => "00011010",22960 => "10100001",22961 => "00000100",22962 => "01110111",22963 => "10010100",22964 => "00000001",22965 => "10111101",22966 => "10111000",22967 => "01100110",22968 => "10111001",22969 => "11110001",22970 => "11011011",22971 => "00100100",22972 => "00101011",22973 => "00110110",22974 => "01110011",22975 => "11001000",22976 => "01000100",22977 => "10100101",22978 => "10101011",22979 => "11101011",22980 => "00010010",22981 => "01111110",22982 => "00001101",22983 => "10111101",22984 => "00101011",22985 => "00111011",22986 => "10100111",22987 => "10010010",22988 => "00010110",22989 => "10110001",22990 => "11100010",22991 => "11101101",22992 => "01100010",22993 => "01000010",22994 => "00111101",22995 => "10110110",22996 => "11111110",22997 => "01001101",22998 => "11000010",22999 => "10110101",23000 => "00110101",23001 => "01010100",23002 => "10110001",23003 => "01011001",23004 => "11001111",23005 => "00111100",23006 => "01101111",23007 => "10101100",23008 => "00111000",23009 => "11101000",23010 => "01011010",23011 => "00010011",23012 => "10000011",23013 => "11110011",23014 => "10100101",23015 => "10100110",23016 => "01100110",23017 => "00001111",23018 => "01001010",23019 => "01100011",23020 => "00000010",23021 => "11100010",23022 => "10010001",23023 => "11000100",23024 => "11000010",23025 => "10100110",23026 => "10110011",23027 => "11110010",23028 => "00101000",23029 => "10001111",23030 => "01011001",23031 => "00001111",23032 => "00111111",23033 => "10000010",23034 => "11100101",23035 => "01001001",23036 => "01000100",23037 => "11111010",23038 => "11101111",23039 => "10110000",23040 => "10110011",23041 => "11001010",23042 => "10010100",23043 => "11111011",23044 => "10101110",23045 => "01110010",23046 => "01011011",23047 => "10110010",23048 => "01100000",23049 => "11110010",23050 => "01101111",23051 => "11101100",23052 => "00000101",23053 => "00010110",23054 => "01010110",23055 => "00000111",23056 => "00110010",23057 => "01100111",23058 => "01011111",23059 => "00100110",23060 => "00111001",23061 => "10011000",23062 => "10110100",23063 => "10001010",23064 => "11111101",23065 => "10011000",23066 => "10111110",23067 => "11011101",23068 => "11101010",23069 => "00001010",23070 => "11110001",23071 => "00101100",23072 => "11100011",23073 => "01111101",23074 => "11011111",23075 => "01100000",23076 => "01111110",23077 => "01111110",23078 => "11010111",23079 => "00000100",23080 => "11101001",23081 => "01101011",23082 => "11011110",23083 => "01110101",23084 => "01010100",23085 => "11010010",23086 => "01100010",23087 => "01111110",23088 => "01110001",23089 => "00001010",23090 => "10111101",23091 => "00100011",23092 => "11011000",23093 => "00101100",23094 => "00110001",23095 => "00000100",23096 => "10110111",23097 => "01011000",23098 => "01010101",23099 => "11011011",23100 => "01111100",23101 => "10110111",23102 => "11010011",23103 => "10111111",23104 => "01010111",23105 => "10011011",23106 => "01000110",23107 => "10110110",23108 => "11100000",23109 => "01101000",23110 => "01100100",23111 => "00010101",23112 => "01101011",23113 => "01100101",23114 => "11000101",23115 => "00001001",23116 => "10011000",23117 => "00000000",23118 => "00111010",23119 => "10100010",23120 => "10011111",23121 => "01000111",23122 => "10010000",23123 => "00101111",23124 => "11101010",23125 => "10100010",23126 => "00000110",23127 => "10010110",23128 => "11010000",23129 => "10010011",23130 => "00011000",23131 => "01111011",23132 => "00001011",23133 => "10011101",23134 => "01000010",23135 => "00001101",23136 => "11100010",23137 => "11000000",23138 => "11010010",23139 => "01111010",23140 => "11100000",23141 => "10110111",23142 => "01111110",23143 => "00001011",23144 => "11010001",23145 => "10110011",23146 => "11000001",23147 => "10101110",23148 => "10011111",23149 => "11001101",23150 => "01110111",23151 => "00010011",23152 => "00101001",23153 => "00011001",23154 => "01010100",23155 => "11110100",23156 => "01111000",23157 => "11011110",23158 => "00111110",23159 => "01100111",23160 => "00101001",23161 => "00111101",23162 => "10110010",23163 => "11111111",23164 => "01011111",23165 => "11011111",23166 => "01000011",23167 => "01111101",23168 => "10101101",23169 => "10111101",23170 => "01010110",23171 => "00011011",23172 => "01011100",23173 => "01101011",23174 => "11101100",23175 => "00111100",23176 => "00011100",23177 => "00101000",23178 => "01111001",23179 => "01001011",23180 => "10011100",23181 => "01010111",23182 => "10000110",23183 => "01010011",23184 => "01111001",23185 => "01100010",23186 => "10110110",23187 => "01101001",23188 => "00011000",23189 => "10001101",23190 => "00101001",23191 => "10001100",23192 => "10100011",23193 => "11011000",23194 => "01011011",23195 => "10101010",23196 => "01000111",23197 => "00100011",23198 => "10000010",23199 => "01010101",23200 => "10110111",23201 => "11101110",23202 => "10011011",23203 => "01100110",23204 => "01101110",23205 => "11000000",23206 => "00101011",23207 => "00110101",23208 => "10100001",23209 => "01000010",23210 => "11101001",23211 => "11110011",23212 => "10100000",23213 => "11001110",23214 => "01000111",23215 => "01100101",23216 => "11011101",23217 => "01001001",23218 => "11001110",23219 => "01011010",23220 => "00101011",23221 => "01011000",23222 => "01101010",23223 => "00101001",23224 => "10100000",23225 => "00101010",23226 => "10101011",23227 => "01101000",23228 => "11101010",23229 => "00001110",23230 => "11001000",23231 => "01100111",23232 => "01110010",23233 => "01000001",23234 => "01111111",23235 => "11011111",23236 => "11100101",23237 => "10001001",23238 => "00110110",23239 => "00111101",23240 => "10011000",23241 => "00110011",23242 => "01001101",23243 => "10010101",23244 => "00101100",23245 => "01110100",23246 => "01011100",23247 => "00111001",23248 => "00100101",23249 => "01110100",23250 => "00010100",23251 => "10001010",23252 => "00111111",23253 => "11011101",23254 => "01101010",23255 => "11100010",23256 => "00010111",23257 => "11011100",23258 => "11010111",23259 => "10010110",23260 => "01101001",23261 => "10111111",23262 => "11011101",23263 => "11011011",23264 => "11111000",23265 => "11100110",23266 => "11001001",23267 => "11010001",23268 => "11010011",23269 => "11111110",23270 => "11011010",23271 => "00110000",23272 => "11010011",23273 => "10000101",23274 => "00111010",23275 => "01100100",23276 => "10111000",23277 => "00101110",23278 => "00000001",23279 => "11101111",23280 => "11000011",23281 => "01011001",23282 => "01000101",23283 => "01101010",23284 => "10100010",23285 => "00100010",23286 => "00101101",23287 => "11100100",23288 => "00110101",23289 => "01111110",23290 => "10010110",23291 => "10001101",23292 => "01110011",23293 => "01101011",23294 => "01001101",23295 => "01111110",23296 => "01010101",23297 => "00101011",23298 => "01011011",23299 => "11000101",23300 => "10010011",23301 => "00001011",23302 => "01110111",23303 => "10110011",23304 => "11000110",23305 => "10001000",23306 => "11010001",23307 => "00000101",23308 => "11110111",23309 => "01100000",23310 => "01111010",23311 => "01001001",23312 => "10001010",23313 => "00110001",23314 => "10111101",23315 => "11110100",23316 => "10011100",23317 => "11010010",23318 => "10111011",23319 => "01011011",23320 => "11111111",23321 => "01101101",23322 => "00100110",23323 => "11000100",23324 => "01101000",23325 => "01101111",23326 => "00100000",23327 => "10011000",23328 => "10000111",23329 => "01110111",23330 => "00101000",23331 => "01110111",23332 => "11000101",23333 => "11001001",23334 => "10100100",23335 => "10111011",23336 => "00100101",23337 => "11110000",23338 => "00000011",23339 => "00111011",23340 => "10111010",23341 => "01000000",23342 => "00010000",23343 => "01011100",23344 => "11001001",23345 => "10110100",23346 => "10100011",23347 => "01101100",23348 => "01000011",23349 => "01111001",23350 => "10101100",23351 => "11001100",23352 => "00100000",23353 => "10110100",23354 => "11101100",23355 => "00111100",23356 => "11010010",23357 => "00000110",23358 => "01010011",23359 => "01101000",23360 => "00110010",23361 => "01001111",23362 => "11100100",23363 => "00001101",23364 => "01010101",23365 => "01101001",23366 => "10101001",23367 => "00111000",23368 => "10010110",23369 => "01111101",23370 => "11101101",23371 => "10011010",23372 => "01110111",23373 => "00100111",23374 => "10001001",23375 => "01100100",23376 => "10110000",23377 => "11001111",23378 => "01101110",23379 => "00100110",23380 => "00100101",23381 => "00000110",23382 => "00000011",23383 => "10101101",23384 => "10111010",23385 => "00001011",23386 => "10110000",23387 => "10000010",23388 => "10101010",23389 => "00000000",23390 => "10010011",23391 => "10001110",23392 => "10110111",23393 => "00010010",23394 => "10100001",23395 => "01110011",23396 => "00000010",23397 => "00011100",23398 => "00001000",23399 => "00101000",23400 => "00110110",23401 => "11110100",23402 => "10011110",23403 => "01110010",23404 => "00001100",23405 => "01011001",23406 => "10001110",23407 => "01101001",23408 => "10000100",23409 => "01111010",23410 => "00100110",23411 => "10001001",23412 => "01000001",23413 => "10110001",23414 => "10111111",23415 => "01110110",23416 => "10001011",23417 => "00011001",23418 => "00011101",23419 => "01010000",23420 => "11110011",23421 => "11011111",23422 => "11100001",23423 => "01101111",23424 => "10011000",23425 => "11100001",23426 => "10101000",23427 => "01101100",23428 => "10110100",23429 => "11000000",23430 => "00001000",23431 => "10110001",23432 => "00010001",23433 => "11010100",23434 => "11001011",23435 => "11111110",23436 => "10101111",23437 => "00001100",23438 => "01010111",23439 => "00100100",23440 => "01010110",23441 => "10100010",23442 => "11100000",23443 => "11001111",23444 => "00110000",23445 => "01101111",23446 => "11000000",23447 => "10100001",23448 => "10110000",23449 => "11000100",23450 => "01111101",23451 => "10101110",23452 => "00100101",23453 => "01101001",23454 => "01011111",23455 => "11000011",23456 => "01010010",23457 => "11101100",23458 => "00001101",23459 => "01001001",23460 => "11001111",23461 => "10101000",23462 => "00101110",23463 => "11101111",23464 => "10101011",23465 => "00100101",23466 => "11010001",23467 => "11110010",23468 => "11110001",23469 => "10000110",23470 => "01110000",23471 => "01101011",23472 => "10101000",23473 => "00110011",23474 => "11101101",23475 => "10011001",23476 => "01101111",23477 => "10000111",23478 => "01011110",23479 => "01100111",23480 => "10010011",23481 => "00011100",23482 => "11110010",23483 => "11010100",23484 => "11010111",23485 => "11100100",23486 => "01010100",23487 => "00000010",23488 => "01101011",23489 => "01100100",23490 => "01010101",23491 => "00101111",23492 => "01110000",23493 => "10111001",23494 => "00011010",23495 => "10011110",23496 => "01111101",23497 => "00110000",23498 => "00001001",23499 => "10110011",23500 => "11101110",23501 => "01011110",23502 => "00000010",23503 => "01010101",23504 => "01001110",23505 => "11111001",23506 => "01000010",23507 => "00011100",23508 => "00001011",23509 => "01100100",23510 => "00100010",23511 => "11101110",23512 => "01101110",23513 => "00010001",23514 => "11101100",23515 => "10101110",23516 => "01110110",23517 => "00100000",23518 => "00000011",23519 => "11110010",23520 => "10110111",23521 => "10110110",23522 => "00100010",23523 => "11100010",23524 => "01111111",23525 => "00000100",23526 => "10001010",23527 => "11000111",23528 => "10110101",23529 => "10110110",23530 => "11101000",23531 => "10000110",23532 => "11100101",23533 => "00110111",23534 => "00011101",23535 => "00000000",23536 => "00001100",23537 => "11100011",23538 => "00001001",23539 => "11100011",23540 => "11100011",23541 => "10010001",23542 => "10000110",23543 => "00110001",23544 => "00101101",23545 => "10111101",23546 => "00011011",23547 => "11100111",23548 => "00111100",23549 => "01000100",23550 => "10010110",23551 => "01000110",23552 => "11000101",23553 => "10111010",23554 => "11010001",23555 => "11011100",23556 => "11011001",23557 => "10100111",23558 => "10101111",23559 => "10101000",23560 => "01111011",23561 => "01010010",23562 => "01011010",23563 => "00101111",23564 => "01100110",23565 => "11000111",23566 => "01111110",23567 => "01010111",23568 => "00110100",23569 => "11111111",23570 => "01100110",23571 => "01100011",23572 => "10111110",23573 => "01011101",23574 => "11001001",23575 => "11000110",23576 => "10010111",23577 => "01111010",23578 => "11011101",23579 => "10101110",23580 => "00010111",23581 => "10110011",23582 => "11110101",23583 => "10111000",23584 => "00010100",23585 => "10101101",23586 => "10111011",23587 => "01010010",23588 => "00001001",23589 => "10100100",23590 => "00100100",23591 => "10000011",23592 => "11111000",23593 => "10110010",23594 => "10110111",23595 => "00010011",23596 => "10010011",23597 => "10010001",23598 => "10011101",23599 => "00100101",23600 => "00101011",23601 => "00001010",23602 => "01001110",23603 => "00001011",23604 => "00010011",23605 => "01000000",23606 => "11000010",23607 => "10100010",23608 => "01011011",23609 => "11101101",23610 => "10001110",23611 => "11100111",23612 => "11101010",23613 => "10111111",23614 => "10011001",23615 => "11101001",23616 => "10100000",23617 => "00001000",23618 => "10011011",23619 => "01001001",23620 => "10101000",23621 => "01000000",23622 => "00011000",23623 => "01110011",23624 => "01010110",23625 => "01000011",23626 => "01010011",23627 => "10101000",23628 => "01111111",23629 => "11100110",23630 => "01010011",23631 => "11100111",23632 => "00110110",23633 => "11111011",23634 => "01101010",23635 => "10011000",23636 => "01011111",23637 => "00010001",23638 => "01100111",23639 => "11011111",23640 => "11011010",23641 => "00101011",23642 => "00010010",23643 => "10101011",23644 => "11001001",23645 => "11011110",23646 => "01111110",23647 => "00101001",23648 => "11100100",23649 => "10010110",23650 => "01110001",23651 => "00100010",23652 => "01010010",23653 => "10010010",23654 => "01001000",23655 => "00100110",23656 => "00011111",23657 => "01000001",23658 => "01111000",23659 => "00101100",23660 => "10100011",23661 => "10011110",23662 => "01010110",23663 => "01001001",23664 => "01000000",23665 => "00010111",23666 => "01000110",23667 => "10011011",23668 => "11010101",23669 => "10101101",23670 => "11000010",23671 => "00110000",23672 => "10110110",23673 => "11111111",23674 => "00011001",23675 => "10011100",23676 => "00100101",23677 => "01011101",23678 => "01001100",23679 => "10101011",23680 => "01100010",23681 => "01111001",23682 => "00011101",23683 => "11001011",23684 => "00111000",23685 => "10101001",23686 => "11111100",23687 => "00000100",23688 => "01000111",23689 => "00110100",23690 => "00011010",23691 => "01010110",23692 => "01100001",23693 => "00110111",23694 => "11100111",23695 => "00010101",23696 => "01011000",23697 => "00101010",23698 => "01110101",23699 => "11010010",23700 => "10011011",23701 => "01111100",23702 => "11001000",23703 => "11100100",23704 => "01010111",23705 => "11011111",23706 => "10001000",23707 => "00010000",23708 => "11100000",23709 => "11011010",23710 => "11100111",23711 => "00010100",23712 => "10000000",23713 => "00110111",23714 => "00011011",23715 => "11111111",23716 => "01000100",23717 => "00001111",23718 => "01100110",23719 => "11110001",23720 => "10010011",23721 => "01100100",23722 => "11000110",23723 => "00001011",23724 => "00100110",23725 => "01001000",23726 => "10111010",23727 => "01110111",23728 => "01010110",23729 => "10001010",23730 => "11001010",23731 => "00011100",23732 => "11010110",23733 => "01000001",23734 => "10000101",23735 => "10001100",23736 => "01110011",23737 => "11101011",23738 => "11101111",23739 => "00101111",23740 => "10010010",23741 => "11000001",23742 => "10011011",23743 => "00011001",23744 => "10000000",23745 => "11000111",23746 => "00111110",23747 => "10010000",23748 => "10011001",23749 => "00111011",23750 => "11000100",23751 => "10101101",23752 => "11100101",23753 => "01100010",23754 => "00010010",23755 => "00000110",23756 => "01000011",23757 => "11001100",23758 => "01011001",23759 => "11100010",23760 => "00001111",23761 => "10101110",23762 => "11000001",23763 => "10111011",23764 => "11010111",23765 => "10101101",23766 => "01111011",23767 => "00101101",23768 => "00101011",23769 => "01111100",23770 => "10101000",23771 => "01010011",23772 => "00101011",23773 => "10100111",23774 => "10111101",23775 => "10100010",23776 => "00111000",23777 => "10001110",23778 => "01101000",23779 => "01110010",23780 => "00100010",23781 => "01110000",23782 => "11101010",23783 => "10110101",23784 => "00001000",23785 => "10100100",23786 => "11101110",23787 => "01100011",23788 => "01010010",23789 => "01010011",23790 => "11100010",23791 => "00000111",23792 => "10000101",23793 => "00110110",23794 => "01100111",23795 => "01010000",23796 => "01100011",23797 => "11001010",23798 => "00100000",23799 => "10101010",23800 => "00010011",23801 => "10001000",23802 => "00011110",23803 => "10100011",23804 => "11011111",23805 => "01000101",23806 => "11101100",23807 => "00111100",23808 => "11000000",23809 => "01110010",23810 => "10001000",23811 => "11011011",23812 => "01001000",23813 => "01001110",23814 => "01101000",23815 => "11011110",23816 => "10000110",23817 => "01110110",23818 => "01101010",23819 => "00100011",23820 => "11010001",23821 => "10000111",23822 => "00010101",23823 => "00100000",23824 => "11010110",23825 => "01111010",23826 => "00000010",23827 => "00001000",23828 => "10001010",23829 => "10101110",23830 => "10000101",23831 => "00110001",23832 => "01110111",23833 => "01100101",23834 => "10011110",23835 => "11111010",23836 => "11011111",23837 => "00011111",23838 => "00001111",23839 => "11110010",23840 => "10011101",23841 => "00110010",23842 => "01111110",23843 => "11000100",23844 => "01110101",23845 => "11011001",23846 => "00101000",23847 => "00111010",23848 => "01011001",23849 => "01110001",23850 => "10000100",23851 => "01110001",23852 => "11011000",23853 => "10000010",23854 => "10011100",23855 => "00100100",23856 => "10101100",23857 => "10000001",23858 => "00100101",23859 => "10011001",23860 => "01011101",23861 => "01010100",23862 => "01011001",23863 => "00011001",23864 => "00101101",23865 => "01100001",23866 => "01011001",23867 => "10001100",23868 => "00010000",23869 => "10101001",23870 => "11001111",23871 => "10010011",23872 => "00001010",23873 => "01110100",23874 => "11100001",23875 => "10001001",23876 => "11000001",23877 => "10100111",23878 => "00111010",23879 => "00101000",23880 => "00011011",23881 => "11000110",23882 => "11000110",23883 => "00001101",23884 => "00111010",23885 => "00111101",23886 => "11101100",23887 => "00100101",23888 => "10011110",23889 => "10001101",23890 => "10111011",23891 => "00000011",23892 => "10010111",23893 => "00011000",23894 => "00010000",23895 => "11100101",23896 => "10110011",23897 => "01100101",23898 => "11110010",23899 => "10100100",23900 => "10110010",23901 => "10001111",23902 => "01001111",23903 => "11001110",23904 => "00110001",23905 => "11110011",23906 => "00100000",23907 => "01000101",23908 => "01100010",23909 => "01011111",23910 => "11110101",23911 => "10101101",23912 => "10000000",23913 => "11001000",23914 => "00101010",23915 => "00111101",23916 => "01110001",23917 => "11101011",23918 => "01010010",23919 => "01010111",23920 => "01101001",23921 => "11100000",23922 => "10000111",23923 => "11001010",23924 => "11000101",23925 => "00110101",23926 => "10000111",23927 => "10000000",23928 => "11100001",23929 => "00000011",23930 => "00110101",23931 => "11110000",23932 => "01100101",23933 => "00110110",23934 => "01111011",23935 => "11010101",23936 => "10011101",23937 => "01000010",23938 => "11011111",23939 => "11011011",23940 => "00111101",23941 => "00001010",23942 => "10010110",23943 => "01001001",23944 => "11010000",23945 => "11011110",23946 => "11100100",23947 => "01101110",23948 => "10010000",23949 => "11010000",23950 => "01101111",23951 => "01101111",23952 => "11110000",23953 => "00101000",23954 => "10111111",23955 => "10000110",23956 => "11000110",23957 => "01000001",23958 => "11011011",23959 => "00100000",23960 => "11010010",23961 => "00110011",23962 => "11101001",23963 => "01011010",23964 => "11010010",23965 => "11100010",23966 => "01000001",23967 => "00000100",23968 => "01100011",23969 => "10111001",23970 => "11110011",23971 => "11110011",23972 => "01111101",23973 => "11100100",23974 => "01101011",23975 => "01010100",23976 => "01000110",23977 => "00110100",23978 => "01011011",23979 => "11011001",23980 => "10100110",23981 => "01011100",23982 => "11010010",23983 => "11000000",23984 => "11001001",23985 => "01000001",23986 => "10100010",23987 => "11111110",23988 => "00000000",23989 => "00111100",23990 => "01100000",23991 => "10001000",23992 => "01000111",23993 => "00010111",23994 => "11000001",23995 => "01111111",23996 => "10111001",23997 => "11100010",23998 => "10100111",23999 => "01011010",24000 => "10100111",24001 => "00100011",24002 => "10001100",24003 => "10110110",24004 => "00100000",24005 => "01001100",24006 => "01011010",24007 => "10111110",24008 => "01010001",24009 => "11011110",24010 => "01100100",24011 => "01001011",24012 => "00110101",24013 => "10000100",24014 => "00001110",24015 => "11010111",24016 => "01100011",24017 => "00010010",24018 => "11000000",24019 => "10010101",24020 => "01011101",24021 => "10001110",24022 => "11010011",24023 => "01101000",24024 => "00100010",24025 => "00001111",24026 => "10000010",24027 => "10010110",24028 => "00100001",24029 => "01010100",24030 => "11000111",24031 => "10001100",24032 => "00110110",24033 => "11101101",24034 => "11010010",24035 => "10000000",24036 => "01110110",24037 => "10000011",24038 => "01111011",24039 => "01110010",24040 => "11001111",24041 => "11101101",24042 => "00011101",24043 => "10010100",24044 => "01111000",24045 => "00000110",24046 => "00100101",24047 => "01001101",24048 => "10000101",24049 => "00001000",24050 => "00110011",24051 => "01100110",24052 => "11111011",24053 => "00101001",24054 => "11010100",24055 => "01010111",24056 => "00010001",24057 => "10001010",24058 => "00110011",24059 => "11111000",24060 => "00111010",24061 => "11001110",24062 => "11101110",24063 => "00110111",24064 => "11110000",24065 => "00100011",24066 => "10010101",24067 => "00101011",24068 => "11110101",24069 => "10100010",24070 => "01000010",24071 => "00111111",24072 => "11000011",24073 => "01000010",24074 => "00000101",24075 => "10001001",24076 => "01011010",24077 => "11001000",24078 => "00101001",24079 => "11000110",24080 => "11010111",24081 => "00111011",24082 => "10011101",24083 => "00001000",24084 => "00111111",24085 => "00111101",24086 => "00110011",24087 => "11100111",24088 => "00100010",24089 => "11000101",24090 => "10101011",24091 => "00111000",24092 => "01111010",24093 => "01111111",24094 => "01110111",24095 => "10001110",24096 => "10111011",24097 => "10101101",24098 => "11000010",24099 => "11010110",24100 => "11010111",24101 => "11100100",24102 => "00111100",24103 => "11011001",24104 => "10100010",24105 => "01100100",24106 => "01101000",24107 => "11000001",24108 => "10110110",24109 => "11100000",24110 => "10001101",24111 => "01110001",24112 => "00010101",24113 => "10000111",24114 => "11110010",24115 => "10011100",24116 => "10000010",24117 => "00001000",24118 => "01001011",24119 => "10011010",24120 => "10101000",24121 => "00110011",24122 => "11000111",24123 => "10010000",24124 => "11011000",24125 => "11011110",24126 => "11000010",24127 => "11001111",24128 => "10010101",24129 => "10011101",24130 => "00101100",24131 => "00001000",24132 => "10001011",24133 => "01000010",24134 => "00010000",24135 => "11010000",24136 => "10101000",24137 => "01101101",24138 => "00101111",24139 => "10010100",24140 => "00011010",24141 => "10110110",24142 => "00111011",24143 => "11001101",24144 => "10000111",24145 => "00110001",24146 => "01011001",24147 => "10101101",24148 => "11100111",24149 => "10011001",24150 => "00000110",24151 => "11000101",24152 => "00010111",24153 => "10011000",24154 => "01001000",24155 => "00111010",24156 => "00001000",24157 => "10010011",24158 => "10110010",24159 => "10010101",24160 => "10001100",24161 => "00101010",24162 => "10001000",24163 => "11001010",24164 => "11110010",24165 => "00101100",24166 => "11010111",24167 => "00000100",24168 => "10110111",24169 => "01011110",24170 => "11100000",24171 => "00110110",24172 => "11001100",24173 => "11011111",24174 => "01101001",24175 => "11100011",24176 => "00010001",24177 => "00001100",24178 => "11100010",24179 => "01011110",24180 => "11010001",24181 => "01110001",24182 => "01100011",24183 => "11001101",24184 => "01100101",24185 => "10110001",24186 => "11101110",24187 => "01010010",24188 => "00010001",24189 => "11101011",24190 => "10110101",24191 => "01000011",24192 => "10010000",24193 => "01011011",24194 => "10111101",24195 => "00011011",24196 => "10000100",24197 => "01011000",24198 => "00110110",24199 => "00001111",24200 => "00100000",24201 => "00010011",24202 => "10000111",24203 => "10100000",24204 => "00011001",24205 => "11111000",24206 => "10111100",24207 => "10100010",24208 => "00000101",24209 => "11110010",24210 => "10101010",24211 => "10111000",24212 => "11001001",24213 => "01101001",24214 => "10010011",24215 => "11011101",24216 => "00011010",24217 => "11101010",24218 => "00010111",24219 => "10111101",24220 => "10110010",24221 => "10010011",24222 => "11010111",24223 => "11101000",24224 => "01001111",24225 => "11101110",24226 => "00001100",24227 => "10101101",24228 => "01000010",24229 => "00101001",24230 => "10001110",24231 => "11110000",24232 => "11011100",24233 => "00000001",24234 => "10001111",24235 => "01100011",24236 => "11010001",24237 => "10100111",24238 => "00111111",24239 => "00111101",24240 => "01001110",24241 => "00010001",24242 => "10100001",24243 => "01100101",24244 => "10010001",24245 => "00011100",24246 => "10111111",24247 => "00001010",24248 => "01100100",24249 => "10101010",24250 => "11001110",24251 => "11011101",24252 => "00011010",24253 => "10110011",24254 => "00110111",24255 => "00100011",24256 => "00001101",24257 => "00101110",24258 => "11010110",24259 => "11101101",24260 => "10100111",24261 => "01000000",24262 => "01100011",24263 => "10000110",24264 => "10000100",24265 => "00100000",24266 => "11110010",24267 => "00100100",24268 => "00101111",24269 => "11011010",24270 => "10111101",24271 => "01001110",24272 => "00000010",24273 => "00110110",24274 => "00111110",24275 => "01100011",24276 => "01011010",24277 => "11011111",24278 => "10010000",24279 => "00110011",24280 => "01001111",24281 => "11000110",24282 => "00000101",24283 => "00111000",24284 => "01110101",24285 => "11010111",24286 => "10001110",24287 => "01011001",24288 => "00101000",24289 => "00100000",24290 => "00010110",24291 => "11100011",24292 => "00011000",24293 => "01000101",24294 => "01100011",24295 => "10111111",24296 => "11000110",24297 => "11110100",24298 => "00100010",24299 => "11110110",24300 => "00101010",24301 => "10010011",24302 => "00101010",24303 => "01001110",24304 => "00110001",24305 => "10100100",24306 => "01101000",24307 => "00010010",24308 => "01101001",24309 => "00101010",24310 => "11011001",24311 => "11111110",24312 => "01000000",24313 => "01001111",24314 => "01011111",24315 => "01011111",24316 => "00000111",24317 => "01010010",24318 => "01101101",24319 => "11000101",24320 => "01011100",24321 => "01100101",24322 => "10001011",24323 => "11000011",24324 => "11000110",24325 => "11001010",24326 => "01110110",24327 => "01011000",24328 => "11001001",24329 => "11101000",24330 => "01101101",24331 => "01100110",24332 => "01100100",24333 => "00100000",24334 => "00111011",24335 => "10001011",24336 => "01111000",24337 => "10000110",24338 => "10010010",24339 => "11010000",24340 => "00011010",24341 => "10100111",24342 => "00111110",24343 => "01101110",24344 => "01110011",24345 => "01001110",24346 => "11100001",24347 => "11011101",24348 => "00111110",24349 => "10001010",24350 => "00000100",24351 => "10101010",24352 => "00000111",24353 => "01011111",24354 => "10001111",24355 => "00110011",24356 => "10110100",24357 => "00111110",24358 => "10111111",24359 => "00111111",24360 => "10111011",24361 => "10001000",24362 => "11000011",24363 => "01001101",24364 => "10100000",24365 => "01010000",24366 => "01100101",24367 => "00011101",24368 => "01001011",24369 => "10101111",24370 => "11111101",24371 => "01001101",24372 => "10111010",24373 => "00011110",24374 => "11111001",24375 => "00101110",24376 => "01011100",24377 => "00101110",24378 => "10101010",24379 => "10110101",24380 => "01011010",24381 => "11111111",24382 => "10111100",24383 => "01000001",24384 => "10001111",24385 => "01000000",24386 => "10001111",24387 => "01101011",24388 => "00111011",24389 => "11100110",24390 => "10100000",24391 => "00011001",24392 => "00011011",24393 => "10000110",24394 => "11100011",24395 => "00100100",24396 => "00110100",24397 => "00011100",24398 => "11101111",24399 => "11011011",24400 => "01101010",24401 => "10001010",24402 => "11101000",24403 => "01111110",24404 => "10100011",24405 => "01100000",24406 => "10110100",24407 => "00010110",24408 => "10110001",24409 => "00110110",24410 => "11110010",24411 => "11001111",24412 => "10111001",24413 => "01110110",24414 => "00000110",24415 => "00100101",24416 => "10000000",24417 => "01011001",24418 => "10100100",24419 => "10010100",24420 => "10000101",24421 => "01010001",24422 => "11110001",24423 => "10111100",24424 => "01001000",24425 => "11010111",24426 => "00000110",24427 => "11101100",24428 => "01000110",24429 => "10100100",24430 => "01010101",24431 => "01101111",24432 => "00111010",24433 => "01110110",24434 => "11101011",24435 => "10000101",24436 => "11111101",24437 => "01101011",24438 => "10001111",24439 => "11011100",24440 => "00110101",24441 => "10010100",24442 => "01001010",24443 => "11111001",24444 => "11101000",24445 => "11010010",24446 => "10001111",24447 => "11001110",24448 => "00100110",24449 => "00010101",24450 => "10111110",24451 => "11110111",24452 => "00111001",24453 => "00001011",24454 => "10110110",24455 => "10010010",24456 => "01101001",24457 => "10011011",24458 => "11000110",24459 => "10110011",24460 => "00010101",24461 => "00101100",24462 => "00111011",24463 => "01010010",24464 => "10011111",24465 => "11010000",24466 => "10111100",24467 => "10101011",24468 => "11100100",24469 => "10110011",24470 => "01000000",24471 => "00010000",24472 => "01111100",24473 => "01000001",24474 => "00000110",24475 => "10001000",24476 => "01101101",24477 => "00110101",24478 => "00100010",24479 => "00001110",24480 => "01001011",24481 => "00011000",24482 => "10000010",24483 => "00100011",24484 => "11100111",24485 => "11100000",24486 => "00101111",24487 => "00000101",24488 => "01000010",24489 => "10001101",24490 => "01111011",24491 => "11001100",24492 => "00010101",24493 => "10000010",24494 => "00111010",24495 => "00100101",24496 => "11101101",24497 => "01111000",24498 => "00010011",24499 => "11001010",24500 => "11100001",24501 => "11111111",24502 => "11111110",24503 => "11001000",24504 => "11001000",24505 => "01010110",24506 => "01110000",24507 => "10011000",24508 => "00011111",24509 => "11011000",24510 => "11110100",24511 => "00110101",24512 => "10011001",24513 => "01100010",24514 => "11001101",24515 => "00111011",24516 => "11100100",24517 => "10101100",24518 => "10000100",24519 => "01011010",24520 => "00011001",24521 => "00000111",24522 => "11001010",24523 => "01000010",24524 => "00010100",24525 => "01110000",24526 => "01011110",24527 => "01110110",24528 => "10000111",24529 => "01011111",24530 => "01110110",24531 => "00101000",24532 => "01110000",24533 => "10111110",24534 => "00100111",24535 => "00001001",24536 => "10110010",24537 => "00100011",24538 => "00011000",24539 => "01110010",24540 => "10010001",24541 => "10111010",24542 => "00110100",24543 => "00111111",24544 => "01011001",24545 => "01111011",24546 => "10111011",24547 => "01111011",24548 => "00101011",24549 => "01010001",24550 => "00010010",24551 => "10100001",24552 => "00010111",24553 => "10100111",24554 => "11010111",24555 => "00011101",24556 => "00111110",24557 => "00011110",24558 => "11100011",24559 => "10110101",24560 => "10000101",24561 => "10110111",24562 => "10111001",24563 => "11010100",24564 => "11101010",24565 => "00111010",24566 => "01101011",24567 => "11001001",24568 => "01100011",24569 => "11001011",24570 => "01011110",24571 => "11010011",24572 => "00000011",24573 => "10101000",24574 => "10011001",24575 => "11010010",24576 => "11001111",24577 => "11101100",24578 => "01100001",24579 => "00010111",24580 => "11110011",24581 => "10000010",24582 => "11101001",24583 => "11001011",24584 => "00011101",24585 => "01111011",24586 => "01111011",24587 => "10001101",24588 => "01101100",24589 => "01111111",24590 => "10011001",24591 => "00010001",24592 => "11101011",24593 => "11111000",24594 => "10001110",24595 => "01101101",24596 => "11011110",24597 => "00010000",24598 => "00101000",24599 => "00100110",24600 => "00111001",24601 => "11111000",24602 => "10001011",24603 => "11110110",24604 => "01001110",24605 => "11000110",24606 => "11110100",24607 => "10111011",24608 => "10010010",24609 => "10100000",24610 => "01000110",24611 => "10100010",24612 => "01101101",24613 => "10111001",24614 => "00100010",24615 => "11011110",24616 => "00010110",24617 => "01001010",24618 => "10010101",24619 => "01010111",24620 => "00110111",24621 => "01110111",24622 => "01100001",24623 => "10101001",24624 => "11111000",24625 => "00101100",24626 => "01111111",24627 => "01110010",24628 => "11011010",24629 => "00101000",24630 => "00100110",24631 => "01000100",24632 => "11111100",24633 => "10000010",24634 => "00100111",24635 => "11110011",24636 => "11000001",24637 => "00101101",24638 => "00011111",24639 => "00001011",24640 => "10011011",24641 => "11010101",24642 => "11110111",24643 => "01110101",24644 => "01100110",24645 => "11111110",24646 => "10111101",24647 => "11111111",24648 => "00011101",24649 => "00111101",24650 => "10101101",24651 => "10110010",24652 => "11111100",24653 => "01010001",24654 => "11101110",24655 => "00101011",24656 => "01001010",24657 => "11011101",24658 => "10000000",24659 => "11101111",24660 => "11111110",24661 => "10101000",24662 => "11111001",24663 => "01011001",24664 => "10100101",24665 => "01000010",24666 => "10110001",24667 => "10100011",24668 => "10001100",24669 => "10001110",24670 => "11011111",24671 => "01111000",24672 => "10110111",24673 => "11111110",24674 => "10100001",24675 => "01111011",24676 => "10010100",24677 => "11111001",24678 => "01001011",24679 => "01101110",24680 => "10101110",24681 => "00010101",24682 => "11110011",24683 => "11110111",24684 => "10000100",24685 => "01010100",24686 => "01110001",24687 => "00100001",24688 => "00011010",24689 => "00000010",24690 => "11111011",24691 => "10110011",24692 => "01100101",24693 => "00100100",24694 => "11001010",24695 => "00101010",24696 => "00010001",24697 => "00001000",24698 => "01111101",24699 => "11110010",24700 => "01100010",24701 => "10011101",24702 => "10101010",24703 => "01001010",24704 => "00010111",24705 => "10110101",24706 => "00001100",24707 => "00010000",24708 => "01001100",24709 => "01001011",24710 => "01011110",24711 => "10101001",24712 => "11110000",24713 => "10111001",24714 => "00111001",24715 => "00101000",24716 => "01010000",24717 => "11010111",24718 => "11100111",24719 => "11100011",24720 => "11101101",24721 => "00010100",24722 => "10100101",24723 => "11010001",24724 => "00100111",24725 => "01101001",24726 => "00011101",24727 => "00100000",24728 => "11011011",24729 => "00010000",24730 => "00001111",24731 => "10101111",24732 => "00101101",24733 => "00110010",24734 => "10001000",24735 => "10101100",24736 => "11100111",24737 => "01000111",24738 => "10011110",24739 => "10101111",24740 => "10101110",24741 => "10101010",24742 => "00011001",24743 => "11100111",24744 => "10011010",24745 => "10011001",24746 => "10111000",24747 => "11000001",24748 => "01011001",24749 => "10100110",24750 => "10000010",24751 => "00101101",24752 => "01001000",24753 => "00100101",24754 => "10011101",24755 => "11001111",24756 => "11111101",24757 => "00000011",24758 => "01111001",24759 => "00001010",24760 => "01110001",24761 => "11001101",24762 => "01110000",24763 => "11011010",24764 => "10100111",24765 => "11000101",24766 => "01001000",24767 => "01100111",24768 => "11010111",24769 => "00000101",24770 => "11101001",24771 => "11100010",24772 => "10111111",24773 => "01101100",24774 => "00100000",24775 => "11000101",24776 => "10101110",24777 => "01010100",24778 => "00100001",24779 => "00001100",24780 => "10010000",24781 => "00011110",24782 => "10001101",24783 => "01011010",24784 => "11100010",24785 => "01010100",24786 => "00101000",24787 => "11110000",24788 => "01010011",24789 => "11100000",24790 => "00101000",24791 => "00100000",24792 => "11001010",24793 => "01000110",24794 => "00011111",24795 => "01100111",24796 => "11111001",24797 => "01000111",24798 => "01001010",24799 => "01001110",24800 => "10100000",24801 => "11000010",24802 => "00000111",24803 => "11111111",24804 => "11010100",24805 => "00000001",24806 => "10101110",24807 => "10110010",24808 => "10100100",24809 => "11011011",24810 => "01111010",24811 => "10001111",24812 => "00010010",24813 => "01010000",24814 => "01110111",24815 => "01000001",24816 => "00111001",24817 => "11011011",24818 => "00110001",24819 => "11111100",24820 => "11100100",24821 => "01011111",24822 => "01100010",24823 => "01000000",24824 => "01110001",24825 => "10111110",24826 => "11111101",24827 => "00000111",24828 => "11001011",24829 => "11100100",24830 => "11001011",24831 => "10011010",24832 => "00110100",24833 => "10001111",24834 => "01100101",24835 => "01010001",24836 => "10110000",24837 => "11000001",24838 => "10010101",24839 => "10111111",24840 => "11001111",24841 => "00011000",24842 => "01110011",24843 => "10010101",24844 => "01000001",24845 => "10001000",24846 => "10101001",24847 => "00001111",24848 => "11000011",24849 => "00110000",24850 => "00101101",24851 => "10010010",24852 => "10110001",24853 => "10101001",24854 => "10001000",24855 => "11110110",24856 => "10010101",24857 => "00111100",24858 => "01101011",24859 => "01011000",24860 => "00101010",24861 => "01001001",24862 => "11010100",24863 => "10100100",24864 => "01100000",24865 => "11110111",24866 => "11001000",24867 => "10111110",24868 => "11000101",24869 => "11011101",24870 => "11001000",24871 => "00000000",24872 => "10110111",24873 => "00001110",24874 => "01110000",24875 => "11100110",24876 => "11100011",24877 => "10111001",24878 => "11111101",24879 => "00110010",24880 => "10101000",24881 => "00010011",24882 => "00110111",24883 => "11000110",24884 => "11010111",24885 => "10001011",24886 => "11101001",24887 => "01010001",24888 => "11010100",24889 => "10100110",24890 => "11110011",24891 => "01001101",24892 => "11001010",24893 => "00110000",24894 => "01000110",24895 => "01011100",24896 => "10010000",24897 => "10000101",24898 => "11011110",24899 => "01001010",24900 => "10011110",24901 => "00001101",24902 => "10111000",24903 => "00011111",24904 => "01100000",24905 => "01111101",24906 => "01001100",24907 => "00000001",24908 => "10001001",24909 => "01011100",24910 => "11010101",24911 => "10111001",24912 => "00101111",24913 => "00000100",24914 => "10111110",24915 => "00111100",24916 => "00000000",24917 => "10001100",24918 => "10110001",24919 => "10001110",24920 => "01010101",24921 => "10110010",24922 => "11110110",24923 => "01100001",24924 => "11100000",24925 => "01111010",24926 => "10000101",24927 => "01011110",24928 => "00110111",24929 => "00110011",24930 => "01000101",24931 => "11011110",24932 => "00100101",24933 => "01101011",24934 => "11000100",24935 => "10110011",24936 => "00001100",24937 => "10111100",24938 => "01011000",24939 => "11011111",24940 => "11000111",24941 => "10011110",24942 => "01000101",24943 => "00010100",24944 => "00110011",24945 => "00001111",24946 => "01110110",24947 => "10011010",24948 => "01010101",24949 => "11111001",24950 => "11101111",24951 => "10010111",24952 => "11110011",24953 => "01000111",24954 => "01111011",24955 => "11001010",24956 => "01100111",24957 => "10101101",24958 => "10111011",24959 => "01111101",24960 => "10011010",24961 => "10001101",24962 => "10000110",24963 => "10000101",24964 => "10110011",24965 => "00110111",24966 => "10011100",24967 => "00010001",24968 => "10000110",24969 => "10101111",24970 => "00010000",24971 => "00101101",24972 => "01011011",24973 => "01110000",24974 => "11001111",24975 => "10001101",24976 => "11000010",24977 => "01010011",24978 => "01101111",24979 => "01000111",24980 => "01111001",24981 => "00111010",24982 => "11100101",24983 => "00100011",24984 => "10001100",24985 => "01011100",24986 => "01110001",24987 => "01000010",24988 => "11010110",24989 => "00011011",24990 => "00001101",24991 => "00110011",24992 => "10110100",24993 => "00100111",24994 => "11111001",24995 => "00111011",24996 => "00100101",24997 => "01011110",24998 => "01010101",24999 => "11001010",25000 => "11010000",25001 => "00101000",25002 => "10011011",25003 => "00101101",25004 => "11110100",25005 => "00011001",25006 => "11010100",25007 => "01011110",25008 => "11100000",25009 => "00000100",25010 => "10110111",25011 => "10111001",25012 => "10111001",25013 => "01000011",25014 => "10001011",25015 => "11011111",25016 => "00011011",25017 => "01100111",25018 => "10111001",25019 => "01000111",25020 => "01000111",25021 => "00000000",25022 => "01010111",25023 => "10011100",25024 => "00000100",25025 => "11111110",25026 => "11100101",25027 => "00011000",25028 => "00110100",25029 => "11101000",25030 => "11110010",25031 => "01010111",25032 => "11111110",25033 => "00101111",25034 => "10001110",25035 => "01001001",25036 => "11001101",25037 => "00100101",25038 => "00000100",25039 => "01000010",25040 => "01101101",25041 => "00110100",25042 => "10111001",25043 => "11011001",25044 => "01011101",25045 => "11111100",25046 => "01111010",25047 => "11000011",25048 => "10001011",25049 => "10000001",25050 => "10001011",25051 => "11010110",25052 => "11011110",25053 => "01100000",25054 => "10011111",25055 => "00110100",25056 => "00100011",25057 => "11110010",25058 => "10110101",25059 => "11101110",25060 => "10110101",25061 => "10011000",25062 => "11011111",25063 => "01000110",25064 => "10111111",25065 => "01000000",25066 => "01101010",25067 => "01111110",25068 => "01000001",25069 => "00000000",25070 => "00011111",25071 => "10111111",25072 => "01111111",25073 => "10110000",25074 => "11101111",25075 => "11001111",25076 => "11101100",25077 => "10011010",25078 => "11110001",25079 => "01000011",25080 => "01000010",25081 => "00000101",25082 => "10010111",25083 => "11110100",25084 => "00010101",25085 => "01101010",25086 => "01000110",25087 => "10101111",25088 => "11100001",25089 => "00011110",25090 => "11000010",25091 => "10011101",25092 => "11011000",25093 => "11101001",25094 => "11100101",25095 => "10011000",25096 => "10110010",25097 => "01110101",25098 => "01110011",25099 => "00101111",25100 => "11110011",25101 => "11000111",25102 => "00100110",25103 => "10010001",25104 => "11111100",25105 => "10010010",25106 => "01000010",25107 => "11001111",25108 => "01001110",25109 => "10101111",25110 => "00100100",25111 => "10010010",25112 => "01001010",25113 => "01001000",25114 => "01011111",25115 => "00111001",25116 => "00111011",25117 => "01011011",25118 => "11001100",25119 => "00010011",25120 => "01000110",25121 => "11101101",25122 => "10101111",25123 => "11010110",25124 => "01011110",25125 => "00110101",25126 => "11011110",25127 => "00001010",25128 => "00011011",25129 => "00011110",25130 => "10000011",25131 => "00001101",25132 => "10110101",25133 => "11010100",25134 => "10101100",25135 => "01010101",25136 => "10111111",25137 => "10001100",25138 => "01110001",25139 => "01110001",25140 => "00100001",25141 => "01000010",25142 => "00000110",25143 => "00000110",25144 => "11101011",25145 => "01001101",25146 => "10110011",25147 => "11000001",25148 => "10001111",25149 => "11110110",25150 => "01110010",25151 => "11001000",25152 => "10000011",25153 => "00100001",25154 => "01011000",25155 => "01101111",25156 => "10100011",25157 => "10101011",25158 => "10110111",25159 => "01111100",25160 => "11110111",25161 => "00110001",25162 => "11100111",25163 => "11010000",25164 => "10011010",25165 => "10010010",25166 => "11100111",25167 => "00100010",25168 => "00010101",25169 => "11101001",25170 => "10011001",25171 => "00001111",25172 => "10010100",25173 => "01110110",25174 => "11001010",25175 => "10010101",25176 => "01000010",25177 => "01010110",25178 => "00010110",25179 => "11000100",25180 => "10111010",25181 => "11110011",25182 => "00001100",25183 => "01110110",25184 => "01000000",25185 => "00110001",25186 => "00110111",25187 => "01100111",25188 => "01111100",25189 => "00101010",25190 => "00110101",25191 => "10100010",25192 => "00100000",25193 => "10010000",25194 => "11011011",25195 => "00010000",25196 => "11101010",25197 => "00100100",25198 => "01110010",25199 => "11110100",25200 => "00001111",25201 => "10101010",25202 => "01010001",25203 => "10000011",25204 => "01000010",25205 => "10010101",25206 => "11111010",25207 => "00100111",25208 => "11111001",25209 => "10011011",25210 => "01101100",25211 => "01011001",25212 => "00001011",25213 => "10011100",25214 => "10001111",25215 => "11101001",25216 => "11111011",25217 => "01001111",25218 => "01010101",25219 => "11101100",25220 => "10100011",25221 => "11011000",25222 => "01101010",25223 => "10000101",25224 => "00010111",25225 => "10000110",25226 => "11111101",25227 => "11100011",25228 => "01100011",25229 => "11001010",25230 => "10110001",25231 => "11111001",25232 => "10001110",25233 => "10000110",25234 => "10000101",25235 => "01110001",25236 => "01000010",25237 => "10100101",25238 => "01000001",25239 => "00100111",25240 => "11110101",25241 => "00010000",25242 => "00000010",25243 => "11001101",25244 => "10010001",25245 => "11110100",25246 => "10010011",25247 => "10011010",25248 => "00110011",25249 => "11011000",25250 => "11001111",25251 => "11100111",25252 => "10000000",25253 => "00110011",25254 => "11110110",25255 => "11100001",25256 => "01010000",25257 => "10110100",25258 => "10000100",25259 => "10110000",25260 => "00011100",25261 => "01000111",25262 => "11101101",25263 => "11000100",25264 => "01110011",25265 => "01100110",25266 => "11101001",25267 => "11010001",25268 => "00110010",25269 => "11000110",25270 => "11011000",25271 => "00111001",25272 => "10100111",25273 => "00011010",25274 => "10110111",25275 => "10110110",25276 => "10111110",25277 => "10001111",25278 => "11111101",25279 => "10000000",25280 => "01000001",25281 => "01001001",25282 => "00101111",25283 => "11101010",25284 => "00000110",25285 => "01100011",25286 => "00110011",25287 => "01001101",25288 => "11100111",25289 => "10101001",25290 => "01100100",25291 => "01001001",25292 => "10001110",25293 => "11110100",25294 => "10111100",25295 => "01100000",25296 => "11100101",25297 => "01011100",25298 => "11000011",25299 => "11011100",25300 => "11011010",25301 => "00000111",25302 => "01100111",25303 => "00100110",25304 => "10101001",25305 => "01110110",25306 => "10000001",25307 => "01011101",25308 => "11001110",25309 => "10000010",25310 => "10101010",25311 => "10111111",25312 => "10101011",25313 => "01110101",25314 => "11110110",25315 => "01100110",25316 => "00111011",25317 => "11111001",25318 => "00001010",25319 => "00101100",25320 => "01100000",25321 => "00100010",25322 => "01111011",25323 => "01110001",25324 => "10011110",25325 => "10011110",25326 => "01101011",25327 => "00110101",25328 => "11101001",25329 => "00110010",25330 => "11011001",25331 => "11111000",25332 => "11011010",25333 => "10110110",25334 => "01111000",25335 => "11100101",25336 => "00100111",25337 => "10000101",25338 => "00110110",25339 => "11000000",25340 => "01100111",25341 => "01111100",25342 => "10111000",25343 => "11011001",25344 => "11111001",25345 => "00011100",25346 => "01011111",25347 => "10111000",25348 => "11110110",25349 => "01111110",25350 => "10011011",25351 => "01110111",25352 => "01001001",25353 => "10100001",25354 => "10001000",25355 => "10000101",25356 => "11001100",25357 => "11011000",25358 => "00010011",25359 => "10000101",25360 => "11011110",25361 => "10011101",25362 => "00101111",25363 => "11110101",25364 => "10010111",25365 => "01100000",25366 => "00101001",25367 => "11010101",25368 => "11011111",25369 => "11110110",25370 => "11000101",25371 => "10100001",25372 => "01110111",25373 => "01100101",25374 => "01000110",25375 => "01101100",25376 => "11010100",25377 => "00101010",25378 => "10100011",25379 => "10111101",25380 => "00010110",25381 => "10110110",25382 => "00101100",25383 => "01011010",25384 => "10110100",25385 => "00010111",25386 => "01110110",25387 => "00000101",25388 => "10011000",25389 => "00010010",25390 => "01010001",25391 => "11110011",25392 => "11000011",25393 => "11110101",25394 => "11111101",25395 => "10011110",25396 => "01100111",25397 => "00100111",25398 => "11101000",25399 => "10111111",25400 => "10010110",25401 => "11101011",25402 => "10110111",25403 => "11001101",25404 => "10010011",25405 => "11010000",25406 => "01110101",25407 => "10110100",25408 => "10110110",25409 => "01011111",25410 => "01001010",25411 => "10010100",25412 => "01100111",25413 => "11000010",25414 => "11000100",25415 => "00101100",25416 => "01001001",25417 => "10111001",25418 => "10011101",25419 => "10001111",25420 => "10110001",25421 => "10100011",25422 => "01101001",25423 => "00000011",25424 => "10010000",25425 => "00101011",25426 => "00110111",25427 => "10010010",25428 => "11011111",25429 => "01000110",25430 => "11001011",25431 => "11001000",25432 => "10001101",25433 => "11000110",25434 => "00100101",25435 => "00011010",25436 => "11001011",25437 => "11100010",25438 => "10000001",25439 => "01111111",25440 => "11110101",25441 => "10010111",25442 => "01000000",25443 => "00111110",25444 => "11010101",25445 => "10110011",25446 => "00001110",25447 => "00111010",25448 => "11000000",25449 => "10000001",25450 => "01100010",25451 => "01110101",25452 => "11010001",25453 => "01001101",25454 => "01110001",25455 => "01100111",25456 => "11011010",25457 => "10111011",25458 => "10011000",25459 => "10011011",25460 => "10101111",25461 => "00110110",25462 => "10000101",25463 => "01001001",25464 => "11001101",25465 => "11001101",25466 => "10001001",25467 => "10010100",25468 => "00001000",25469 => "01001001",25470 => "01100011",25471 => "01101110",25472 => "10100111",25473 => "00001101",25474 => "00001111",25475 => "10110111",25476 => "01110000",25477 => "11100111",25478 => "11001001",25479 => "00001000",25480 => "00000101",25481 => "11000100",25482 => "11001111",25483 => "01101001",25484 => "10001100",25485 => "01001110",25486 => "11100001",25487 => "00000101",25488 => "01011010",25489 => "01100010",25490 => "00111100",25491 => "11100001",25492 => "10100001",25493 => "00111100",25494 => "00110010",25495 => "11100100",25496 => "11111111",25497 => "00010111",25498 => "01011001",25499 => "00011101",25500 => "01000111",25501 => "01110100",25502 => "01011001",25503 => "00110101",25504 => "10111000",25505 => "01111000",25506 => "10110111",25507 => "00110001",25508 => "00110110",25509 => "11011001",25510 => "11001010",25511 => "00110111",25512 => "11111100",25513 => "11110111",25514 => "11101101",25515 => "00110011",25516 => "00110101",25517 => "10111101",25518 => "00001111",25519 => "01110011",25520 => "10101101",25521 => "10010110",25522 => "11100000",25523 => "10001011",25524 => "10001010",25525 => "11010000",25526 => "01100111",25527 => "10001101",25528 => "00010010",25529 => "00000101",25530 => "11011000",25531 => "11011100",25532 => "01000111",25533 => "00001100",25534 => "10000010",25535 => "11001000",25536 => "00110010",25537 => "10011100",25538 => "11100000",25539 => "01010010",25540 => "10000011",25541 => "11010001",25542 => "00110000",25543 => "00101110",25544 => "11010011",25545 => "01100110",25546 => "01010010",25547 => "00111001",25548 => "11011100",25549 => "00011100",25550 => "00000010",25551 => "11100011",25552 => "11110111",25553 => "10100101",25554 => "10011100",25555 => "10101001",25556 => "00001111",25557 => "10010010",25558 => "00010001",25559 => "10010101",25560 => "01101110",25561 => "01101111",25562 => "00001001",25563 => "10100010",25564 => "00000101",25565 => "10011001",25566 => "11001010",25567 => "10101010",25568 => "10010011",25569 => "11100111",25570 => "11001011",25571 => "11000111",25572 => "00100101",25573 => "10000011",25574 => "11011001",25575 => "00000101",25576 => "11110111",25577 => "00010000",25578 => "01011011",25579 => "01001110",25580 => "00001000",25581 => "11111001",25582 => "01111101",25583 => "01110110",25584 => "01101101",25585 => "10010111",25586 => "11111110",25587 => "10011111",25588 => "01101000",25589 => "01101010",25590 => "00101110",25591 => "00001111",25592 => "01110000",25593 => "10011100",25594 => "00110001",25595 => "01011000",25596 => "01010000",25597 => "01110010",25598 => "10000101",25599 => "00011110",25600 => "01110101",25601 => "11101111",25602 => "00010110",25603 => "00001001",25604 => "00011110",25605 => "11110110",25606 => "01100010",25607 => "10100001",25608 => "01111111",25609 => "11101101",25610 => "00000001",25611 => "00000001",25612 => "00010000",25613 => "11001010",25614 => "11001010",25615 => "11101101",25616 => "00110001",25617 => "10011101",25618 => "01101110",25619 => "01101000",25620 => "00010111",25621 => "00100011",25622 => "10001000",25623 => "11001110",25624 => "11000001",25625 => "10101011",25626 => "00010010",25627 => "11001100",25628 => "10100110",25629 => "10010001",25630 => "00111110",25631 => "00001111",25632 => "00011110",25633 => "01011010",25634 => "00000000",25635 => "00101011",25636 => "11010011",25637 => "00011100",25638 => "11101100",25639 => "01111011",25640 => "11001100",25641 => "01101000",25642 => "10100110",25643 => "00110100",25644 => "11100111",25645 => "11100111",25646 => "01110111",25647 => "10100001",25648 => "01010110",25649 => "10011001",25650 => "11010001",25651 => "10101010",25652 => "01000011",25653 => "00100111",25654 => "10001001",25655 => "10000010",25656 => "11110001",25657 => "11001010",25658 => "00000111",25659 => "00000011",25660 => "00110101",25661 => "11010111",25662 => "11110010",25663 => "10110101",25664 => "11100010",25665 => "10100111",25666 => "11000101",25667 => "10100000",25668 => "11011010",25669 => "01001000",25670 => "11110000",25671 => "10000111",25672 => "00101000",25673 => "01110010",25674 => "01100111",25675 => "10100100",25676 => "10111101",25677 => "00011000",25678 => "11001110",25679 => "10111010",25680 => "00011111",25681 => "01100111",25682 => "11100010",25683 => "11111100",25684 => "10100001",25685 => "10110110",25686 => "01011010",25687 => "00000101",25688 => "11111010",25689 => "00011000",25690 => "11100100",25691 => "00010100",25692 => "10011111",25693 => "10001000",25694 => "10111000",25695 => "10100110",25696 => "10100001",25697 => "11010110",25698 => "01010101",25699 => "10001001",25700 => "00000100",25701 => "00110000",25702 => "00111110",25703 => "10000100",25704 => "00111111",25705 => "10001001",25706 => "11100111",25707 => "10100101",25708 => "01001000",25709 => "01101101",25710 => "00110000",25711 => "01100100",25712 => "00010011",25713 => "10110101",25714 => "01101011",25715 => "11111001",25716 => "11010111",25717 => "11000000",25718 => "11010111",25719 => "10000111",25720 => "10101011",25721 => "00110111",25722 => "11000010",25723 => "11100010",25724 => "00001111",25725 => "01100101",25726 => "01001011",25727 => "00011110",25728 => "01111011",25729 => "11001101",25730 => "10101000",25731 => "00001100",25732 => "10100110",25733 => "00010110",25734 => "10010000",25735 => "00110110",25736 => "10111101",25737 => "01011010",25738 => "10010010",25739 => "00000000",25740 => "01010000",25741 => "11111101",25742 => "00011001",25743 => "01110000",25744 => "11010110",25745 => "00101010",25746 => "01110111",25747 => "11010000",25748 => "00100111",25749 => "11001010",25750 => "11111101",25751 => "10100001",25752 => "11010110",25753 => "10100110",25754 => "11100011",25755 => "10101110",25756 => "10011001",25757 => "01000111",25758 => "01111000",25759 => "00011110",25760 => "10100111",25761 => "10010000",25762 => "10110101",25763 => "01100110",25764 => "01011011",25765 => "10001001",25766 => "11000111",25767 => "11011110",25768 => "10110010",25769 => "11000110",25770 => "11010100",25771 => "11000100",25772 => "10011110",25773 => "10000110",25774 => "11111000",25775 => "01110010",25776 => "00100011",25777 => "00001000",25778 => "11110110",25779 => "10111100",25780 => "11101001",25781 => "01011001",25782 => "00001101",25783 => "11111000",25784 => "11100100",25785 => "11101000",25786 => "10000001",25787 => "00111101",25788 => "00111010",25789 => "01101110",25790 => "01010101",25791 => "00000111",25792 => "01010110",25793 => "01110110",25794 => "01011001",25795 => "11111011",25796 => "11101100",25797 => "00111000",25798 => "10111110",25799 => "01001010",25800 => "10101000",25801 => "00000111",25802 => "01000010",25803 => "11011111",25804 => "10101110",25805 => "10010000",25806 => "01001100",25807 => "01100000",25808 => "11000110",25809 => "01011111",25810 => "01111110",25811 => "01111010",25812 => "00001101",25813 => "00110010",25814 => "10011000",25815 => "01000110",25816 => "11100110",25817 => "10001010",25818 => "00100111",25819 => "00010000",25820 => "00100100",25821 => "10011111",25822 => "10111110",25823 => "11101011",25824 => "00011101",25825 => "11111100",25826 => "11000001",25827 => "00100001",25828 => "01011111",25829 => "10111000",25830 => "00110101",25831 => "10110011",25832 => "10101011",25833 => "10011000",25834 => "11100000",25835 => "11111011",25836 => "11100001",25837 => "00000100",25838 => "01001000",25839 => "00000110",25840 => "10001011",25841 => "11000101",25842 => "11110000",25843 => "10011100",25844 => "01111010",25845 => "01110100",25846 => "00011000",25847 => "11111000",25848 => "10101000",25849 => "00000001",25850 => "10100110",25851 => "00001100",25852 => "11101100",25853 => "10000000",25854 => "11011100",25855 => "01110101",25856 => "01000100",25857 => "00010100",25858 => "11100111",25859 => "11111110",25860 => "11001110",25861 => "00011111",25862 => "10010101",25863 => "00010100",25864 => "01011010",25865 => "10010001",25866 => "01001010",25867 => "00101110",25868 => "00001011",25869 => "00001000",25870 => "01111100",25871 => "11100101",25872 => "00000011",25873 => "01111011",25874 => "11000111",25875 => "10110010",25876 => "01010000",25877 => "10111011",25878 => "10101110",25879 => "10010011",25880 => "01101000",25881 => "00001001",25882 => "01110100",25883 => "11101010",25884 => "10000100",25885 => "01110110",25886 => "00000111",25887 => "11100000",25888 => "00011101",25889 => "00011100",25890 => "11011011",25891 => "11100010",25892 => "10101010",25893 => "11101011",25894 => "00101110",25895 => "11001111",25896 => "00000001",25897 => "11101110",25898 => "10000011",25899 => "10011011",25900 => "10110111",25901 => "11011001",25902 => "01000100",25903 => "00111001",25904 => "00111111",25905 => "01000100",25906 => "00001011",25907 => "00110100",25908 => "00110001",25909 => "01101001",25910 => "00010010",25911 => "11100011",25912 => "11010110",25913 => "11111000",25914 => "01011010",25915 => "01000001",25916 => "00110001",25917 => "11110111",25918 => "10001110",25919 => "10101100",25920 => "01010000",25921 => "01100110",25922 => "01010011",25923 => "01100110",25924 => "00110010",25925 => "11010011",25926 => "10111101",25927 => "00000000",25928 => "10110101",25929 => "00001011",25930 => "10101000",25931 => "01110000",25932 => "10110011",25933 => "10101110",25934 => "10000101",25935 => "01111011",25936 => "00001001",25937 => "00010011",25938 => "10010000",25939 => "11000111",25940 => "00010110",25941 => "10110100",25942 => "00010000",25943 => "10111011",25944 => "10011110",25945 => "10100101",25946 => "11111110",25947 => "01001110",25948 => "01111100",25949 => "01010001",25950 => "11101010",25951 => "00111001",25952 => "11101110",25953 => "00010000",25954 => "00000010",25955 => "10100100",25956 => "11011000",25957 => "00001110",25958 => "00011000",25959 => "11101000",25960 => "11110000",25961 => "01101110",25962 => "01011000",25963 => "10010000",25964 => "01000100",25965 => "11011001",25966 => "11001011",25967 => "01010101",25968 => "11100000",25969 => "11011000",25970 => "01111110",25971 => "10011100",25972 => "00101101",25973 => "00001000",25974 => "01101111",25975 => "10100101",25976 => "10111111",25977 => "11000111",25978 => "11100101",25979 => "01101011",25980 => "11111000",25981 => "10000001",25982 => "00111101",25983 => "11011000",25984 => "10100111",25985 => "11001101",25986 => "00100100",25987 => "11101111",25988 => "11001001",25989 => "10101100",25990 => "00100100",25991 => "01010100",25992 => "00000101",25993 => "00000011",25994 => "01001010",25995 => "10100110",25996 => "00001100",25997 => "11100010",25998 => "00011000",25999 => "11011111",26000 => "11001110",26001 => "10101100",26002 => "11100111",26003 => "10011111",26004 => "11110101",26005 => "10100100",26006 => "00101001",26007 => "11111110",26008 => "10111001",26009 => "10000100",26010 => "00010000",26011 => "01000101",26012 => "11011110",26013 => "01001100",26014 => "01001000",26015 => "01100011",26016 => "01000111",26017 => "01100000",26018 => "00100000",26019 => "10111100",26020 => "10111100",26021 => "00100100",26022 => "00100111",26023 => "10000000",26024 => "00110101",26025 => "01011010",26026 => "00001001",26027 => "01010010",26028 => "10110110",26029 => "01010101",26030 => "01000111",26031 => "10010100",26032 => "01100100",26033 => "11011011",26034 => "10001110",26035 => "01010010",26036 => "01101101",26037 => "01111011",26038 => "01111101",26039 => "11111100",26040 => "00000001",26041 => "11100001",26042 => "11011110",26043 => "01010000",26044 => "00101111",26045 => "10001000",26046 => "00100110",26047 => "11111110",26048 => "11010110",26049 => "00110110",26050 => "01110000",26051 => "00110000",26052 => "00010010",26053 => "01111000",26054 => "00101110",26055 => "11010001",26056 => "10001010",26057 => "00001001",26058 => "11100110",26059 => "01000101",26060 => "01101011",26061 => "11111100",26062 => "00101101",26063 => "00010010",26064 => "01111111",26065 => "10111110",26066 => "01010100",26067 => "11111001",26068 => "00100010",26069 => "00100110",26070 => "11100001",26071 => "10111000",26072 => "00111000",26073 => "10000111",26074 => "11100101",26075 => "11110000",26076 => "10000100",26077 => "11011000",26078 => "10000100",26079 => "01000001",26080 => "11111101",26081 => "01011100",26082 => "00100100",26083 => "00101100",26084 => "00111100",26085 => "01100110",26086 => "11011010",26087 => "01101001",26088 => "11010000",26089 => "11101101",26090 => "01110001",26091 => "01000000",26092 => "11110010",26093 => "10100010",26094 => "00011100",26095 => "11111001",26096 => "01110101",26097 => "01101100",26098 => "01000110",26099 => "01011110",26100 => "00101101",26101 => "11111100",26102 => "11101110",26103 => "11110000",26104 => "10000110",26105 => "10001111",26106 => "01011001",26107 => "01010100",26108 => "11111100",26109 => "01011000",26110 => "10000111",26111 => "01000100",26112 => "00110100",26113 => "00000110",26114 => "11101010",26115 => "00000110",26116 => "10101011",26117 => "11111100",26118 => "10000101",26119 => "01001110",26120 => "01001110",26121 => "11001011",26122 => "01101111",26123 => "00100010",26124 => "01110101",26125 => "00101110",26126 => "00101001",26127 => "11000001",26128 => "11001110",26129 => "01001100",26130 => "00011101",26131 => "10100010",26132 => "01010001",26133 => "00000111",26134 => "11011011",26135 => "11100010",26136 => "10010110",26137 => "00111101",26138 => "00010111",26139 => "01011100",26140 => "11111011",26141 => "11101101",26142 => "11101101",26143 => "10111001",26144 => "11001100",26145 => "00100111",26146 => "00010111",26147 => "11100010",26148 => "01010101",26149 => "11001111",26150 => "01000100",26151 => "00100101",26152 => "11010011",26153 => "01010110",26154 => "01000101",26155 => "11000011",26156 => "01111111",26157 => "01010011",26158 => "10010011",26159 => "10100010",26160 => "01011100",26161 => "00001111",26162 => "10011100",26163 => "11101110",26164 => "00001001",26165 => "01100011",26166 => "01111011",26167 => "10010001",26168 => "01111010",26169 => "01101000",26170 => "01111001",26171 => "01000001",26172 => "00100001",26173 => "11100000",26174 => "00001111",26175 => "10110100",26176 => "01100110",26177 => "01101011",26178 => "00011100",26179 => "00111100",26180 => "10100101",26181 => "11010010",26182 => "01000100",26183 => "00111010",26184 => "00111001",26185 => "00111000",26186 => "01011011",26187 => "01011000",26188 => "00100011",26189 => "10101000",26190 => "10011111",26191 => "10000001",26192 => "11010011",26193 => "00111110",26194 => "00111011",26195 => "01111011",26196 => "11110111",26197 => "10001101",26198 => "01010110",26199 => "10101110",26200 => "00011010",26201 => "11101010",26202 => "01011111",26203 => "01011001",26204 => "11100101",26205 => "11101001",26206 => "01100010",26207 => "11101011",26208 => "11110101",26209 => "01111011",26210 => "10010010",26211 => "10000001",26212 => "01000011",26213 => "01011110",26214 => "00010000",26215 => "11111010",26216 => "01101110",26217 => "10100110",26218 => "10110010",26219 => "10110010",26220 => "01100011",26221 => "10001010",26222 => "11111110",26223 => "11011110",26224 => "10110000",26225 => "11110010",26226 => "10000100",26227 => "01000100",26228 => "01101100",26229 => "01100100",26230 => "00011101",26231 => "10101011",26232 => "11110011",26233 => "01111011",26234 => "11011011",26235 => "01011010",26236 => "11111110",26237 => "11000100",26238 => "01111110",26239 => "01110001",26240 => "01010101",26241 => "10100100",26242 => "00110000",26243 => "00011111",26244 => "10101101",26245 => "00010000",26246 => "11010010",26247 => "10110000",26248 => "10110110",26249 => "00110110",26250 => "10111001",26251 => "11101101",26252 => "01101011",26253 => "10101010",26254 => "00001100",26255 => "00111010",26256 => "01001010",26257 => "11011011",26258 => "11001011",26259 => "00100101",26260 => "00101000",26261 => "10010011",26262 => "01100110",26263 => "10000011",26264 => "10001100",26265 => "11110000",26266 => "00000010",26267 => "11100100",26268 => "01001111",26269 => "00100100",26270 => "11001100",26271 => "11101011",26272 => "11011110",26273 => "10100001",26274 => "10110000",26275 => "01111101",26276 => "01000001",26277 => "10111011",26278 => "00011111",26279 => "00110110",26280 => "01000110",26281 => "11100110",26282 => "01101000",26283 => "10010000",26284 => "11001110",26285 => "11100000",26286 => "00101111",26287 => "11011011",26288 => "01000111",26289 => "10101111",26290 => "00101101",26291 => "10100101",26292 => "01101000",26293 => "11010011",26294 => "00010001",26295 => "00000000",26296 => "01110000",26297 => "00101101",26298 => "11000010",26299 => "10010001",26300 => "11001111",26301 => "11101010",26302 => "11000000",26303 => "01011110",26304 => "01110111",26305 => "00001010",26306 => "11001011",26307 => "01000000",26308 => "01010010",26309 => "01111001",26310 => "10110011",26311 => "00101100",26312 => "00100101",26313 => "00101001",26314 => "00011111",26315 => "01100110",26316 => "00110000",26317 => "10101101",26318 => "11100101",26319 => "11101101",26320 => "00111010",26321 => "01011011",26322 => "01110100",26323 => "11001000",26324 => "01111110",26325 => "01111011",26326 => "11010010",26327 => "11100010",26328 => "11101111",26329 => "00100011",26330 => "01100011",26331 => "00101100",26332 => "11110001",26333 => "01111011",26334 => "10100011",26335 => "01001110",26336 => "11011001",26337 => "10100001",26338 => "10011110",26339 => "00010101",26340 => "10000110",26341 => "01010100",26342 => "01001110",26343 => "11111010",26344 => "00110111",26345 => "01100100",26346 => "01110101",26347 => "01100010",26348 => "10101111",26349 => "11101100",26350 => "11110110",26351 => "00110100",26352 => "00000001",26353 => "10100110",26354 => "11111010",26355 => "01011000",26356 => "00111101",26357 => "10111111",26358 => "00011001",26359 => "00000100",26360 => "10101010",26361 => "01110110",26362 => "10100000",26363 => "10100011",26364 => "00100101",26365 => "00001111",26366 => "00011111",26367 => "00010110",26368 => "01111011",26369 => "00101111",26370 => "11011110",26371 => "11110000",26372 => "11000111",26373 => "01101100",26374 => "00110011",26375 => "10011001",26376 => "11010001",26377 => "00011110",26378 => "00101100",26379 => "11011111",26380 => "01011101",26381 => "10001110",26382 => "01111110",26383 => "11111001",26384 => "00111000",26385 => "01011011",26386 => "01010011",26387 => "11100010",26388 => "10101111",26389 => "10100011",26390 => "00110000",26391 => "10111000",26392 => "00100010",26393 => "00010010",26394 => "10000000",26395 => "10111010",26396 => "11101110",26397 => "01100000",26398 => "10010111",26399 => "00000001",26400 => "01100110",26401 => "10000011",26402 => "10001010",26403 => "10011101",26404 => "00000100",26405 => "10100111",26406 => "11001011",26407 => "10100011",26408 => "11100101",26409 => "10110110",26410 => "01111110",26411 => "11110101",26412 => "00100110",26413 => "00110100",26414 => "11110110",26415 => "10100010",26416 => "00111001",26417 => "11110100",26418 => "01010111",26419 => "01100000",26420 => "10011111",26421 => "11011000",26422 => "11011110",26423 => "00111110",26424 => "00000101",26425 => "11001001",26426 => "10011011",26427 => "01000000",26428 => "00101011",26429 => "00101001",26430 => "00100101",26431 => "00100000",26432 => "10001000",26433 => "01100111",26434 => "11100010",26435 => "01001000",26436 => "11100000",26437 => "01001011",26438 => "11001011",26439 => "10011011",26440 => "10000110",26441 => "01100011",26442 => "10011111",26443 => "00010010",26444 => "01001100",26445 => "01000011",26446 => "10001010",26447 => "00101110",26448 => "01011010",26449 => "11101011",26450 => "00011011",26451 => "10011110",26452 => "10010011",26453 => "11010001",26454 => "10111001",26455 => "10100111",26456 => "10001000",26457 => "11110000",26458 => "01100101",26459 => "11111011",26460 => "10011100",26461 => "01110001",26462 => "00110011",26463 => "10011100",26464 => "11011000",26465 => "00111111",26466 => "11000111",26467 => "11101000",26468 => "01101111",26469 => "11100010",26470 => "11010000",26471 => "01100010",26472 => "00011010",26473 => "00001001",26474 => "11000111",26475 => "01100010",26476 => "11100010",26477 => "10011100",26478 => "00101110",26479 => "00100010",26480 => "01110111",26481 => "00011110",26482 => "01010010",26483 => "01110011",26484 => "10110001",26485 => "00101111",26486 => "01011010",26487 => "11000011",26488 => "01001010",26489 => "01000000",26490 => "11001101",26491 => "01100011",26492 => "10111111",26493 => "01010110",26494 => "10101001",26495 => "10101011",26496 => "10000011",26497 => "00101000",26498 => "11110111",26499 => "00010110",26500 => "11111011",26501 => "10011010",26502 => "00101010",26503 => "10111000",26504 => "01110110",26505 => "10100111",26506 => "11111010",26507 => "00101111",26508 => "11010101",26509 => "01000000",26510 => "00010110",26511 => "10100100",26512 => "01010000",26513 => "00000111",26514 => "11100001",26515 => "01000101",26516 => "00100010",26517 => "10001110",26518 => "01001000",26519 => "01001101",26520 => "01111110",26521 => "11101000",26522 => "00100000",26523 => "00111001",26524 => "01100101",26525 => "11111001",26526 => "11100101",26527 => "10011001",26528 => "10011111",26529 => "01010111",26530 => "11001101",26531 => "01000100",26532 => "11001001",26533 => "00011011",26534 => "01010100",26535 => "11011001",26536 => "01011000",26537 => "10110011",26538 => "10001101",26539 => "10010100",26540 => "00111000",26541 => "10101100",26542 => "01001111",26543 => "11000001",26544 => "10110101",26545 => "11000100",26546 => "11101000",26547 => "11001111",26548 => "11001000",26549 => "10000001",26550 => "00011101",26551 => "00110001",26552 => "11100101",26553 => "11101101",26554 => "00101001",26555 => "00100000",26556 => "11100111",26557 => "01011000",26558 => "10101000",26559 => "01111110",26560 => "01000011",26561 => "01111101",26562 => "00111000",26563 => "10100011",26564 => "11110010",26565 => "01000000",26566 => "10011010",26567 => "01010111",26568 => "11010010",26569 => "00100001",26570 => "01001011",26571 => "00010111",26572 => "10000011",26573 => "11111100",26574 => "10110001",26575 => "00000111",26576 => "11101001",26577 => "11100000",26578 => "01001101",26579 => "10011011",26580 => "00011111",26581 => "00111110",26582 => "11001011",26583 => "11111000",26584 => "00010101",26585 => "01001100",26586 => "10000001",26587 => "00010100",26588 => "10010010",26589 => "00100100",26590 => "10010111",26591 => "01110111",26592 => "10011001",26593 => "11110001",26594 => "10100001",26595 => "00100101",26596 => "00011100",26597 => "01000011",26598 => "11100111",26599 => "11011101",26600 => "01100011",26601 => "00000100",26602 => "11110101",26603 => "10100001",26604 => "01100101",26605 => "11001100",26606 => "01000010",26607 => "00110001",26608 => "10100100",26609 => "01100001",26610 => "00011010",26611 => "10001100",26612 => "00110100",26613 => "01000001",26614 => "00000010",26615 => "01101000",26616 => "01111001",26617 => "11100011",26618 => "11001101",26619 => "10110111",26620 => "01101100",26621 => "11100111",26622 => "10110011",26623 => "00011111",26624 => "10001110",26625 => "01011000",26626 => "00111001",26627 => "10001110",26628 => "11001110",26629 => "10011110",26630 => "11100001",26631 => "01110010",26632 => "00000010",26633 => "00101110",26634 => "11101111",26635 => "00011100",26636 => "01010001",26637 => "10001110",26638 => "01000010",26639 => "00000000",26640 => "10111011",26641 => "00010111",26642 => "01000010",26643 => "10000110",26644 => "10101100",26645 => "10110101",26646 => "00101010",26647 => "10100111",26648 => "10011101",26649 => "01100101",26650 => "11000101",26651 => "01000010",26652 => "11110100",26653 => "01010000",26654 => "01011110",26655 => "10110010",26656 => "01011000",26657 => "11100110",26658 => "10110011",26659 => "11110100",26660 => "11111001",26661 => "11000001",26662 => "10100101",26663 => "10010011",26664 => "01111100",26665 => "11100100",26666 => "11001101",26667 => "01000110",26668 => "00001110",26669 => "00100000",26670 => "01100101",26671 => "01011110",26672 => "01010111",26673 => "01111100",26674 => "01011111",26675 => "10001000",26676 => "11101110",26677 => "10000010",26678 => "01110100",26679 => "00010101",26680 => "00000001",26681 => "10110011",26682 => "00101010",26683 => "00011010",26684 => "11010101",26685 => "01101000",26686 => "01001000",26687 => "11011110",26688 => "00011111",26689 => "10000000",26690 => "00111111",26691 => "10001010",26692 => "01100110",26693 => "00000110",26694 => "11011011",26695 => "01101110",26696 => "11101000",26697 => "00011000",26698 => "01100110",26699 => "10000111",26700 => "11111011",26701 => "11101011",26702 => "11101001",26703 => "01011101",26704 => "01100001",26705 => "10001010",26706 => "01011000",26707 => "01000100",26708 => "11001101",26709 => "10100000",26710 => "11010010",26711 => "01100110",26712 => "11000000",26713 => "11111111",26714 => "00100011",26715 => "00010010",26716 => "01100011",26717 => "10011001",26718 => "01110110",26719 => "01100100",26720 => "00011001",26721 => "01100100",26722 => "11100011",26723 => "00111110",26724 => "11101101",26725 => "10111110",26726 => "11010010",26727 => "01000101",26728 => "11011100",26729 => "11011010",26730 => "11100100",26731 => "01010100",26732 => "00010011",26733 => "10011001",26734 => "01111010",26735 => "10000001",26736 => "10011110",26737 => "11001001",26738 => "11110111",26739 => "11111111",26740 => "01011000",26741 => "11011101",26742 => "10010000",26743 => "01100000",26744 => "10100000",26745 => "10010000",26746 => "01011110",26747 => "01001111",26748 => "01011011",26749 => "10100000",26750 => "01111011",26751 => "10101001",26752 => "01110100",26753 => "10010101",26754 => "11110000",26755 => "11010001",26756 => "11000110",26757 => "00011100",26758 => "11010010",26759 => "01111011",26760 => "01011010",26761 => "00101011",26762 => "11001011",26763 => "10110010",26764 => "00110101",26765 => "11101001",26766 => "00010101",26767 => "01001110",26768 => "01100110",26769 => "00000101",26770 => "01000001",26771 => "00011101",26772 => "00100101",26773 => "11101010",26774 => "00100000",26775 => "01001010",26776 => "10101001",26777 => "00101001",26778 => "00101100",26779 => "11110100",26780 => "10001010",26781 => "11000010",26782 => "10101001",26783 => "00111001",26784 => "10111010",26785 => "01001101",26786 => "11110110",26787 => "10000011",26788 => "10011001",26789 => "11010010",26790 => "01101001",26791 => "10010000",26792 => "01101011",26793 => "01000010",26794 => "00100001",26795 => "11110011",26796 => "11001011",26797 => "00101111",26798 => "01011100",26799 => "10001011",26800 => "10111000",26801 => "11100110",26802 => "11011001",26803 => "10100001",26804 => "10101000",26805 => "01001010",26806 => "11011001",26807 => "00100101",26808 => "11101011",26809 => "11001100",26810 => "00010000",26811 => "01011101",26812 => "00110101",26813 => "00001011",26814 => "10111011",26815 => "01011011",26816 => "11010001",26817 => "00110010",26818 => "00110111",26819 => "01000011",26820 => "01001101",26821 => "00001010",26822 => "11000010",26823 => "10011101",26824 => "01100110",26825 => "00011111",26826 => "10110110",26827 => "00100110",26828 => "10101001",26829 => "00001000",26830 => "10100111",26831 => "01010100",26832 => "10011110",26833 => "01010100",26834 => "10000011",26835 => "00110011",26836 => "01100101",26837 => "00100100",26838 => "11011011",26839 => "01010000",26840 => "00011110",26841 => "00100101",26842 => "00101000",26843 => "11011101",26844 => "01110011",26845 => "11010001",26846 => "11010101",26847 => "00000100",26848 => "11111101",26849 => "11011111",26850 => "11101010",26851 => "11111110",26852 => "01110011",26853 => "00001100",26854 => "10100110",26855 => "10001011",26856 => "01010101",26857 => "01010100",26858 => "10110011",26859 => "00100001",26860 => "01110100",26861 => "01111000",26862 => "00100010",26863 => "11100000",26864 => "00001000",26865 => "00001001",26866 => "00000101",26867 => "10110010",26868 => "11101101",26869 => "11001011",26870 => "11011000",26871 => "10011010",26872 => "11101000",26873 => "01001000",26874 => "11111110",26875 => "10001010",26876 => "01101110",26877 => "11001011",26878 => "01101011",26879 => "11011111",26880 => "00111110",26881 => "11100011",26882 => "00001100",26883 => "00011101",26884 => "01110110",26885 => "01110010",26886 => "00001000",26887 => "00110001",26888 => "10001100",26889 => "01001000",26890 => "11010100",26891 => "10100010",26892 => "11100101",26893 => "01110010",26894 => "01101011",26895 => "00000111",26896 => "10000000",26897 => "10011111",26898 => "00000111",26899 => "10111101",26900 => "10110111",26901 => "01001111",26902 => "11111111",26903 => "10001101",26904 => "01010100",26905 => "01111010",26906 => "00111001",26907 => "01100100",26908 => "00111011",26909 => "10001111",26910 => "01100110",26911 => "01100110",26912 => "11011101",26913 => "00000010",26914 => "01001110",26915 => "00111100",26916 => "01101100",26917 => "00100100",26918 => "11101000",26919 => "01011001",26920 => "00010100",26921 => "11100110",26922 => "11010111",26923 => "11000101",26924 => "10000000",26925 => "00100110",26926 => "11011101",26927 => "00101100",26928 => "11010101",26929 => "10010001",26930 => "10110001",26931 => "10111111",26932 => "00101110",26933 => "01000011",26934 => "00010001",26935 => "01111011",26936 => "11011100",26937 => "10111001",26938 => "10100110",26939 => "11100001",26940 => "01100001",26941 => "11010110",26942 => "00111111",26943 => "01001100",26944 => "01101100",26945 => "00001000",26946 => "00000011",26947 => "00010011",26948 => "01011011",26949 => "10001110",26950 => "01001011",26951 => "01111100",26952 => "00100110",26953 => "00100110",26954 => "00010001",26955 => "11111110",26956 => "11110101",26957 => "10000110",26958 => "00110001",26959 => "01110110",26960 => "10111110",26961 => "00010001",26962 => "10100100",26963 => "11101110",26964 => "00100110",26965 => "11011011",26966 => "11000110",26967 => "00100011",26968 => "10001001",26969 => "11101111",26970 => "10000101",26971 => "00011010",26972 => "00011100",26973 => "10100111",26974 => "10000110",26975 => "01001011",26976 => "01111100",26977 => "11010101",26978 => "10000001",26979 => "01001000",26980 => "00000111",26981 => "01011010",26982 => "01101000",26983 => "01010010",26984 => "11100011",26985 => "10100001",26986 => "01111000",26987 => "00001100",26988 => "10001110",26989 => "10100011",26990 => "10100011",26991 => "01110111",26992 => "01000101",26993 => "01010100",26994 => "01000101",26995 => "11111110",26996 => "10011010",26997 => "01111001",26998 => "00101100",26999 => "11111000",27000 => "00101011",27001 => "11111000",27002 => "01110001",27003 => "11001001",27004 => "01101110",27005 => "00101111",27006 => "00000001",27007 => "10001000",27008 => "00100010",27009 => "01100000",27010 => "10100100",27011 => "11001101",27012 => "00100100",27013 => "01100101",27014 => "00001101",27015 => "01101101",27016 => "11101010",27017 => "00100011",27018 => "10110101",27019 => "00101001",27020 => "11010001",27021 => "11001101",27022 => "00011111",27023 => "10001011",27024 => "01001111",27025 => "11100100",27026 => "10000000",27027 => "01010000",27028 => "01001000",27029 => "10010111",27030 => "00001100",27031 => "00011010",27032 => "01001000",27033 => "10111010",27034 => "00000100",27035 => "11111101",27036 => "10011100",27037 => "10110010",27038 => "10010000",27039 => "10001101",27040 => "11011111",27041 => "00011000",27042 => "01011010",27043 => "10000101",27044 => "00010000",27045 => "10001001",27046 => "01010111",27047 => "10011001",27048 => "10010101",27049 => "00010001",27050 => "01010100",27051 => "00110010",27052 => "11110010",27053 => "11001100",27054 => "00100011",27055 => "10010000",27056 => "11001101",27057 => "01110010",27058 => "00100001",27059 => "00000000",27060 => "00011111",27061 => "00000010",27062 => "01011011",27063 => "10011010",27064 => "10101100",27065 => "00100010",27066 => "01100011",27067 => "01011110",27068 => "11011111",27069 => "00110010",27070 => "01110001",27071 => "10010100",27072 => "10011101",27073 => "01111111",27074 => "11100000",27075 => "01000010",27076 => "10010100",27077 => "00001001",27078 => "01010010",27079 => "00000110",27080 => "10101011",27081 => "00111100",27082 => "00111011",27083 => "01011100",27084 => "11001101",27085 => "00100111",27086 => "01100100",27087 => "00101001",27088 => "11110101",27089 => "00100101",27090 => "11010111",27091 => "01101011",27092 => "10101110",27093 => "11110010",27094 => "10001110",27095 => "01001100",27096 => "01100000",27097 => "11010110",27098 => "10101011",27099 => "11001000",27100 => "00111000",27101 => "11000001",27102 => "00001010",27103 => "11100100",27104 => "11001000",27105 => "11110000",27106 => "01011011",27107 => "11011111",27108 => "10111111",27109 => "01111010",27110 => "01010011",27111 => "01101001",27112 => "10111101",27113 => "01011010",27114 => "10011111",27115 => "00010110",27116 => "10001110",27117 => "11010101",27118 => "11110011",27119 => "00100001",27120 => "11110011",27121 => "11110011",27122 => "10011011",27123 => "01100000",27124 => "00010101",27125 => "01111111",27126 => "11111011",27127 => "10001000",27128 => "01101100",27129 => "10011010",27130 => "10011101",27131 => "11001100",27132 => "11000011",27133 => "01101010",27134 => "00010110",27135 => "11110001",27136 => "11011111",27137 => "01000001",27138 => "10111011",27139 => "11001110",27140 => "11111001",27141 => "01001000",27142 => "11100110",27143 => "10010001",27144 => "00000010",27145 => "01101011",27146 => "00010110",27147 => "01110100",27148 => "00111010",27149 => "10110111",27150 => "00100111",27151 => "01001100",27152 => "01010110",27153 => "01001001",27154 => "11000010",27155 => "10010000",27156 => "10111100",27157 => "01001101",27158 => "10111100",27159 => "10110010",27160 => "11000001",27161 => "10000001",27162 => "01001010",27163 => "10010001",27164 => "00110001",27165 => "00010011",27166 => "11010001",27167 => "11111101",27168 => "00110010",27169 => "01100001",27170 => "00110101",27171 => "10110001",27172 => "00101001",27173 => "11101000",27174 => "10000101",27175 => "01011010",27176 => "11010100",27177 => "11101001",27178 => "10100010",27179 => "00011100",27180 => "11100100",27181 => "00111011",27182 => "10111111",27183 => "01010000",27184 => "11110011",27185 => "00111110",27186 => "11110111",27187 => "01001110",27188 => "11111001",27189 => "01101110",27190 => "01011010",27191 => "11000001",27192 => "10001010",27193 => "11110000",27194 => "10110110",27195 => "10101110",27196 => "00011101",27197 => "00010001",27198 => "10111001",27199 => "10010100",27200 => "00010111",27201 => "10001100",27202 => "01000011",27203 => "10011111",27204 => "10000000",27205 => "10100000",27206 => "10101111",27207 => "11011011",27208 => "11010001",27209 => "01001110",27210 => "10110001",27211 => "10111110",27212 => "01101100",27213 => "01101001",27214 => "10100001",27215 => "10010101",27216 => "10011010",27217 => "01001101",27218 => "11011011",27219 => "11001111",27220 => "10100101",27221 => "10000011",27222 => "00011001",27223 => "11000100",27224 => "11011111",27225 => "01011001",27226 => "10010110",27227 => "11101101",27228 => "01101111",27229 => "01100010",27230 => "01111010",27231 => "10001111",27232 => "00001101",27233 => "00110010",27234 => "00110111",27235 => "01101000",27236 => "11111010",27237 => "11110111",27238 => "00111010",27239 => "11001001",27240 => "00011110",27241 => "10011011",27242 => "00011011",27243 => "00100000",27244 => "11101101",27245 => "10010010",27246 => "01000000",27247 => "11111111",27248 => "01011100",27249 => "11101100",27250 => "11101000",27251 => "00001110",27252 => "01001001",27253 => "10000001",27254 => "01110010",27255 => "00111110",27256 => "10101101",27257 => "01001011",27258 => "01011011",27259 => "11011011",27260 => "10101000",27261 => "01101101",27262 => "11011001",27263 => "11100001",27264 => "01110010",27265 => "01011001",27266 => "11000001",27267 => "00100000",27268 => "10011010",27269 => "10111001",27270 => "01010010",27271 => "00100111",27272 => "10110101",27273 => "11101100",27274 => "01010000",27275 => "10110011",27276 => "00000011",27277 => "01011010",27278 => "11101001",27279 => "11100101",27280 => "11000111",27281 => "11010100",27282 => "11111100",27283 => "11000111",27284 => "00110101",27285 => "11100010",27286 => "11000100",27287 => "10110111",27288 => "10000110",27289 => "10111011",27290 => "11101101",27291 => "11111000",27292 => "01100110",27293 => "01100111",27294 => "01011101",27295 => "10110100",27296 => "11000111",27297 => "00100011",27298 => "11001000",27299 => "10011100",27300 => "01000101",27301 => "00000011",27302 => "00110010",27303 => "10110000",27304 => "10001110",27305 => "10101100",27306 => "00100001",27307 => "10011001",27308 => "00110101",27309 => "00010100",27310 => "11111111",27311 => "11110010",27312 => "01111101",27313 => "11111000",27314 => "01010111",27315 => "11010111",27316 => "10000001",27317 => "11100100",27318 => "11111101",27319 => "10011010",27320 => "11100010",27321 => "11000001",27322 => "00000101",27323 => "11111110",27324 => "11001011",27325 => "00011010",27326 => "10011011",27327 => "01000011",27328 => "10000111",27329 => "01001011",27330 => "10011010",27331 => "10110110",27332 => "00001010",27333 => "11011001",27334 => "10101110",27335 => "11110111",27336 => "01010001",27337 => "00101010",27338 => "10000000",27339 => "00111101",27340 => "10001001",27341 => "11010100",27342 => "11100101",27343 => "10101011",27344 => "11100110",27345 => "10011011",27346 => "10111001",27347 => "01001000",27348 => "00100100",27349 => "00101110",27350 => "11010000",27351 => "00010001",27352 => "01111111",27353 => "00101001",27354 => "00100011",27355 => "01001001",27356 => "11011100",27357 => "11011010",27358 => "00000010",27359 => "11110111",27360 => "10011010",27361 => "00011111",27362 => "00000111",27363 => "01100101",27364 => "10000001",27365 => "00101110",27366 => "00010110",27367 => "01001011",27368 => "01000010",27369 => "01110000",27370 => "00101100",27371 => "00100011",27372 => "10010101",27373 => "00100001",27374 => "11101001",27375 => "01101101",27376 => "10100101",27377 => "11100010",27378 => "00011101",27379 => "00010100",27380 => "10110100",27381 => "01000101",27382 => "00111101",27383 => "00001001",27384 => "01110000",27385 => "11011010",27386 => "10101111",27387 => "01000110",27388 => "00100100",27389 => "00110111",27390 => "10101011",27391 => "00110101",27392 => "11010111",27393 => "10010011",27394 => "10111000",27395 => "00011011",27396 => "00110011",27397 => "11010001",27398 => "01000011",27399 => "11001011",27400 => "11110100",27401 => "01011011",27402 => "00101000",27403 => "00110001",27404 => "10001101",27405 => "00010001",27406 => "10000101",27407 => "10101100",27408 => "00001000",27409 => "00000010",27410 => "11110000",27411 => "11001010",27412 => "11100101",27413 => "00110100",27414 => "10110100",27415 => "10101100",27416 => "11010101",27417 => "01001111",27418 => "00111010",27419 => "00100100",27420 => "00011011",27421 => "01100000",27422 => "11001010",27423 => "01110001",27424 => "01001101",27425 => "00011000",27426 => "01000111",27427 => "10111001",27428 => "00110101",27429 => "11000001",27430 => "01001110",27431 => "10110000",27432 => "00000011",27433 => "01100101",27434 => "00111100",27435 => "01111001",27436 => "01100111",27437 => "00011010",27438 => "11111011",27439 => "10000100",27440 => "01000001",27441 => "10001010",27442 => "01100111",27443 => "11110001",27444 => "11010100",27445 => "10001101",27446 => "11110011",27447 => "00100011",27448 => "00000100",27449 => "10110110",27450 => "11111011",27451 => "00000100",27452 => "00111111",27453 => "10100010",27454 => "11110011",27455 => "10100110",27456 => "10011011",27457 => "11001011",27458 => "01001100",27459 => "01000011",27460 => "11010001",27461 => "10000000",27462 => "10111001",27463 => "11110001",27464 => "10011011",27465 => "01100111",27466 => "01000011",27467 => "00100010",27468 => "11101111",27469 => "10011100",27470 => "00010101",27471 => "00011110",27472 => "11010100",27473 => "00011000",27474 => "00111001",27475 => "01110001",27476 => "11100010",27477 => "10000011",27478 => "01011001",27479 => "10111011",27480 => "00110010",27481 => "10101100",27482 => "11011001",27483 => "01111101",27484 => "01000000",27485 => "10110000",27486 => "11000111",27487 => "11100101",27488 => "10100010",27489 => "01101101",27490 => "00010111",27491 => "01000011",27492 => "11010001",27493 => "10101111",27494 => "00010101",27495 => "11101101",27496 => "10011000",27497 => "10100111",27498 => "01110111",27499 => "10011111",27500 => "01101011",27501 => "10001000",27502 => "01011110",27503 => "10110100",27504 => "01011110",27505 => "11101100",27506 => "01000010",27507 => "01001011",27508 => "00100101",27509 => "01000100",27510 => "01110001",27511 => "11111001",27512 => "11010000",27513 => "01100101",27514 => "01011100",27515 => "11100001",27516 => "01010101",27517 => "00111010",27518 => "11000100",27519 => "11010010",27520 => "10010010",27521 => "00110101",27522 => "01001110",27523 => "00111101",27524 => "01010110",27525 => "00111000",27526 => "11001100",27527 => "00110000",27528 => "10000010",27529 => "00000001",27530 => "10101100",27531 => "10100001",27532 => "10101110",27533 => "11001110",27534 => "01100111",27535 => "11100100",27536 => "00011101",27537 => "00011000",27538 => "00011000",27539 => "11010010",27540 => "00001110",27541 => "00000101",27542 => "00110110",27543 => "11001010",27544 => "01001100",27545 => "00111000",27546 => "01000100",27547 => "11110111",27548 => "11101000",27549 => "11111101",27550 => "10010000",27551 => "00110011",27552 => "10100100",27553 => "00110111",27554 => "11000000",27555 => "10111110",27556 => "11010110",27557 => "00101010",27558 => "11110101",27559 => "00100101",27560 => "00111000",27561 => "01100011",27562 => "11000110",27563 => "11000100",27564 => "10011100",27565 => "01010001",27566 => "01100011",27567 => "11110101",27568 => "00011001",27569 => "11000000",27570 => "01000010",27571 => "00101010",27572 => "11011111",27573 => "11111111",27574 => "10001101",27575 => "10110100",27576 => "01111010",27577 => "01011010",27578 => "01111011",27579 => "11010100",27580 => "11010101",27581 => "10100111",27582 => "10100110",27583 => "10001011",27584 => "10000001",27585 => "11010010",27586 => "11000111",27587 => "11001001",27588 => "10111101",27589 => "10111101",27590 => "00101010",27591 => "00101111",27592 => "00110110",27593 => "10110111",27594 => "10111010",27595 => "00101111",27596 => "01010100",27597 => "10010111",27598 => "10101010",27599 => "11000100",27600 => "01110000",27601 => "11001101",27602 => "10110011",27603 => "00010011",27604 => "00100010",27605 => "01100001",27606 => "11000001",27607 => "11010000",27608 => "11001010",27609 => "10100011",27610 => "10100001",27611 => "00010100",27612 => "00010001",27613 => "01100001",27614 => "01101011",27615 => "01011000",27616 => "11010100",27617 => "01110110",27618 => "00011110",27619 => "01111111",27620 => "10100011",27621 => "00110010",27622 => "11110011",27623 => "10010110",27624 => "01000111",27625 => "01001010",27626 => "00000100",27627 => "11101000",27628 => "01011011",27629 => "10000110",27630 => "10010110",27631 => "10110100",27632 => "01001001",27633 => "10000101",27634 => "01010100",27635 => "01010101",27636 => "01111011",27637 => "01000110",27638 => "01011000",27639 => "01100101",27640 => "00110111",27641 => "10101100",27642 => "01110100",27643 => "00011111",27644 => "11001111",27645 => "10111011",27646 => "00110000",27647 => "10111100",27648 => "10000011",27649 => "01110011",27650 => "11101100",27651 => "01100000",27652 => "01000110",27653 => "01001000",27654 => "00001100",27655 => "10111101",27656 => "00100111",27657 => "10110000",27658 => "10001010",27659 => "00101110",27660 => "01011000",27661 => "00001101",27662 => "10110111",27663 => "00111000",27664 => "01100010",27665 => "11011000",27666 => "11101000",27667 => "01100111",27668 => "01001100",27669 => "11101111",27670 => "01010100",27671 => "00100011",27672 => "01100111",27673 => "00001100",27674 => "01011011",27675 => "00001001",27676 => "10101101",27677 => "10111011",27678 => "11001110",27679 => "11010111",27680 => "11001000",27681 => "10000100",27682 => "10011000",27683 => "01000010",27684 => "10100110",27685 => "10011111",27686 => "10001010",27687 => "11101001",27688 => "10000111",27689 => "00011000",27690 => "01010101",27691 => "11111100",27692 => "11100101",27693 => "01111100",27694 => "10110111",27695 => "01101100",27696 => "11011001",27697 => "11111101",27698 => "01100010",27699 => "00001100",27700 => "10000000",27701 => "10001111",27702 => "01100110",27703 => "00000101",27704 => "00100000",27705 => "01101100",27706 => "10110111",27707 => "01101101",27708 => "11011110",27709 => "10101110",27710 => "00110001",27711 => "10111001",27712 => "00000110",27713 => "00101100",27714 => "10001001",27715 => "01011111",27716 => "01100100",27717 => "10100100",27718 => "00001101",27719 => "10010000",27720 => "00001011",27721 => "00110101",27722 => "00000100",27723 => "10100111",27724 => "11111000",27725 => "00110000",27726 => "00101001",27727 => "00100110",27728 => "11000000",27729 => "00001110",27730 => "10110011",27731 => "01101100",27732 => "00000011",27733 => "10011100",27734 => "11100010",27735 => "00111110",27736 => "10111100",27737 => "00000000",27738 => "00001101",27739 => "00100101",27740 => "11111010",27741 => "01010000",27742 => "10111111",27743 => "01011000",27744 => "01011110",27745 => "11011101",27746 => "00011101",27747 => "11001000",27748 => "11000111",27749 => "10001011",27750 => "01101110",27751 => "00110111",27752 => "01111000",27753 => "10000100",27754 => "11110110",27755 => "01110111",27756 => "01000110",27757 => "11011100",27758 => "11011010",27759 => "01100101",27760 => "11100100",27761 => "01111000",27762 => "01110010",27763 => "00011101",27764 => "11001001",27765 => "10001010",27766 => "10101000",27767 => "11100000",27768 => "01010011",27769 => "00011010",27770 => "00101001",27771 => "10100110",27772 => "10011100",27773 => "01001101",27774 => "10001110",27775 => "11010100",27776 => "11101001",27777 => "10011001",27778 => "01100111",27779 => "11110011",27780 => "01001001",27781 => "10100100",27782 => "00011011",27783 => "01011000",27784 => "00100010",27785 => "01101000",27786 => "10010110",27787 => "10100110",27788 => "11101010",27789 => "00011100",27790 => "00101101",27791 => "10001011",27792 => "10110010",27793 => "11100100",27794 => "11000110",27795 => "11001110",27796 => "11010010",27797 => "00000011",27798 => "01111000",27799 => "01001101",27800 => "10100010",27801 => "10011110",27802 => "11110011",27803 => "10100111",27804 => "10100011",27805 => "10111010",27806 => "11110100",27807 => "01010001",27808 => "10100111",27809 => "00000110",27810 => "00011011",27811 => "00110001",27812 => "10100111",27813 => "01100011",27814 => "00101111",27815 => "10001110",27816 => "01001000",27817 => "00111000",27818 => "00010111",27819 => "10010001",27820 => "11011101",27821 => "00110101",27822 => "11000110",27823 => "01000001",27824 => "11011011",27825 => "10111100",27826 => "10111101",27827 => "10100000",27828 => "00000001",27829 => "11110001",27830 => "10011010",27831 => "11101010",27832 => "00010010",27833 => "10011101",27834 => "11011101",27835 => "10011101",27836 => "11101100",27837 => "01000010",27838 => "10100001",27839 => "01011110",27840 => "00101010",27841 => "10000010",27842 => "10101111",27843 => "01111111",27844 => "10110001",27845 => "01101001",27846 => "11010101",27847 => "01101100",27848 => "11001010",27849 => "10010100",27850 => "11100001",27851 => "11110001",27852 => "10100101",27853 => "11010001",27854 => "00100010",27855 => "01011000",27856 => "11111010",27857 => "10101010",27858 => "01100000",27859 => "00000001",27860 => "00101001",27861 => "10001101",27862 => "10011100",27863 => "10110110",27864 => "01100100",27865 => "01100101",27866 => "11111001",27867 => "11100110",27868 => "00100101",27869 => "01101100",27870 => "10001100",27871 => "01101001",27872 => "00010011",27873 => "10100011",27874 => "01100011",27875 => "01110001",27876 => "10101101",27877 => "11111000",27878 => "00111100",27879 => "10000100",27880 => "11100101",27881 => "10010101",27882 => "11111000",27883 => "00110001",27884 => "10111011",27885 => "10111011",27886 => "11111001",27887 => "10000100",27888 => "11011110",27889 => "11100000",27890 => "11111011",27891 => "00011110",27892 => "10110011",27893 => "10111110",27894 => "01101000",27895 => "11000110",27896 => "01101100",27897 => "11110001",27898 => "11000110",27899 => "10100111",27900 => "00101101",27901 => "11001100",27902 => "01010101",27903 => "01000110",27904 => "11111001",27905 => "00111111",27906 => "11101100",27907 => "11101000",27908 => "01011101",27909 => "11011011",27910 => "00110101",27911 => "11001110",27912 => "10100110",27913 => "11011110",27914 => "00010000",27915 => "10100111",27916 => "01011001",27917 => "00100111",27918 => "10110111",27919 => "01101011",27920 => "10011110",27921 => "01101101",27922 => "01111100",27923 => "01110111",27924 => "00111101",27925 => "10011110",27926 => "01101100",27927 => "10111011",27928 => "00111000",27929 => "01010001",27930 => "01100110",27931 => "10000000",27932 => "11000111",27933 => "00000100",27934 => "10101110",27935 => "00101101",27936 => "01000010",27937 => "01011110",27938 => "01101010",27939 => "11000011",27940 => "11010111",27941 => "01111001",27942 => "00110111",27943 => "10110110",27944 => "01010011",27945 => "11100000",27946 => "01101000",27947 => "00111100",27948 => "00100001",27949 => "00111001",27950 => "11101011",27951 => "00111011",27952 => "00011111",27953 => "11100011",27954 => "00101101",27955 => "01110111",27956 => "01011100",27957 => "01100010",27958 => "11000111",27959 => "11111101",27960 => "00011110",27961 => "01001011",27962 => "11110100",27963 => "01011111",27964 => "11101100",27965 => "10110111",27966 => "10011001",27967 => "01111110",27968 => "10000000",27969 => "01111110",27970 => "11100000",27971 => "00100100",27972 => "11100001",27973 => "01001100",27974 => "10000001",27975 => "10001011",27976 => "11011001",27977 => "11111110",27978 => "10110001",27979 => "01010000",27980 => "11010100",27981 => "10110000",27982 => "10010011",27983 => "11111000",27984 => "10010101",27985 => "00011000",27986 => "11011010",27987 => "11010011",27988 => "01011100",27989 => "01101010",27990 => "10010101",27991 => "01010000",27992 => "00110101",27993 => "01011010",27994 => "10011010",27995 => "10010110",27996 => "11111000",27997 => "10010101",27998 => "01101011",27999 => "00000111",28000 => "11000011",28001 => "10101101",28002 => "10010011",28003 => "10110000",28004 => "00110101",28005 => "11001010",28006 => "10000100",28007 => "11101111",28008 => "00100010",28009 => "01000101",28010 => "10011001",28011 => "11101101",28012 => "11101000",28013 => "11010110",28014 => "11000010",28015 => "00110000",28016 => "01100100",28017 => "00011111",28018 => "01011100",28019 => "01100110",28020 => "00101100",28021 => "00001101",28022 => "11110110",28023 => "11100010",28024 => "01111011",28025 => "00110111",28026 => "11100011",28027 => "11000011",28028 => "00111110",28029 => "00100110",28030 => "11000101",28031 => "11101000",28032 => "00011111",28033 => "00011100",28034 => "01001000",28035 => "11101001",28036 => "11001011",28037 => "11011100",28038 => "11010001",28039 => "01001001",28040 => "10100001",28041 => "11010111",28042 => "10110101",28043 => "10011011",28044 => "00000011",28045 => "11011001",28046 => "00010100",28047 => "00110101",28048 => "01010101",28049 => "11110101",28050 => "10110001",28051 => "11000001",28052 => "01100011",28053 => "01010010",28054 => "01011010",28055 => "10000110",28056 => "01001010",28057 => "10011000",28058 => "00110111",28059 => "00010010",28060 => "01000010",28061 => "01010001",28062 => "00001010",28063 => "00010001",28064 => "11011111",28065 => "10000001",28066 => "01101101",28067 => "10110000",28068 => "00001111",28069 => "10001010",28070 => "10011100",28071 => "00010001",28072 => "10101010",28073 => "01110100",28074 => "01001001",28075 => "11111111",28076 => "00111010",28077 => "01100101",28078 => "00101101",28079 => "00000100",28080 => "00000100",28081 => "01110001",28082 => "01100000",28083 => "01001100",28084 => "01001010",28085 => "00000011",28086 => "00011100",28087 => "11001110",28088 => "11011010",28089 => "11111011",28090 => "11101100",28091 => "00111111",28092 => "00001111",28093 => "01110111",28094 => "01110110",28095 => "11010111",28096 => "00010111",28097 => "00001100",28098 => "00010000",28099 => "01011001",28100 => "00111101",28101 => "01000000",28102 => "00100010",28103 => "01101000",28104 => "01100000",28105 => "01100001",28106 => "10100100",28107 => "10101100",28108 => "11110101",28109 => "01011010",28110 => "10000111",28111 => "11101100",28112 => "01001001",28113 => "10000110",28114 => "01011010",28115 => "11110010",28116 => "10101011",28117 => "01010101",28118 => "11111001",28119 => "01011110",28120 => "00111101",28121 => "11000010",28122 => "11100001",28123 => "11010100",28124 => "10100000",28125 => "01011110",28126 => "10001010",28127 => "00110101",28128 => "01101110",28129 => "11111011",28130 => "11100000",28131 => "01101110",28132 => "11011010",28133 => "11000110",28134 => "11010011",28135 => "01111111",28136 => "00001101",28137 => "01111000",28138 => "00011111",28139 => "00110111",28140 => "01010000",28141 => "00010111",28142 => "01100101",28143 => "00111010",28144 => "11011011",28145 => "11011110",28146 => "10100100",28147 => "11011011",28148 => "11001001",28149 => "01000110",28150 => "11101000",28151 => "00100101",28152 => "00001001",28153 => "10101101",28154 => "10010010",28155 => "11100110",28156 => "00000111",28157 => "11111010",28158 => "11010001",28159 => "00001010",28160 => "10110100",28161 => "10010001",28162 => "00100111",28163 => "11010101",28164 => "00111010",28165 => "11100110",28166 => "10101000",28167 => "10010001",28168 => "11100000",28169 => "10101001",28170 => "01111111",28171 => "11100111",28172 => "10100011",28173 => "11001000",28174 => "00011000",28175 => "00010001",28176 => "00110111",28177 => "10101000",28178 => "11100010",28179 => "01000010",28180 => "00011010",28181 => "11001000",28182 => "11000010",28183 => "11101001",28184 => "11110100",28185 => "00111010",28186 => "10001000",28187 => "01011110",28188 => "01111010",28189 => "11101110",28190 => "00111110",28191 => "01110001",28192 => "01100110",28193 => "00100101",28194 => "01111011",28195 => "00010100",28196 => "01000110",28197 => "10111011",28198 => "00000010",28199 => "11001000",28200 => "10100000",28201 => "00010110",28202 => "00100001",28203 => "00100101",28204 => "01001010",28205 => "00000010",28206 => "01011000",28207 => "10010100",28208 => "11000111",28209 => "01000010",28210 => "10100111",28211 => "10011100",28212 => "00010001",28213 => "00100000",28214 => "11110000",28215 => "10010101",28216 => "01100010",28217 => "00101100",28218 => "01111011",28219 => "11000111",28220 => "10111111",28221 => "01101110",28222 => "11111011",28223 => "00111110",28224 => "01010100",28225 => "11010001",28226 => "01000001",28227 => "00010110",28228 => "10011010",28229 => "11100101",28230 => "11110110",28231 => "00110001",28232 => "10011100",28233 => "01001100",28234 => "10010111",28235 => "01001110",28236 => "00101111",28237 => "11001110",28238 => "10011111",28239 => "10100000",28240 => "01010101",28241 => "00111001",28242 => "00011111",28243 => "11011000",28244 => "00010000",28245 => "01001110",28246 => "10110000",28247 => "00001101",28248 => "00100111",28249 => "01110011",28250 => "00011001",28251 => "10000001",28252 => "11000110",28253 => "00011010",28254 => "11011101",28255 => "01010011",28256 => "01010011",28257 => "11101111",28258 => "00010110",28259 => "00000111",28260 => "00000001",28261 => "11100110",28262 => "10110010",28263 => "11001010",28264 => "00000100",28265 => "00101010",28266 => "11010001",28267 => "11000001",28268 => "11101100",28269 => "11010101",28270 => "10110111",28271 => "00010001",28272 => "10000011",28273 => "00101011",28274 => "00110110",28275 => "00010100",28276 => "11011011",28277 => "11011001",28278 => "10000100",28279 => "10100000",28280 => "00000001",28281 => "01111101",28282 => "00011010",28283 => "01011001",28284 => "10111000",28285 => "10000110",28286 => "10100110",28287 => "10011001",28288 => "11000011",28289 => "11011011",28290 => "00011010",28291 => "10010000",28292 => "01101101",28293 => "00011010",28294 => "00010101",28295 => "11101001",28296 => "11000001",28297 => "11110110",28298 => "01001011",28299 => "11010000",28300 => "11101101",28301 => "11001101",28302 => "01100000",28303 => "10000101",28304 => "10001011",28305 => "01101100",28306 => "11000001",28307 => "00000110",28308 => "10010000",28309 => "10100100",28310 => "00001111",28311 => "01100000",28312 => "10110001",28313 => "10111011",28314 => "00111001",28315 => "01110111",28316 => "01111000",28317 => "00001100",28318 => "10100011",28319 => "11000111",28320 => "11010011",28321 => "10110100",28322 => "10111110",28323 => "01000111",28324 => "11111100",28325 => "01100111",28326 => "01010111",28327 => "00001100",28328 => "11111000",28329 => "10100100",28330 => "01111010",28331 => "01100000",28332 => "11000001",28333 => "00010000",28334 => "10100001",28335 => "10001001",28336 => "11011100",28337 => "01101001",28338 => "11110000",28339 => "11010000",28340 => "10011001",28341 => "11111100",28342 => "10001100",28343 => "11001000",28344 => "11100111",28345 => "11100111",28346 => "10111101",28347 => "10100001",28348 => "10100011",28349 => "11101100",28350 => "11001011",28351 => "01111010",28352 => "11100011",28353 => "01001000",28354 => "11001001",28355 => "00111011",28356 => "10111101",28357 => "10010010",28358 => "11111011",28359 => "10110001",28360 => "01100100",28361 => "10100001",28362 => "01110000",28363 => "01011100",28364 => "11011010",28365 => "00001011",28366 => "10010001",28367 => "01011010",28368 => "11100100",28369 => "11100000",28370 => "11110000",28371 => "01111100",28372 => "11111011",28373 => "11100010",28374 => "00110100",28375 => "00111101",28376 => "01000011",28377 => "10001000",28378 => "10101011",28379 => "01111001",28380 => "10001011",28381 => "10011100",28382 => "00010110",28383 => "11110001",28384 => "01110011",28385 => "01010000",28386 => "00110111",28387 => "01010110",28388 => "01101010",28389 => "00101001",28390 => "11100101",28391 => "10101000",28392 => "01010101",28393 => "11100101",28394 => "10111000",28395 => "11000000",28396 => "01101100",28397 => "10110101",28398 => "10110000",28399 => "11110011",28400 => "10011010",28401 => "10011100",28402 => "11111101",28403 => "10000100",28404 => "01101100",28405 => "01011101",28406 => "01001010",28407 => "01000101",28408 => "01101111",28409 => "00101111",28410 => "00101111",28411 => "10011010",28412 => "00001001",28413 => "10100001",28414 => "00101100",28415 => "10010100",28416 => "01001001",28417 => "11011101",28418 => "10101111",28419 => "00101010",28420 => "10111011",28421 => "11110000",28422 => "10011110",28423 => "10110101",28424 => "00111100",28425 => "10100110",28426 => "10011111",28427 => "01011111",28428 => "01011001",28429 => "01000010",28430 => "01011110",28431 => "00110110",28432 => "01000010",28433 => "10000010",28434 => "11110101",28435 => "00111111",28436 => "11000110",28437 => "00101111",28438 => "10001011",28439 => "00011100",28440 => "01100010",28441 => "11101101",28442 => "00000110",28443 => "01010110",28444 => "00001000",28445 => "00011111",28446 => "10011110",28447 => "10011110",28448 => "11110111",28449 => "11000101",28450 => "01001011",28451 => "00000111",28452 => "11111100",28453 => "10111011",28454 => "00010111",28455 => "01110110",28456 => "00100111",28457 => "10010111",28458 => "11110101",28459 => "00010110",28460 => "10011111",28461 => "11010100",28462 => "01110001",28463 => "01100100",28464 => "00010110",28465 => "11111101",28466 => "01001001",28467 => "01010100",28468 => "11010010",28469 => "10100010",28470 => "00110100",28471 => "10000001",28472 => "00010000",28473 => "10010100",28474 => "10101101",28475 => "00011100",28476 => "00110010",28477 => "11000001",28478 => "10110000",28479 => "01000001",28480 => "00101111",28481 => "00001111",28482 => "01101010",28483 => "11000001",28484 => "01011000",28485 => "10011000",28486 => "10011100",28487 => "10100000",28488 => "00000011",28489 => "11001111",28490 => "01101000",28491 => "00110000",28492 => "01010110",28493 => "01000010",28494 => "01001110",28495 => "11111001",28496 => "10100100",28497 => "00101000",28498 => "10001010",28499 => "10101010",28500 => "10111111",28501 => "11011011",28502 => "01000011",28503 => "00110101",28504 => "10111100",28505 => "10001111",28506 => "11000100",28507 => "01010011",28508 => "01000001",28509 => "00001101",28510 => "10111010",28511 => "11001001",28512 => "10000100",28513 => "10010000",28514 => "10101110",28515 => "11011111",28516 => "11001011",28517 => "11111000",28518 => "00111000",28519 => "00101000",28520 => "00100111",28521 => "00011101",28522 => "01111000",28523 => "11001111",28524 => "10001100",28525 => "10001100",28526 => "11110101",28527 => "11011011",28528 => "10010001",28529 => "00011001",28530 => "11001110",28531 => "11111011",28532 => "00110111",28533 => "01000101",28534 => "01001000",28535 => "01101110",28536 => "10011011",28537 => "11100001",28538 => "00010100",28539 => "01100101",28540 => "00100111",28541 => "11110011",28542 => "00111001",28543 => "00100011",28544 => "11010011",28545 => "00000000",28546 => "10011101",28547 => "01010011",28548 => "01010110",28549 => "11110101",28550 => "00110011",28551 => "10000000",28552 => "01111011",28553 => "11111110",28554 => "00101011",28555 => "11111110",28556 => "01001010",28557 => "01001000",28558 => "10001110",28559 => "00111100",28560 => "10000111",28561 => "11000100",28562 => "00010011",28563 => "10010100",28564 => "01101101",28565 => "11111100",28566 => "11101011",28567 => "00000001",28568 => "01110000",28569 => "10011010",28570 => "10011101",28571 => "01011000",28572 => "11000111",28573 => "00100101",28574 => "10101111",28575 => "01101000",28576 => "01011100",28577 => "00010000",28578 => "10000100",28579 => "00011011",28580 => "10001000",28581 => "01010101",28582 => "10001000",28583 => "00010111",28584 => "10101111",28585 => "11001101",28586 => "01000111",28587 => "01000110",28588 => "10011010",28589 => "11111000",28590 => "11100101",28591 => "00000001",28592 => "11001010",28593 => "00001111",28594 => "11100110",28595 => "01011010",28596 => "00000001",28597 => "11111001",28598 => "10110011",28599 => "10110010",28600 => "01111010",28601 => "11111010",28602 => "10101000",28603 => "01000000",28604 => "01010100",28605 => "00101001",28606 => "11111011",28607 => "11001111",28608 => "00011010",28609 => "01011100",28610 => "00011111",28611 => "00100111",28612 => "01011110",28613 => "01101111",28614 => "00100101",28615 => "00000100",28616 => "11101010",28617 => "11011010",28618 => "01001000",28619 => "11010111",28620 => "10001110",28621 => "10001110",28622 => "10010100",28623 => "01111110",28624 => "00110101",28625 => "01000011",28626 => "01110010",28627 => "10100001",28628 => "11110000",28629 => "10001100",28630 => "11111110",28631 => "10010101",28632 => "00010101",28633 => "10010000",28634 => "01100000",28635 => "00110111",28636 => "10010011",28637 => "11010001",28638 => "10010101",28639 => "01110011",28640 => "00011001",28641 => "01110011",28642 => "11001001",28643 => "10001110",28644 => "10111101",28645 => "11101001",28646 => "01100100",28647 => "10011111",28648 => "00011001",28649 => "11100100",28650 => "11000011",28651 => "01010110",28652 => "01001100",28653 => "00010001",28654 => "11100001",28655 => "00011010",28656 => "10000111",28657 => "00110101",28658 => "01010011",28659 => "00000000",28660 => "11110110",28661 => "00110010",28662 => "01101010",28663 => "11111110",28664 => "11011100",28665 => "01111000",28666 => "10111011",28667 => "01101100",28668 => "01000111",28669 => "00010010",28670 => "01000000",28671 => "11001011",28672 => "11110111",28673 => "01110111",28674 => "00110100",28675 => "01111111",28676 => "10010011",28677 => "00110100",28678 => "01110100",28679 => "00101111",28680 => "11100010",28681 => "00001001",28682 => "00010000",28683 => "11101010",28684 => "00010011",28685 => "00101101",28686 => "00000110",28687 => "10011000",28688 => "11011001",28689 => "10010001",28690 => "00110110",28691 => "11110111",28692 => "01101101",28693 => "01000001",28694 => "00000000",28695 => "00110001",28696 => "10010000",28697 => "00111111",28698 => "01001110",28699 => "01001000",28700 => "01001001",28701 => "01101111",28702 => "00011001",28703 => "00011001",28704 => "10011011",28705 => "11001100",28706 => "10010010",28707 => "10010101",28708 => "10001111",28709 => "11011000",28710 => "10010101",28711 => "00100100",28712 => "01001110",28713 => "10111001",28714 => "10100010",28715 => "10010101",28716 => "01001100",28717 => "10100101",28718 => "10100000",28719 => "00010010",28720 => "11001000",28721 => "01100111",28722 => "10100101",28723 => "01000110",28724 => "01010110",28725 => "00110111",28726 => "01101110",28727 => "11110010",28728 => "10000111",28729 => "11010100",28730 => "10100100",28731 => "11010001",28732 => "10111011",28733 => "10110101",28734 => "01100010",28735 => "11111000",28736 => "01000101",28737 => "10010101",28738 => "01111110",28739 => "00100000",28740 => "11010110",28741 => "01010000",28742 => "00100011",28743 => "00100100",28744 => "01100100",28745 => "11111011",28746 => "00000100",28747 => "11000001",28748 => "01010001",28749 => "11011011",28750 => "00001100",28751 => "00101111",28752 => "11001100",28753 => "01011100",28754 => "11100100",28755 => "00110100",28756 => "01100010",28757 => "01000010",28758 => "10000000",28759 => "10010010",28760 => "01000110",28761 => "00111001",28762 => "00001111",28763 => "01000111",28764 => "00111010",28765 => "00010110",28766 => "10101100",28767 => "11000100",28768 => "01110010",28769 => "11010000",28770 => "11010101",28771 => "10111011",28772 => "01000000",28773 => "01001101",28774 => "00000110",28775 => "10010011",28776 => "11011001",28777 => "01000000",28778 => "11100000",28779 => "11100000",28780 => "11111100",28781 => "01101101",28782 => "11101101",28783 => "01111101",28784 => "01110000",28785 => "10000001",28786 => "00110111",28787 => "00011110",28788 => "10001111",28789 => "01111011",28790 => "11111001",28791 => "01011111",28792 => "01010011",28793 => "00111010",28794 => "11001010",28795 => "11110011",28796 => "01111111",28797 => "11010001",28798 => "01010010",28799 => "01000101",28800 => "01111010",28801 => "01101110",28802 => "11110101",28803 => "10000000",28804 => "01101110",28805 => "00000001",28806 => "11101010",28807 => "01001101",28808 => "11011101",28809 => "01100100",28810 => "00001110",28811 => "00011001",28812 => "01000101",28813 => "00001111",28814 => "01101100",28815 => "01000100",28816 => "11000011",28817 => "11100001",28818 => "10010000",28819 => "11010111",28820 => "11011010",28821 => "11101110",28822 => "01110001",28823 => "00000010",28824 => "11011001",28825 => "01011000",28826 => "00111010",28827 => "11011000",28828 => "00000010",28829 => "10100001",28830 => "10001001",28831 => "10111001",28832 => "00011001",28833 => "00101011",28834 => "00011111",28835 => "00010001",28836 => "11110111",28837 => "10101101",28838 => "11000111",28839 => "11000110",28840 => "10011000",28841 => "00011100",28842 => "11110101",28843 => "00000101",28844 => "11011001",28845 => "11110001",28846 => "01100010",28847 => "10111010",28848 => "10111001",28849 => "01100010",28850 => "10000001",28851 => "10100110",28852 => "10011001",28853 => "01001011",28854 => "11111100",28855 => "11100010",28856 => "10110001",28857 => "01110111",28858 => "00101000",28859 => "01111111",28860 => "01110000",28861 => "11000111",28862 => "00000000",28863 => "00110100",28864 => "11110000",28865 => "01000011",28866 => "01110101",28867 => "00110010",28868 => "00000101",28869 => "11101100",28870 => "10100100",28871 => "11001110",28872 => "10110010",28873 => "00010100",28874 => "01100110",28875 => "00010101",28876 => "11000110",28877 => "10001010",28878 => "01010111",28879 => "11101111",28880 => "11000010",28881 => "11000100",28882 => "01111001",28883 => "00111110",28884 => "10011111",28885 => "11000100",28886 => "10110001",28887 => "10010101",28888 => "10010000",28889 => "01111110",28890 => "00001010",28891 => "01100111",28892 => "00011011",28893 => "10100011",28894 => "11000010",28895 => "01111111",28896 => "10111010",28897 => "10111100",28898 => "11110101",28899 => "00001000",28900 => "11000110",28901 => "01000000",28902 => "00000100",28903 => "00110111",28904 => "00110000",28905 => "11000000",28906 => "10111010",28907 => "10000001",28908 => "00011000",28909 => "11111101",28910 => "01011111",28911 => "11110011",28912 => "01000110",28913 => "01011010",28914 => "01111100",28915 => "01111010",28916 => "01101101",28917 => "00001110",28918 => "10011101",28919 => "11101100",28920 => "10100000",28921 => "11000110",28922 => "11010011",28923 => "11011111",28924 => "10001101",28925 => "00100101",28926 => "10011100",28927 => "11101000",28928 => "01010010",28929 => "10001110",28930 => "01001110",28931 => "01011110",28932 => "11000111",28933 => "01000110",28934 => "01100111",28935 => "00001010",28936 => "01101110",28937 => "00001010",28938 => "01010011",28939 => "11010111",28940 => "10111010",28941 => "10000001",28942 => "01000110",28943 => "00111011",28944 => "10001111",28945 => "01111101",28946 => "10101001",28947 => "10101001",28948 => "11010111",28949 => "11110000",28950 => "10011101",28951 => "00111011",28952 => "11000100",28953 => "01110100",28954 => "10101011",28955 => "11010000",28956 => "00011111",28957 => "11010101",28958 => "00010010",28959 => "00000101",28960 => "11001001",28961 => "11010110",28962 => "10100111",28963 => "10010100",28964 => "01111011",28965 => "01100010",28966 => "10000101",28967 => "01001010",28968 => "00011101",28969 => "01111010",28970 => "00001110",28971 => "11100010",28972 => "10010110",28973 => "11000000",28974 => "00101011",28975 => "11000010",28976 => "10010110",28977 => "11010101",28978 => "11110000",28979 => "01110010",28980 => "01001110",28981 => "10111011",28982 => "00000010",28983 => "01100100",28984 => "00010110",28985 => "01010011",28986 => "10000101",28987 => "10101110",28988 => "01010001",28989 => "01110101",28990 => "11010000",28991 => "00010111",28992 => "01110000",28993 => "10100101",28994 => "01110101",28995 => "00000100",28996 => "00110011",28997 => "11011010",28998 => "01110010",28999 => "00001100",29000 => "01000000",29001 => "00001011",29002 => "10110100",29003 => "01111111",29004 => "01101101",29005 => "11000001",29006 => "01100100",29007 => "10000011",29008 => "01100011",29009 => "10001000",29010 => "10010111",29011 => "11011111",29012 => "10100000",29013 => "10101011",29014 => "00100001",29015 => "11011101",29016 => "01000101",29017 => "00011111",29018 => "10011110",29019 => "10000111",29020 => "00111000",29021 => "01010001",29022 => "11100101",29023 => "10110001",29024 => "10001010",29025 => "00001001",29026 => "10110010",29027 => "01110111",29028 => "00110101",29029 => "00101000",29030 => "11011011",29031 => "11111111",29032 => "11111101",29033 => "11110101",29034 => "10101011",29035 => "01100111",29036 => "01001000",29037 => "10111011",29038 => "01110100",29039 => "01010111",29040 => "11001001",29041 => "11010101",29042 => "00011000",29043 => "11000111",29044 => "10111001",29045 => "00001100",29046 => "01110000",29047 => "01110101",29048 => "11111010",29049 => "00100110",29050 => "01010111",29051 => "00010100",29052 => "01000010",29053 => "10010001",29054 => "00110111",29055 => "01011100",29056 => "00011100",29057 => "11001111",29058 => "11101100",29059 => "01110111",29060 => "00101010",29061 => "10110010",29062 => "11011110",29063 => "10001100",29064 => "00100000",29065 => "11110101",29066 => "10110111",29067 => "11011110",29068 => "10010111",29069 => "01010011",29070 => "11110001",29071 => "10000011",29072 => "01110000",29073 => "00000100",29074 => "11001110",29075 => "00011110",29076 => "00011101",29077 => "00000111",29078 => "11000000",29079 => "10010000",29080 => "00011100",29081 => "10111001",29082 => "10100010",29083 => "00001010",29084 => "01100011",29085 => "11100100",29086 => "01011100",29087 => "11001001",29088 => "01011000",29089 => "01101101",29090 => "11000000",29091 => "11010001",29092 => "11101001",29093 => "01100101",29094 => "00110001",29095 => "10110000",29096 => "11111110",29097 => "10100111",29098 => "00011000",29099 => "01111011",29100 => "01011100",29101 => "01100101",29102 => "01010100",29103 => "00011100",29104 => "10111110",29105 => "01111000",29106 => "01000010",29107 => "00101110",29108 => "10010110",29109 => "11010111",29110 => "01100011",29111 => "01011100",29112 => "10011110",29113 => "10111100",29114 => "01010110",29115 => "01001001",29116 => "01110111",29117 => "01001110",29118 => "00000011",29119 => "00001101",29120 => "11000000",29121 => "11111111",29122 => "01011010",29123 => "01011110",29124 => "00101001",29125 => "10000101",29126 => "00100111",29127 => "00010110",29128 => "01111110",29129 => "10100110",29130 => "00110011",29131 => "11100101",29132 => "00110010",29133 => "11100000",29134 => "11001111",29135 => "00001000",29136 => "10110111",29137 => "10100010",29138 => "10110011",29139 => "01000000",29140 => "00111011",29141 => "10100001",29142 => "01110110",29143 => "10000100",29144 => "00001101",29145 => "01110011",29146 => "11101001",29147 => "10000111",29148 => "00110111",29149 => "10110101",29150 => "10111000",29151 => "00111111",29152 => "00000011",29153 => "01110100",29154 => "01001010",29155 => "01100011",29156 => "11001110",29157 => "00101000",29158 => "10100000",29159 => "00111100",29160 => "11110000",29161 => "00100100",29162 => "00000001",29163 => "11001110",29164 => "11101001",29165 => "01100011",29166 => "10001101",29167 => "01100100",29168 => "10011000",29169 => "11001101",29170 => "00010011",29171 => "01111101",29172 => "11001000",29173 => "00110101",29174 => "11110000",29175 => "00111000",29176 => "01111010",29177 => "11000011",29178 => "00101011",29179 => "01011010",29180 => "00010100",29181 => "10000000",29182 => "00111000",29183 => "11100011",29184 => "00001110",29185 => "00000010",29186 => "10010110",29187 => "00011101",29188 => "01000110",29189 => "10000110",29190 => "00111000",29191 => "00001100",29192 => "00011111",29193 => "10010001",29194 => "01001001",29195 => "10001110",29196 => "01111111",29197 => "01110001",29198 => "00100100",29199 => "10111100",29200 => "11110110",29201 => "00101110",29202 => "10100111",29203 => "01101000",29204 => "00110101",29205 => "00111010",29206 => "11011001",29207 => "11010000",29208 => "00100110",29209 => "01010010",29210 => "11011011",29211 => "11110100",29212 => "10010001",29213 => "01000001",29214 => "11011011",29215 => "10000101",29216 => "00001011",29217 => "01111001",29218 => "01110000",29219 => "01010111",29220 => "01011001",29221 => "11111101",29222 => "00011101",29223 => "00101001",29224 => "11010011",29225 => "10101001",29226 => "11100111",29227 => "01011100",29228 => "10100010",29229 => "00010001",29230 => "11001011",29231 => "01101101",29232 => "10111010",29233 => "01111100",29234 => "10101111",29235 => "10011011",29236 => "10011111",29237 => "11110101",29238 => "11001100",29239 => "11101100",29240 => "01001010",29241 => "01110110",29242 => "00110111",29243 => "01101001",29244 => "00010100",29245 => "00100100",29246 => "00011101",29247 => "00001111",29248 => "01110101",29249 => "01000001",29250 => "11101110",29251 => "00010101",29252 => "10011011",29253 => "01000110",29254 => "00100001",29255 => "11110011",29256 => "11110111",29257 => "00100001",29258 => "01000010",29259 => "10001101",29260 => "00100110",29261 => "00101010",29262 => "01011010",29263 => "10100110",29264 => "00000011",29265 => "00110111",29266 => "00000101",29267 => "11111111",29268 => "11010010",29269 => "10110110",29270 => "10001111",29271 => "11000111",29272 => "01010010",29273 => "11001100",29274 => "00110101",29275 => "11100011",29276 => "01011010",29277 => "11000100",29278 => "10101011",29279 => "00110111",29280 => "01111000",29281 => "01100011",29282 => "01101110",29283 => "10100010",29284 => "01001110",29285 => "01111100",29286 => "10110010",29287 => "11000011",29288 => "01101000",29289 => "01001100",29290 => "00010101",29291 => "01010001",29292 => "00011110",29293 => "10001001",29294 => "00000101",29295 => "10010011",29296 => "01101110",29297 => "10011000",29298 => "00100000",29299 => "01001111",29300 => "11101100",29301 => "10111100",29302 => "10110111",29303 => "11100000",29304 => "01111111",29305 => "11010101",29306 => "01100110",29307 => "01011001",29308 => "01110111",29309 => "01101011",29310 => "01110010",29311 => "10001100",29312 => "01001100",29313 => "00110100",29314 => "00101010",29315 => "10011000",29316 => "10101010",29317 => "10111110",29318 => "11001110",29319 => "01110011",29320 => "00101000",29321 => "11010000",29322 => "10100001",29323 => "00000110",29324 => "01010111",29325 => "00001011",29326 => "01001011",29327 => "11011011",29328 => "00110010",29329 => "10110001",29330 => "10000101",29331 => "01100101",29332 => "10111110",29333 => "00101000",29334 => "01100101",29335 => "01011110",29336 => "01010101",29337 => "01100010",29338 => "11111011",29339 => "00011101",29340 => "00110100",29341 => "00100000",29342 => "00001010",29343 => "01110001",29344 => "00001000",29345 => "10100000",29346 => "00110011",29347 => "00000000",29348 => "11000011",29349 => "11010011",29350 => "01000000",29351 => "11001110",29352 => "10100100",29353 => "00001000",29354 => "01101011",29355 => "10100001",29356 => "01100101",29357 => "00001100",29358 => "01110011",29359 => "11010100",29360 => "01101101",29361 => "01010110",29362 => "00101110",29363 => "10110010",29364 => "00011101",29365 => "01100100",29366 => "00001100",29367 => "01011110",29368 => "00111011",29369 => "11011111",29370 => "01101011",29371 => "01100101",29372 => "01100010",29373 => "01000110",29374 => "01011011",29375 => "01011101",29376 => "01010001",29377 => "10111010",29378 => "10100010",29379 => "11101010",29380 => "11001111",29381 => "01111110",29382 => "01010001",29383 => "10010000",29384 => "01101000",29385 => "10000001",29386 => "00011010",29387 => "10100111",29388 => "00100010",29389 => "10101111",29390 => "00011101",29391 => "10111010",29392 => "10101001",29393 => "11011000",29394 => "01100101",29395 => "10110110",29396 => "10111000",29397 => "00111111",29398 => "11010000",29399 => "00000111",29400 => "11000111",29401 => "00010010",29402 => "01111000",29403 => "00101110",29404 => "01111111",29405 => "00001010",29406 => "01010101",29407 => "10111101",29408 => "11110110",29409 => "01010001",29410 => "00100110",29411 => "10111101",29412 => "11111101",29413 => "01011111",29414 => "01001101",29415 => "00111100",29416 => "01000000",29417 => "01000001",29418 => "01010101",29419 => "01000111",29420 => "10101000",29421 => "00110110",29422 => "01000110",29423 => "11111111",29424 => "01010111",29425 => "11110010",29426 => "10111100",29427 => "10000010",29428 => "00111011",29429 => "10100101",29430 => "10101001",29431 => "00100011",29432 => "01101111",29433 => "10010010",29434 => "11001010",29435 => "10101000",29436 => "01011011",29437 => "00010111",29438 => "10110101",29439 => "11101101",29440 => "10111110",29441 => "01111000",29442 => "00100111",29443 => "01001011",29444 => "11001101",29445 => "00100001",29446 => "00100101",29447 => "11111100",29448 => "10010101",29449 => "11011010",29450 => "10010011",29451 => "00110001",29452 => "00010011",29453 => "10001010",29454 => "01010111",29455 => "10101011",29456 => "00101111",29457 => "11000101",29458 => "11110000",29459 => "00101100",29460 => "10011111",29461 => "10011001",29462 => "10001010",29463 => "11010111",29464 => "00111001",29465 => "11011001",29466 => "10101111",29467 => "00011100",29468 => "10110101",29469 => "00111000",29470 => "00110001",29471 => "10000000",29472 => "10000110",29473 => "01111011",29474 => "11110010",29475 => "11011100",29476 => "10110111",29477 => "01101001",29478 => "01101000",29479 => "01110100",29480 => "10000101",29481 => "11111010",29482 => "00100111",29483 => "11101010",29484 => "11111011",29485 => "11011101",29486 => "01110001",29487 => "10011101",29488 => "00001110",29489 => "10010100",29490 => "00001110",29491 => "00100101",29492 => "11111000",29493 => "11110100",29494 => "01110000",29495 => "11010000",29496 => "00010001",29497 => "00001111",29498 => "00011110",29499 => "10011110",29500 => "11000010",29501 => "11110111",29502 => "11111011",29503 => "11010100",29504 => "01011001",29505 => "00101111",29506 => "00100011",29507 => "01110100",29508 => "10010010",29509 => "10001111",29510 => "01010110",29511 => "01010011",29512 => "11000110",29513 => "10001001",29514 => "01101111",29515 => "01111100",29516 => "00111011",29517 => "01001001",29518 => "10010101",29519 => "10110010",29520 => "01110011",29521 => "10000111",29522 => "11110001",29523 => "11110010",29524 => "10010001",29525 => "10111000",29526 => "11101100",29527 => "01110101",29528 => "10110111",29529 => "01000110",29530 => "10001000",29531 => "00111010",29532 => "01101101",29533 => "00010001",29534 => "11000111",29535 => "01101110",29536 => "10011100",29537 => "10000010",29538 => "10111000",29539 => "01011000",29540 => "10101001",29541 => "00001001",29542 => "00111110",29543 => "11110010",29544 => "00001101",29545 => "00110000",29546 => "00000111",29547 => "00010111",29548 => "00100110",29549 => "00010101",29550 => "10011101",29551 => "01110100",29552 => "01010010",29553 => "10000110",29554 => "10101110",29555 => "10101011",29556 => "11100110",29557 => "10001110",29558 => "01011010",29559 => "10011000",29560 => "10111110",29561 => "00110011",29562 => "00001111",29563 => "01100100",29564 => "10100000",29565 => "11010001",29566 => "00001011",29567 => "00100001",29568 => "10010111",29569 => "00100011",29570 => "00001111",29571 => "11011010",29572 => "11100011",29573 => "00111100",29574 => "01011101",29575 => "00100111",29576 => "10010011",29577 => "01101001",29578 => "00101110",29579 => "00011000",29580 => "00011000",29581 => "00001001",29582 => "11100010",29583 => "11111011",29584 => "01011101",29585 => "00000000",29586 => "00011010",29587 => "01111111",29588 => "10111010",29589 => "01001101",29590 => "11011110",29591 => "00110101",29592 => "11011100",29593 => "11111000",29594 => "10101000",29595 => "10000011",29596 => "10011111",29597 => "10110000",29598 => "11100010",29599 => "00110001",29600 => "00111111",29601 => "11000011",29602 => "10001011",29603 => "10101111",29604 => "01110000",29605 => "01110001",29606 => "00011010",29607 => "00010100",29608 => "11010100",29609 => "11000111",29610 => "10110111",29611 => "00001000",29612 => "10110100",29613 => "10101100",29614 => "00001000",29615 => "11000001",29616 => "00100010",29617 => "10000010",29618 => "11010100",29619 => "10110011",29620 => "01100001",29621 => "11110000",29622 => "10101101",29623 => "11011111",29624 => "10010000",29625 => "10001111",29626 => "01111000",29627 => "01110011",29628 => "10100001",29629 => "01001000",29630 => "10111100",29631 => "11000001",29632 => "11010101",29633 => "00000110",29634 => "01001111",29635 => "11001000",29636 => "00000110",29637 => "11100010",29638 => "00001111",29639 => "10000011",29640 => "00101111",29641 => "01110011",29642 => "11001111",29643 => "00010101",29644 => "11000101",29645 => "01011010",29646 => "00010111",29647 => "10001101",29648 => "10111011",29649 => "00111001",29650 => "01011010",29651 => "11111000",29652 => "01100110",29653 => "01010000",29654 => "11100010",29655 => "11101101",29656 => "11001001",29657 => "00010101",29658 => "11000011",29659 => "00011011",29660 => "11111011",29661 => "11000111",29662 => "10010110",29663 => "00000101",29664 => "11101111",29665 => "01011001",29666 => "01110010",29667 => "10011001",29668 => "10001001",29669 => "00101100",29670 => "10001111",29671 => "01000010",29672 => "01111010",29673 => "10111111",29674 => "00001101",29675 => "11111011",29676 => "11100001",29677 => "00111111",29678 => "10100110",29679 => "00000001",29680 => "10000100",29681 => "10111110",29682 => "01111000",29683 => "10000101",29684 => "01110100",29685 => "11010100",29686 => "01001010",29687 => "00000011",29688 => "00100101",29689 => "00011010",29690 => "11000010",29691 => "00010011",29692 => "00100101",29693 => "10000110",29694 => "00111000",29695 => "10111001",29696 => "10100010",29697 => "00010111",29698 => "01101011",29699 => "10111100",29700 => "11010110",29701 => "00100101",29702 => "11110101",29703 => "01101011",29704 => "00000111",29705 => "00011111",29706 => "01001100",29707 => "10001001",29708 => "10000111",29709 => "00110110",29710 => "01111111",29711 => "01100001",29712 => "11000100",29713 => "01110101",29714 => "10000110",29715 => "10001111",29716 => "11010011",29717 => "11110101",29718 => "11110000",29719 => "01010101",29720 => "01011010",29721 => "10111010",29722 => "01100101",29723 => "11010000",29724 => "00000111",29725 => "10110000",29726 => "01111000",29727 => "01101100",29728 => "00110010",29729 => "11100101",29730 => "01001001",29731 => "10011000",29732 => "00001101",29733 => "00100010",29734 => "11001011",29735 => "01111000",29736 => "01011101",29737 => "11111101",29738 => "10000000",29739 => "10011101",29740 => "00011010",29741 => "01111000",29742 => "10110001",29743 => "11110101",29744 => "11110100",29745 => "11001111",29746 => "11111101",29747 => "01010010",29748 => "01001101",29749 => "10001011",29750 => "01100101",29751 => "10011011",29752 => "01101101",29753 => "00100101",29754 => "01000100",29755 => "00011010",29756 => "00110011",29757 => "10011000",29758 => "10100100",29759 => "01000101",29760 => "10000100",29761 => "00011010",29762 => "01101111",29763 => "01000010",29764 => "00010101",29765 => "00011110",29766 => "10011100",29767 => "00101110",29768 => "00001111",29769 => "10001011",29770 => "01100110",29771 => "10100011",29772 => "10001000",29773 => "11011110",29774 => "10010011",29775 => "00110100",29776 => "00000010",29777 => "10101001",29778 => "01100101",29779 => "11001111",29780 => "00110110",29781 => "01100000",29782 => "00100100",29783 => "11101001",29784 => "11011110",29785 => "00001111",29786 => "01100110",29787 => "01001111",29788 => "11000100",29789 => "00110011",29790 => "10110110",29791 => "11001010",29792 => "00111010",29793 => "11111000",29794 => "10111110",29795 => "01011111",29796 => "10101100",29797 => "01100101",29798 => "01101100",29799 => "00110101",29800 => "11000100",29801 => "10110010",29802 => "11110011",29803 => "01110101",29804 => "01110011",29805 => "10000001",29806 => "10000010",29807 => "00110001",29808 => "11011011",29809 => "10011111",29810 => "00000010",29811 => "10110000",29812 => "11110110",29813 => "01011101",29814 => "10011011",29815 => "10010111",29816 => "10011001",29817 => "11001101",29818 => "01011110",29819 => "01110100",29820 => "11110001",29821 => "00000111",29822 => "10111000",29823 => "11001010",29824 => "01100100",29825 => "00001010",29826 => "01010111",29827 => "01011100",29828 => "00000000",29829 => "10010011",29830 => "11100110",29831 => "11000011",29832 => "10110000",29833 => "01000111",29834 => "10011101",29835 => "00010001",29836 => "10010100",29837 => "11111101",29838 => "11111011",29839 => "11111111",29840 => "10010001",29841 => "00000111",29842 => "00111001",29843 => "11001000",29844 => "11011010",29845 => "10111011",29846 => "01011010",29847 => "11101000",29848 => "00000001",29849 => "11100011",29850 => "01101000",29851 => "11101101",29852 => "11101110",29853 => "01010111",29854 => "11110100",29855 => "01101011",29856 => "11111110",29857 => "10010001",29858 => "00100011",29859 => "10110011",29860 => "10000110",29861 => "11010000",29862 => "11001111",29863 => "10111001",29864 => "10010000",29865 => "01100000",29866 => "00011010",29867 => "00001111",29868 => "10111001",29869 => "10010110",29870 => "01011000",29871 => "01111100",29872 => "00101000",29873 => "01001001",29874 => "10010010",29875 => "00101101",29876 => "11110110",29877 => "10001011",29878 => "01101011",29879 => "01101001",29880 => "00011000",29881 => "11011010",29882 => "11101100",29883 => "00110001",29884 => "00111100",29885 => "10101111",29886 => "10101110",29887 => "00100100",29888 => "11100011",29889 => "10001010",29890 => "11111010",29891 => "00011001",29892 => "01011101",29893 => "01100010",29894 => "11010000",29895 => "11100110",29896 => "10011110",29897 => "11110101",29898 => "01010110",29899 => "00111110",29900 => "10101000",29901 => "11010001",29902 => "11110011",29903 => "01101101",29904 => "11111011",29905 => "10101011",29906 => "11000100",29907 => "01111111",29908 => "11011100",29909 => "10010100",29910 => "11011011",29911 => "11001101",29912 => "00101000",29913 => "01101110",29914 => "11100101",29915 => "10010010",29916 => "11110101",29917 => "00110001",29918 => "10001001",29919 => "10101011",29920 => "11000111",29921 => "10110001",29922 => "10011100",29923 => "10101110",29924 => "10111100",29925 => "11000001",29926 => "01010110",29927 => "10100011",29928 => "01010101",29929 => "11100001",29930 => "00000110",29931 => "10101111",29932 => "10000110",29933 => "10110001",29934 => "10100010",29935 => "10001010",29936 => "11001000",29937 => "00011100",29938 => "00011110",29939 => "11000010",29940 => "00110001",29941 => "01101101",29942 => "01110011",29943 => "10100111",29944 => "10101110",29945 => "10000000",29946 => "00100101",29947 => "00010111",29948 => "11010101",29949 => "11110010",29950 => "00101100",29951 => "00101011",29952 => "01110000",29953 => "11010001",29954 => "01111010",29955 => "10001110",29956 => "00110001",29957 => "00011101",29958 => "11001000",29959 => "10100000",29960 => "11001101",29961 => "11100011",29962 => "01110011",29963 => "00110100",29964 => "00111111",29965 => "10010100",29966 => "00010000",29967 => "01010100",29968 => "10010101",29969 => "10010110",29970 => "11001101",29971 => "11011011",29972 => "01010010",29973 => "11001110",29974 => "11000001",29975 => "00101000",29976 => "11100110",29977 => "10001110",29978 => "00011011",29979 => "11111001",29980 => "11100010",29981 => "01011000",29982 => "10111100",29983 => "01111111",29984 => "11001001",29985 => "11100101",29986 => "11110101",29987 => "11110000",29988 => "00010111",29989 => "00001110",29990 => "10001001",29991 => "00011010",29992 => "01111111",29993 => "01100001",29994 => "10110100",29995 => "00110001",29996 => "01100001",29997 => "11110101",29998 => "00100111",29999 => "11101000",30000 => "11101011",30001 => "01010110",30002 => "10111110",30003 => "11001001",30004 => "00000011",30005 => "11110010",30006 => "00110001",30007 => "00010001",30008 => "11000010",30009 => "11000110",30010 => "10110000",30011 => "00101010",30012 => "10011111",30013 => "11001110",30014 => "10011000",30015 => "01110000",30016 => "00000110",30017 => "01000110",30018 => "00100010",30019 => "00101010",30020 => "01001100",30021 => "11110110",30022 => "10001001",30023 => "11000110",30024 => "10011110",30025 => "01110001",30026 => "00101011",30027 => "00011101",30028 => "01101111",30029 => "01000101",30030 => "01000001",30031 => "00011011",30032 => "11001000",30033 => "01000011",30034 => "10110000",30035 => "01100001",30036 => "10111110",30037 => "00100011",30038 => "10100000",30039 => "11101110",30040 => "01101100",30041 => "10100000",30042 => "00000100",30043 => "11101010",30044 => "10010100",30045 => "01101000",30046 => "00111000",30047 => "01011001",30048 => "11110100",30049 => "01001110",30050 => "00001001",30051 => "00111000",30052 => "10000000",30053 => "00011000",30054 => "10100001",30055 => "01011101",30056 => "10000111",30057 => "10011001",30058 => "01001101",30059 => "10001101",30060 => "11011000",30061 => "01000001",30062 => "01000100",30063 => "00101111",30064 => "11001110",30065 => "11101101",30066 => "10100010",30067 => "11101111",30068 => "11100111",30069 => "10000111",30070 => "00000010",30071 => "11000101",30072 => "10100100",30073 => "10110101",30074 => "01001011",30075 => "10010011",30076 => "11010100",30077 => "11001011",30078 => "00101110",30079 => "11101000",30080 => "00100110",30081 => "11111100",30082 => "00000110",30083 => "01110000",30084 => "10010100",30085 => "00101100",30086 => "00001000",30087 => "10000101",30088 => "01111010",30089 => "10100110",30090 => "11000101",30091 => "00010000",30092 => "10011010",30093 => "01100101",30094 => "10101110",30095 => "01010100",30096 => "01001101",30097 => "01001101",30098 => "11110010",30099 => "01001010",30100 => "10100001",30101 => "01000101",30102 => "11011010",30103 => "10111011",30104 => "00101000",30105 => "00000000",30106 => "00100110",30107 => "01111000",30108 => "01110001",30109 => "00001011",30110 => "11010100",30111 => "00110011",30112 => "00100011",30113 => "10001010",30114 => "10010011",30115 => "11001000",30116 => "00011000",30117 => "01001100",30118 => "11101100",30119 => "11011101",30120 => "10100101",30121 => "01011011",30122 => "00100000",30123 => "10110001",30124 => "00010011",30125 => "01101001",30126 => "10110001",30127 => "10001111",30128 => "11000100",30129 => "10110101",30130 => "01111001",30131 => "00000110",30132 => "00110010",30133 => "00110010",30134 => "10001110",30135 => "10110010",30136 => "00101110",30137 => "01110000",30138 => "01110100",30139 => "10011001",30140 => "01100011",30141 => "11100011",30142 => "11110010",30143 => "10101010",30144 => "00101001",30145 => "01010111",30146 => "11111010",30147 => "01101001",30148 => "11101010",30149 => "01000110",30150 => "11100010",30151 => "01111101",30152 => "00001011",30153 => "10100111",30154 => "11001010",30155 => "11111110",30156 => "11000101",30157 => "10111000",30158 => "10110000",30159 => "10101000",30160 => "01000010",30161 => "10011101",30162 => "10101010",30163 => "11011101",30164 => "11110000",30165 => "10100010",30166 => "10011000",30167 => "00000111",30168 => "11011101",30169 => "10011101",30170 => "01100100",30171 => "00101111",30172 => "11101111",30173 => "01001110",30174 => "11001001",30175 => "01011110",30176 => "11011101",30177 => "10000101",30178 => "10010101",30179 => "01011010",30180 => "00010101",30181 => "01011010",30182 => "11101010",30183 => "01101011",30184 => "11000000",30185 => "10101001",30186 => "01101101",30187 => "00000111",30188 => "01000101",30189 => "11111010",30190 => "10101010",30191 => "01111011",30192 => "00101001",30193 => "10110010",30194 => "01010011",30195 => "10111100",30196 => "00011110",30197 => "00000010",30198 => "11011110",30199 => "01101001",30200 => "10100100",30201 => "11001101",30202 => "11100011",30203 => "11011111",30204 => "10100010",30205 => "00110010",30206 => "01101001",30207 => "00001010",30208 => "00010000",30209 => "01100000",30210 => "01110011",30211 => "10001001",30212 => "11000101",30213 => "01010100",30214 => "10010010",30215 => "11001110",30216 => "00101110",30217 => "00110010",30218 => "00001001",30219 => "00110010",30220 => "01001010",30221 => "01101101",30222 => "01011000",30223 => "10010011",30224 => "00111010",30225 => "10001111",30226 => "01010101",30227 => "10000101",30228 => "11011010",30229 => "11100011",30230 => "01000011",30231 => "10010010",30232 => "00011001",30233 => "10111100",30234 => "01000100",30235 => "11010011",30236 => "11110000",30237 => "01110001",30238 => "11001011",30239 => "10010001",30240 => "10110100",30241 => "10001011",30242 => "11010111",30243 => "01010011",30244 => "11110001",30245 => "00011001",30246 => "00110010",30247 => "00001000",30248 => "00000000",30249 => "10001110",30250 => "00111110",30251 => "11001011",30252 => "11000100",30253 => "11110111",30254 => "11011100",30255 => "11110101",30256 => "10101100",30257 => "01101111",30258 => "00110001",30259 => "01001101",30260 => "10100101",30261 => "01100110",30262 => "01001001",30263 => "11101101",30264 => "10110100",30265 => "01110111",30266 => "11101110",30267 => "00000011",30268 => "00100100",30269 => "10001100",30270 => "10011101",30271 => "00111000",30272 => "11000110",30273 => "11111101",30274 => "00101001",30275 => "00101010",30276 => "00110100",30277 => "01101001",30278 => "10101101",30279 => "01100011",30280 => "10011111",30281 => "01101001",30282 => "11010010",30283 => "10101111",30284 => "11110010",30285 => "10101111",30286 => "01001010",30287 => "00001010",30288 => "11100111",30289 => "01100001",30290 => "01110101",30291 => "01111010",30292 => "10010011",30293 => "11010000",30294 => "00100010",30295 => "11101001",30296 => "01111111",30297 => "00010100",30298 => "10000110",30299 => "11010111",30300 => "00110110",30301 => "01001001",30302 => "11001101",30303 => "01010111",30304 => "01011100",30305 => "10000111",30306 => "11111101",30307 => "10101010",30308 => "10111110",30309 => "01110111",30310 => "01101011",30311 => "00100000",30312 => "01111110",30313 => "00001010",30314 => "00001100",30315 => "10101001",30316 => "10010000",30317 => "10100001",30318 => "10111100",30319 => "11010010",30320 => "10010001",30321 => "00000010",30322 => "00100001",30323 => "10000100",30324 => "00000010",30325 => "11000011",30326 => "00101011",30327 => "01000011",30328 => "11101010",30329 => "10101110",30330 => "10111111",30331 => "01110100",30332 => "11000100",30333 => "11101000",30334 => "00110000",30335 => "10010100",30336 => "10001000",30337 => "11000110",30338 => "11110111",30339 => "00000000",30340 => "00101100",30341 => "01110111",30342 => "00000100",30343 => "00010000",30344 => "00100100",30345 => "11100011",30346 => "11010100",30347 => "10000011",30348 => "11110111",30349 => "10000011",30350 => "01011011",30351 => "01000100",30352 => "10001011",30353 => "10010110",30354 => "01010001",30355 => "01011010",30356 => "00011111",30357 => "00010000",30358 => "00001010",30359 => "01000000",30360 => "01000001",30361 => "01101011",30362 => "00000000",30363 => "11010001",30364 => "11101111",30365 => "11100000",30366 => "00000110",30367 => "11111011",30368 => "01110110",30369 => "10011001",30370 => "10111111",30371 => "01011011",30372 => "01100011",30373 => "11000000",30374 => "00000010",30375 => "11001100",30376 => "00100101",30377 => "10111101",30378 => "00111100",30379 => "01111100",30380 => "10110110",30381 => "01010101",30382 => "00010010",30383 => "00101111",30384 => "01101101",30385 => "00101011",30386 => "10100101",30387 => "00111010",30388 => "11001111",30389 => "00111000",30390 => "10110110",30391 => "11110011",30392 => "10101110",30393 => "10010000",30394 => "10000000",30395 => "00001010",30396 => "11101100",30397 => "11011100",30398 => "10011111",30399 => "10010101",30400 => "11111001",30401 => "00011110",30402 => "01010110",30403 => "11110100",30404 => "10011101",30405 => "00001110",30406 => "00110101",30407 => "10011101",30408 => "11011100",30409 => "00111100",30410 => "00010001",30411 => "11101100",30412 => "00010100",30413 => "11001001",30414 => "11011010",30415 => "11100011",30416 => "10010001",30417 => "00110000",30418 => "01101100",30419 => "01101101",30420 => "11101000",30421 => "10111011",30422 => "10000111",30423 => "11001001",30424 => "01010110",30425 => "11000010",30426 => "00110010",30427 => "00100101",30428 => "01010010",30429 => "01101010",30430 => "00101000",30431 => "11011011",30432 => "10110100",30433 => "10011000",30434 => "11011011",30435 => "01101100",30436 => "00111011",30437 => "00110101",30438 => "01110110",30439 => "10111010",30440 => "01111100",30441 => "11010000",30442 => "11101111",30443 => "11110011",30444 => "11111100",30445 => "01101110",30446 => "01110000",30447 => "10111110",30448 => "00110110",30449 => "11111111",30450 => "11001010",30451 => "01100000",30452 => "10101101",30453 => "00011000",30454 => "00000011",30455 => "11110011",30456 => "01011101",30457 => "11101101",30458 => "01111101",30459 => "11111010",30460 => "10111011",30461 => "01110101",30462 => "01110110",30463 => "11111011",30464 => "00100001",30465 => "11001010",30466 => "01111100",30467 => "01101010",30468 => "01000010",30469 => "01011000",30470 => "11101110",30471 => "00010000",30472 => "11010110",30473 => "11100110",30474 => "11110100",30475 => "11010001",30476 => "10001111",30477 => "11011011",30478 => "11001101",30479 => "00010001",30480 => "10111001",30481 => "00010110",30482 => "00001011",30483 => "10100101",30484 => "01001110",30485 => "01000000",30486 => "01010011",30487 => "01100100",30488 => "00111000",30489 => "01011011",30490 => "00111101",30491 => "00111010",30492 => "01010000",30493 => "10011011",30494 => "00001001",30495 => "11101001",30496 => "01101011",30497 => "01011100",30498 => "11100011",30499 => "11100111",30500 => "01110111",30501 => "01100010",30502 => "11100101",30503 => "01010100",30504 => "01111001",30505 => "11101110",30506 => "00111011",30507 => "01111000",30508 => "10100001",30509 => "11111010",30510 => "10110100",30511 => "11100000",30512 => "10000000",30513 => "11001110",30514 => "01101101",30515 => "10000011",30516 => "01000110",30517 => "10101110",30518 => "10101011",30519 => "01011001",30520 => "00111010",30521 => "10101010",30522 => "10000100",30523 => "10001011",30524 => "11000110",30525 => "00010101",30526 => "11100001",30527 => "01011000",30528 => "11111101",30529 => "11101110",30530 => "01011000",30531 => "00111111",30532 => "11101000",30533 => "00011011",30534 => "01101001",30535 => "11001110",30536 => "00110011",30537 => "11110110",30538 => "10100010",30539 => "10011011",30540 => "10101101",30541 => "11111100",30542 => "00010010",30543 => "10101000",30544 => "01011111",30545 => "00011111",30546 => "00010101",30547 => "00100001",30548 => "01001011",30549 => "11000000",30550 => "00000000",30551 => "10111010",30552 => "01010100",30553 => "11110010",30554 => "11010111",30555 => "01011111",30556 => "11110011",30557 => "10011011",30558 => "11111111",30559 => "10100001",30560 => "10110010",30561 => "01000101",30562 => "01011011",30563 => "00100011",30564 => "11101010",30565 => "01001000",30566 => "11001010",30567 => "10010111",30568 => "10000100",30569 => "00000001",30570 => "00000100",30571 => "10101000",30572 => "11011000",30573 => "11110100",30574 => "00100111",30575 => "01101111",30576 => "11101100",30577 => "00111110",30578 => "01010100",30579 => "00111010",30580 => "01010100",30581 => "10010011",30582 => "00101001",30583 => "11011100",30584 => "11011001",30585 => "00101001",30586 => "00111100",30587 => "10001011",30588 => "00010000",30589 => "01001110",30590 => "10010111",30591 => "00010101",30592 => "10100000",30593 => "00001001",30594 => "10100111",30595 => "11101101",30596 => "01001111",30597 => "11010010",30598 => "01011100",30599 => "11110010",30600 => "10100010",30601 => "11001100",30602 => "11010101",30603 => "10100010",30604 => "11101000",30605 => "01011000",30606 => "01110101",30607 => "01010110",30608 => "00101111",30609 => "11111100",30610 => "11000101",30611 => "11001101",30612 => "10100010",30613 => "01011100",30614 => "00000101",30615 => "10000001",30616 => "11001111",30617 => "11101100",30618 => "10101101",30619 => "11100000",30620 => "01100001",30621 => "01011011",30622 => "01011000",30623 => "10110011",30624 => "01101010",30625 => "10101001",30626 => "11110111",30627 => "01001101",30628 => "01010100",30629 => "11101010",30630 => "10000111",30631 => "11100110",30632 => "11110001",30633 => "10001000",30634 => "10011101",30635 => "11111100",30636 => "11011101",30637 => "10111011",30638 => "00010110",30639 => "00010111",30640 => "10101010",30641 => "11011000",30642 => "01100100",30643 => "01000101",30644 => "11101000",30645 => "01110101",30646 => "01011110",30647 => "11101001",30648 => "00111100",30649 => "00001000",30650 => "10010010",30651 => "10111011",30652 => "11111101",30653 => "00111011",30654 => "00011000",30655 => "11101001",30656 => "00011000",30657 => "01111100",30658 => "11101111",30659 => "10101111",30660 => "00010111",30661 => "11110111",30662 => "01111100",30663 => "00100110",30664 => "10111010",30665 => "00011011",30666 => "11111000",30667 => "11111011",30668 => "00101000",30669 => "00110011",30670 => "01011100",30671 => "00101011",30672 => "11101101",30673 => "10010111",30674 => "00100110",30675 => "10011011",30676 => "11010011",30677 => "11011011",30678 => "00001111",30679 => "01101110",30680 => "00011101",30681 => "01000111",30682 => "01111111",30683 => "11100001",30684 => "00010001",30685 => "11111011",30686 => "11111010",30687 => "10000001",30688 => "01000011",30689 => "10101111",30690 => "01011110",30691 => "01010101",30692 => "01000000",30693 => "11110010",30694 => "00101101",30695 => "11011101",30696 => "10101000",30697 => "01011001",30698 => "01100111",30699 => "01010111",30700 => "01111010",30701 => "01110011",30702 => "01011100",30703 => "10100111",30704 => "11101100",30705 => "01101110",30706 => "00100100",30707 => "00110011",30708 => "00001110",30709 => "00000010",30710 => "10110000",30711 => "11110000",30712 => "00111100",30713 => "00110011",30714 => "00110110",30715 => "10111000",30716 => "10100110",30717 => "11100000",30718 => "00001101",30719 => "10110110",30720 => "01111001",30721 => "11101001",30722 => "00000011",30723 => "11011111",30724 => "10000110",30725 => "10100010",30726 => "00010000",30727 => "00110101",30728 => "00100100",30729 => "01101110",30730 => "01100110",30731 => "11101111",30732 => "10100101",30733 => "11111000",30734 => "01001110",30735 => "10000000",30736 => "01101100",30737 => "11010001",30738 => "00010011",30739 => "01001001",30740 => "11111010",30741 => "00011111",30742 => "10011101",30743 => "01111011",30744 => "00010000",30745 => "00001101",30746 => "11100011",30747 => "10101010",30748 => "11011101",30749 => "10010001",30750 => "10000011",30751 => "01101101",30752 => "00010101",30753 => "01000111",30754 => "10111110",30755 => "11101110",30756 => "00110010",30757 => "01010000",30758 => "11111001",30759 => "01000101",30760 => "00011001",30761 => "00000001",30762 => "10000000",30763 => "10111001",30764 => "01101000",30765 => "11011101",30766 => "10100111",30767 => "00110100",30768 => "00100101",30769 => "00110111",30770 => "00011100",30771 => "01000000",30772 => "10000001",30773 => "11000010",30774 => "11111110",30775 => "00110000",30776 => "10000101",30777 => "10011100",30778 => "01001010",30779 => "10011010",30780 => "01110100",30781 => "01110001",30782 => "01001010",30783 => "01101100",30784 => "10110001",30785 => "00001000",30786 => "10110101",30787 => "01111000",30788 => "01010100",30789 => "01010011",30790 => "01010011",30791 => "01001101",30792 => "11011101",30793 => "01000001",30794 => "01111111",30795 => "00101101",30796 => "01011100",30797 => "01100100",30798 => "10100101",30799 => "11100000",30800 => "00001001",30801 => "10110100",30802 => "01000100",30803 => "11111101",30804 => "11100000",30805 => "11001100",30806 => "00010110",30807 => "11100101",30808 => "10100100",30809 => "10000100",30810 => "00001011",30811 => "10000000",30812 => "00110001",30813 => "01001000",30814 => "01011010",30815 => "00111011",30816 => "01001111",30817 => "01010110",30818 => "10110010",30819 => "00110011",30820 => "10110100",30821 => "11111011",30822 => "11001110",30823 => "10111101",30824 => "01001000",30825 => "00101001",30826 => "00100111",30827 => "10111011",30828 => "01110101",30829 => "11000001",30830 => "00111010",30831 => "10110110",30832 => "10001011",30833 => "00010001",30834 => "11101101",30835 => "01100000",30836 => "10101011",30837 => "00100101",30838 => "01001001",30839 => "01011001",30840 => "10100100",30841 => "11000101",30842 => "10111110",30843 => "00001001",30844 => "10011000",30845 => "01110001",30846 => "00011010",30847 => "00100100",30848 => "11110010",30849 => "10100111",30850 => "10011110",30851 => "11111101",30852 => "01100011",30853 => "00110110",30854 => "11100101",30855 => "10110110",30856 => "01000110",30857 => "10010111",30858 => "11111001",30859 => "01101100",30860 => "10011001",30861 => "01101010",30862 => "10100101",30863 => "01010111",30864 => "11110000",30865 => "01111001",30866 => "11000110",30867 => "01001000",30868 => "00101011",30869 => "00010010",30870 => "01100101",30871 => "10100001",30872 => "01100100",30873 => "10100111",30874 => "01011101",30875 => "10111011",30876 => "01111011",30877 => "10010010",30878 => "00100101",30879 => "10111100",30880 => "00000010",30881 => "11110111",30882 => "01111101",30883 => "01000101",30884 => "00111000",30885 => "11110100",30886 => "10110110",30887 => "11100001",30888 => "10010100",30889 => "11010100",30890 => "00010101",30891 => "01000000",30892 => "01111110",30893 => "01000011",30894 => "00101100",30895 => "00100010",30896 => "01000101",30897 => "00011110",30898 => "01101110",30899 => "10101001",30900 => "00101100",30901 => "01000010",30902 => "01010111",30903 => "11011100",30904 => "10111110",30905 => "11011010",30906 => "10010011",30907 => "01000100",30908 => "10001110",30909 => "10011010",30910 => "00011000",30911 => "01010111",30912 => "00001100",30913 => "11011100",30914 => "11110101",30915 => "11110111",30916 => "10111000",30917 => "11101101",30918 => "10101001",30919 => "11010101",30920 => "11100010",30921 => "10011101",30922 => "00110101",30923 => "01101101",30924 => "11100000",30925 => "11010001",30926 => "10001111",30927 => "01001000",30928 => "11001110",30929 => "00001100",30930 => "01111110",30931 => "01011010",30932 => "00110001",30933 => "11110010",30934 => "10100001",30935 => "00001010",30936 => "11011010",30937 => "01000110",30938 => "11001101",30939 => "00111011",30940 => "10111010",30941 => "11110001",30942 => "10011000",30943 => "11101001",30944 => "01011100",30945 => "10101000",30946 => "10001110",30947 => "00101111",30948 => "00100111",30949 => "11001111",30950 => "10110001",30951 => "10011101",30952 => "01001000",30953 => "11011011",30954 => "01100011",30955 => "00110100",30956 => "11000111",30957 => "01111010",30958 => "01110001",30959 => "00101111",30960 => "11110010",30961 => "01000010",30962 => "00101011",30963 => "00000111",30964 => "00100111",30965 => "01111010",30966 => "11001101",30967 => "11011111",30968 => "01011110",30969 => "11000011",30970 => "10111110",30971 => "01001101",30972 => "11111001",30973 => "01111010",30974 => "01001110",30975 => "00111111",30976 => "10111011",30977 => "11110000",30978 => "11001000",30979 => "10011011",30980 => "00000011",30981 => "11100100",30982 => "00111011",30983 => "00100100",30984 => "11001001",30985 => "00101000",30986 => "10010100",30987 => "10010100",30988 => "01111111",30989 => "00001010",30990 => "01011011",30991 => "11110010",30992 => "10100001",30993 => "00011111",30994 => "01100110",30995 => "00100000",30996 => "10001010",30997 => "00111000",30998 => "01101000",30999 => "00000000",31000 => "11000010",31001 => "00011011",31002 => "00000110",31003 => "00110010",31004 => "10110001",31005 => "00101111",31006 => "00101111",31007 => "01010000",31008 => "00111111",31009 => "10010010",31010 => "11101101",31011 => "01010010",31012 => "11100000",31013 => "10011010",31014 => "01000100",31015 => "10110010",31016 => "00011011",31017 => "00111110",31018 => "11110000",31019 => "10111110",31020 => "00110101",31021 => "01111100",31022 => "00011101",31023 => "00011001",31024 => "10101110",31025 => "10101101",31026 => "10101000",31027 => "10101000",31028 => "11011011",31029 => "00101000",31030 => "10100110",31031 => "00100100",31032 => "10011110",31033 => "00001010",31034 => "10110101",31035 => "00010011",31036 => "01011100",31037 => "11111000",31038 => "00111111",31039 => "10101100",31040 => "01101111",31041 => "11011110",31042 => "00101101",31043 => "10000101",31044 => "00110100",31045 => "10001110",31046 => "01110100",31047 => "00000111",31048 => "10000011",31049 => "10010001",31050 => "11111000",31051 => "11101001",31052 => "11000110",31053 => "10010111",31054 => "11110011",31055 => "11110110",31056 => "11010100",31057 => "11100111",31058 => "10011000",31059 => "00101100",31060 => "01011001",31061 => "01000111",31062 => "10000110",31063 => "11101001",31064 => "01110110",31065 => "00011110",31066 => "00110100",31067 => "01000111",31068 => "00010011",31069 => "11110111",31070 => "00111101",31071 => "11100001",31072 => "00110110",31073 => "11101100",31074 => "10010011",31075 => "01010110",31076 => "01101101",31077 => "01011011",31078 => "00000000",31079 => "01001110",31080 => "11100011",31081 => "01111111",31082 => "11100010",31083 => "10111010",31084 => "01001110",31085 => "11001111",31086 => "10101111",31087 => "00111000",31088 => "11110101",31089 => "11000011",31090 => "10110000",31091 => "01110010",31092 => "10101100",31093 => "00100000",31094 => "11101100",31095 => "11100011",31096 => "00100000",31097 => "11111010",31098 => "00010101",31099 => "10011001",31100 => "10110010",31101 => "10001100",31102 => "00110011",31103 => "11011010",31104 => "00000000",31105 => "11101001",31106 => "11100011",31107 => "00001100",31108 => "11010001",31109 => "00001111",31110 => "00000101",31111 => "11100110",31112 => "01111101",31113 => "10001100",31114 => "00010101",31115 => "10101111",31116 => "11000111",31117 => "01100100",31118 => "01000011",31119 => "10110100",31120 => "10100011",31121 => "11100111",31122 => "00111101",31123 => "11001001",31124 => "10110110",31125 => "11110100",31126 => "01011010",31127 => "01000101",31128 => "01101111",31129 => "00101110",31130 => "00010101",31131 => "01011100",31132 => "11101000",31133 => "01101000",31134 => "01111011",31135 => "11110101",31136 => "11000010",31137 => "10100100",31138 => "01011000",31139 => "11111100",31140 => "00110010",31141 => "11110000",31142 => "10111000",31143 => "10101000",31144 => "01000001",31145 => "10010011",31146 => "01101101",31147 => "00100110",31148 => "00100011",31149 => "01100111",31150 => "11110001",31151 => "11110011",31152 => "01101110",31153 => "01100110",31154 => "01000110",31155 => "01001110",31156 => "10001111",31157 => "10110001",31158 => "11100111",31159 => "10010110",31160 => "10101011",31161 => "01111001",31162 => "11000110",31163 => "00110010",31164 => "11000101",31165 => "01001000",31166 => "11101101",31167 => "00110101",31168 => "00100110",31169 => "10000010",31170 => "10001110",31171 => "10010000",31172 => "11010000",31173 => "00111000",31174 => "01100010",31175 => "00101101",31176 => "00000111",31177 => "11110110",31178 => "01110001",31179 => "10101011",31180 => "11001000",31181 => "01110101",31182 => "10100001",31183 => "11110100",31184 => "10001111",31185 => "11000010",31186 => "01101100",31187 => "10011000",31188 => "10010111",31189 => "11110010",31190 => "01100100",31191 => "00000011",31192 => "01010011",31193 => "00110000",31194 => "00000001",31195 => "11110000",31196 => "11101100",31197 => "10000100",31198 => "01010101",31199 => "10000101",31200 => "10100111",31201 => "00000100",31202 => "00000101",31203 => "01010110",31204 => "01101010",31205 => "10111101",31206 => "11101111",31207 => "11011100",31208 => "00111100",31209 => "01100110",31210 => "00111011",31211 => "11011100",31212 => "00000111",31213 => "10101100",31214 => "10111101",31215 => "01011001",31216 => "11110101",31217 => "00110110",31218 => "10101010",31219 => "01001111",31220 => "01101011",31221 => "00101010",31222 => "10010100",31223 => "11100000",31224 => "10111111",31225 => "00011011",31226 => "11101111",31227 => "10000100",31228 => "00011111",31229 => "00010011",31230 => "01100100",31231 => "00001110",31232 => "00001111",31233 => "00011101",31234 => "11001001",31235 => "11001011",31236 => "11110101",31237 => "10011100",31238 => "01001000",31239 => "10001100",31240 => "00010000",31241 => "10100100",31242 => "00010001",31243 => "11011111",31244 => "10011000",31245 => "10110111",31246 => "01000110",31247 => "00110111",31248 => "11100010",31249 => "01100101",31250 => "10000101",31251 => "11100000",31252 => "11011111",31253 => "10001101",31254 => "00000011",31255 => "00100001",31256 => "01000001",31257 => "11010011",31258 => "10011111",31259 => "01010100",31260 => "11011010",31261 => "11011011",31262 => "01011100",31263 => "10001111",31264 => "01100110",31265 => "00111000",31266 => "01101101",31267 => "00111111",31268 => "00001010",31269 => "10010011",31270 => "01001110",31271 => "01101101",31272 => "00110010",31273 => "01111000",31274 => "10011110",31275 => "01001101",31276 => "10010001",31277 => "00010110",31278 => "10100100",31279 => "00111010",31280 => "00000101",31281 => "11001000",31282 => "01110010",31283 => "00101111",31284 => "00100010",31285 => "00010110",31286 => "11001010",31287 => "01100101",31288 => "00110011",31289 => "01100100",31290 => "10100101",31291 => "10100110",31292 => "10000001",31293 => "01100100",31294 => "00010011",31295 => "11000011",31296 => "00101001",31297 => "11111100",31298 => "11001011",31299 => "11001010",31300 => "10111000",31301 => "00100000",31302 => "00001000",31303 => "01101000",31304 => "10110011",31305 => "00111110",31306 => "10011110",31307 => "00011111",31308 => "00011101",31309 => "11100110",31310 => "01010000",31311 => "11111000",31312 => "00011010",31313 => "10010000",31314 => "01100011",31315 => "10010101",31316 => "00110000",31317 => "00000110",31318 => "01011110",31319 => "01000010",31320 => "01011000",31321 => "11111110",31322 => "01101110",31323 => "01110000",31324 => "01101111",31325 => "10000011",31326 => "01110110",31327 => "11111100",31328 => "11100010",31329 => "00010100",31330 => "10000001",31331 => "11011011",31332 => "11101100",31333 => "00001111",31334 => "00101000",31335 => "10000110",31336 => "00010001",31337 => "00110000",31338 => "10111011",31339 => "01001101",31340 => "00110110",31341 => "00011101",31342 => "10111010",31343 => "00110100",31344 => "00001010",31345 => "01101111",31346 => "01010110",31347 => "00010000",31348 => "01011101",31349 => "10001111",31350 => "01001111",31351 => "10111011",31352 => "01010100",31353 => "10111111",31354 => "11100101",31355 => "00011000",31356 => "11110101",31357 => "00110101",31358 => "11011111",31359 => "11001011",31360 => "10001000",31361 => "11011001",31362 => "11110110",31363 => "00010011",31364 => "11110110",31365 => "11111101",31366 => "10110011",31367 => "10000010",31368 => "00010111",31369 => "11111000",31370 => "00000010",31371 => "01100100",31372 => "10001010",31373 => "11011001",31374 => "00111111",31375 => "10101101",31376 => "01001111",31377 => "00101011",31378 => "10110101",31379 => "10010000",31380 => "01110001",31381 => "11111011",31382 => "00010011",31383 => "11111010",31384 => "11000111",31385 => "11110010",31386 => "11001011",31387 => "00101110",31388 => "11110100",31389 => "00100001",31390 => "01011000",31391 => "11001101",31392 => "01100000",31393 => "10011000",31394 => "01110101",31395 => "01110111",31396 => "00011110",31397 => "11100000",31398 => "00111101",31399 => "00101011",31400 => "11111011",31401 => "01111111",31402 => "01110101",31403 => "01101011",31404 => "01110000",31405 => "00000100",31406 => "10000111",31407 => "01101001",31408 => "10100011",31409 => "11001111",31410 => "10110011",31411 => "11001101",31412 => "11111111",31413 => "01101111",31414 => "11100010",31415 => "11000101",31416 => "01110111",31417 => "01111000",31418 => "01001100",31419 => "11101110",31420 => "11000101",31421 => "00111110",31422 => "01000111",31423 => "01111100",31424 => "01011110",31425 => "01000000",31426 => "00001101",31427 => "01000100",31428 => "00110100",31429 => "01100010",31430 => "11101011",31431 => "10111111",31432 => "01100110",31433 => "10010010",31434 => "10010111",31435 => "11100011",31436 => "11101100",31437 => "01101100",31438 => "01010011",31439 => "10111111",31440 => "01001101",31441 => "10000111",31442 => "11101110",31443 => "11011010",31444 => "01101000",31445 => "00000010",31446 => "10111111",31447 => "01101110",31448 => "01011010",31449 => "00110110",31450 => "00000110",31451 => "10011100",31452 => "11000001",31453 => "11011111",31454 => "00000010",31455 => "11101101",31456 => "10001110",31457 => "11111101",31458 => "00100000",31459 => "10011010",31460 => "00011100",31461 => "00110111",31462 => "00111100",31463 => "01001000",31464 => "01010100",31465 => "11100110",31466 => "01111111",31467 => "10000111",31468 => "11010101",31469 => "00101101",31470 => "11011100",31471 => "00011010",31472 => "00111111",31473 => "00011111",31474 => "01111011",31475 => "01000111",31476 => "11111110",31477 => "10100110",31478 => "11011010",31479 => "00101000",31480 => "00110011",31481 => "01100011",31482 => "11011001",31483 => "10000011",31484 => "10100111",31485 => "10110100",31486 => "01100110",31487 => "01001101",31488 => "10011010",31489 => "00100001",31490 => "10100001",31491 => "10100011",31492 => "10010101",31493 => "01100011",31494 => "01110110",31495 => "00011001",31496 => "01001000",31497 => "10111101",31498 => "00110101",31499 => "00111001",31500 => "11110000",31501 => "01001010",31502 => "11000110",31503 => "01011110",31504 => "00001010",31505 => "10101111",31506 => "10110101",31507 => "01001101",31508 => "11011001",31509 => "01000101",31510 => "11000101",31511 => "01101100",31512 => "00011111",31513 => "11101111",31514 => "00001110",31515 => "00001010",31516 => "10000000",31517 => "01011001",31518 => "11000001",31519 => "11111011",31520 => "10000010",31521 => "00110010",31522 => "11010111",31523 => "00011011",31524 => "10000111",31525 => "00010110",31526 => "00000110",31527 => "11011111",31528 => "10010011",31529 => "11000101",31530 => "11100011",31531 => "10001100",31532 => "11101100",31533 => "00011101",31534 => "00000011",31535 => "01111111",31536 => "01000000",31537 => "11100101",31538 => "10100011",31539 => "11011111",31540 => "00001100",31541 => "01011101",31542 => "10011010",31543 => "11101100",31544 => "11011011",31545 => "00111011",31546 => "00011001",31547 => "11010101",31548 => "11101010",31549 => "10010011",31550 => "01001011",31551 => "11011111",31552 => "10111110",31553 => "11000101",31554 => "11010110",31555 => "00001011",31556 => "01101100",31557 => "00011010",31558 => "01001111",31559 => "10010001",31560 => "01111100",31561 => "00010001",31562 => "10110001",31563 => "00110000",31564 => "00001101",31565 => "11000011",31566 => "00100101",31567 => "01000110",31568 => "10110101",31569 => "11010001",31570 => "10010100",31571 => "11010100",31572 => "01001000",31573 => "10001110",31574 => "01011001",31575 => "00011101",31576 => "00100101",31577 => "01110111",31578 => "00001100",31579 => "10110010",31580 => "00001011",31581 => "01011001",31582 => "01010100",31583 => "11101010",31584 => "10001100",31585 => "00001000",31586 => "01000010",31587 => "01101110",31588 => "10011000",31589 => "11100110",31590 => "11111010",31591 => "01101110",31592 => "00000110",31593 => "00001110",31594 => "11100000",31595 => "11101111",31596 => "11010000",31597 => "11111011",31598 => "00110111",31599 => "01010001",31600 => "10001100",31601 => "10011110",31602 => "10111011",31603 => "10110011",31604 => "10111010",31605 => "10100100",31606 => "10011111",31607 => "00010000",31608 => "10111001",31609 => "00000000",31610 => "00100111",31611 => "01010011",31612 => "00000100",31613 => "00100101",31614 => "00010011",31615 => "01101001",31616 => "11100011",31617 => "10100011",31618 => "10101010",31619 => "10001111",31620 => "10110111",31621 => "11111011",31622 => "10001100",31623 => "11000101",31624 => "10101111",31625 => "01000101",31626 => "11011101",31627 => "00111110",31628 => "00101010",31629 => "11001010",31630 => "00001000",31631 => "10110100",31632 => "11100101",31633 => "00111001",31634 => "00010000",31635 => "11010100",31636 => "11000100",31637 => "00000010",31638 => "10110001",31639 => "00011101",31640 => "11101110",31641 => "00100001",31642 => "11001100",31643 => "00001001",31644 => "00011101",31645 => "01110001",31646 => "11110100",31647 => "01110011",31648 => "01001000",31649 => "00011101",31650 => "10010110",31651 => "01111101",31652 => "00100111",31653 => "10001100",31654 => "01001101",31655 => "10110001",31656 => "11101010",31657 => "10110011",31658 => "00100101",31659 => "00011000",31660 => "01111001",31661 => "10101100",31662 => "10011100",31663 => "11001110",31664 => "01100101",31665 => "10111000",31666 => "01001000",31667 => "10001111",31668 => "01001010",31669 => "10001010",31670 => "01111000",31671 => "01101100",31672 => "10011010",31673 => "00110110",31674 => "01011110",31675 => "00101101",31676 => "11100101",31677 => "00000100",31678 => "01010010",31679 => "11100011",31680 => "00111011",31681 => "10000000",31682 => "01100011",31683 => "10110010",31684 => "01100001",31685 => "10110010",31686 => "01010100",31687 => "01001100",31688 => "10000100",31689 => "00111011",31690 => "10000011",31691 => "00110111",31692 => "11000001",31693 => "00011101",31694 => "11010101",31695 => "10011011",31696 => "01001111",31697 => "01110100",31698 => "01101000",31699 => "10010111",31700 => "10011010",31701 => "10011001",31702 => "11011001",31703 => "11001111",31704 => "11001011",31705 => "10000001",31706 => "01011000",31707 => "11101011",31708 => "11101111",31709 => "10011010",31710 => "10010101",31711 => "00001111",31712 => "01111101",31713 => "10011100",31714 => "10100111",31715 => "11110000",31716 => "10001001",31717 => "00001010",31718 => "01110101",31719 => "00100111",31720 => "10001001",31721 => "01101101",31722 => "01100010",31723 => "10011010",31724 => "10000011",31725 => "00011110",31726 => "11110111",31727 => "10011101",31728 => "11100010",31729 => "11110000",31730 => "11011000",31731 => "10011100",31732 => "10100111",31733 => "00001001",31734 => "10011100",31735 => "01010110",31736 => "11101011",31737 => "00011101",31738 => "01000011",31739 => "10001110",31740 => "00101001",31741 => "11001111",31742 => "11110000",31743 => "11111011",31744 => "01110000",31745 => "11001111",31746 => "11011110",31747 => "00001001",31748 => "00100001",31749 => "00011111",31750 => "01111000",31751 => "00000011",31752 => "01101100",31753 => "11000111",31754 => "11010111",31755 => "11000111",31756 => "10011100",31757 => "10101111",31758 => "10100111",31759 => "00101101",31760 => "01110110",31761 => "10001000",31762 => "01100010",31763 => "00011100",31764 => "10000010",31765 => "01010011",31766 => "01100010",31767 => "10010101",31768 => "11101011",31769 => "00001110",31770 => "00000010",31771 => "11101101",31772 => "00010000",31773 => "11111111",31774 => "10100101",31775 => "00010100",31776 => "00111010",31777 => "11010100",31778 => "01111000",31779 => "11101101",31780 => "01010100",31781 => "11100010",31782 => "00010011",31783 => "11010111",31784 => "11011110",31785 => "11100110",31786 => "11111001",31787 => "10111010",31788 => "00111100",31789 => "01001011",31790 => "10110111",31791 => "10110000",31792 => "11101011",31793 => "00111010",31794 => "10101100",31795 => "10010111",31796 => "01111000",31797 => "00110011",31798 => "11011011",31799 => "10101111",31800 => "00111001",31801 => "10001000",31802 => "00100101",31803 => "01000110",31804 => "11001001",31805 => "01101001",31806 => "10000001",31807 => "01010001",31808 => "01011010",31809 => "10110111",31810 => "00000101",31811 => "10101011",31812 => "01010110",31813 => "11000011",31814 => "10111100",31815 => "11101111",31816 => "11101111",31817 => "00100011",31818 => "01110010",31819 => "10111100",31820 => "01001001",31821 => "10011111",31822 => "01001011",31823 => "01100111",31824 => "11110101",31825 => "11000000",31826 => "11010010",31827 => "11110110",31828 => "01010001",31829 => "10101101",31830 => "10101111",31831 => "10011001",31832 => "10011000",31833 => "10111100",31834 => "11111010",31835 => "11100000",31836 => "01111100",31837 => "11111101",31838 => "10101011",31839 => "10111111",31840 => "11110011",31841 => "10000110",31842 => "01001001",31843 => "01111100",31844 => "01110111",31845 => "01001000",31846 => "10001100",31847 => "00100010",31848 => "11111000",31849 => "11000010",31850 => "01101110",31851 => "00101010",31852 => "11000110",31853 => "01000100",31854 => "11110000",31855 => "01001000",31856 => "00011110",31857 => "11101010",31858 => "11011010",31859 => "00010100",31860 => "00110101",31861 => "10110001",31862 => "10100001",31863 => "01100110",31864 => "10101010",31865 => "01001000",31866 => "11101100",31867 => "01111000",31868 => "01000101",31869 => "10011010",31870 => "00010001",31871 => "10101001",31872 => "11111111",31873 => "11100011",31874 => "10000000",31875 => "01010110",31876 => "10101101",31877 => "10001011",31878 => "11101110",31879 => "00011010",31880 => "00001110",31881 => "01000000",31882 => "00001000",31883 => "00101111",31884 => "00101101",31885 => "10100010",31886 => "11100000",31887 => "00000010",31888 => "01011001",31889 => "10111010",31890 => "01110110",31891 => "10100101",31892 => "11101000",31893 => "01011000",31894 => "10111100",31895 => "01011100",31896 => "01110000",31897 => "11011110",31898 => "01110101",31899 => "00100001",31900 => "00111110",31901 => "10001110",31902 => "11001010",31903 => "10111101",31904 => "11110010",31905 => "01010100",31906 => "01110001",31907 => "10101000",31908 => "01100010",31909 => "01111101",31910 => "11101011",31911 => "10110101",31912 => "10001001",31913 => "00111110",31914 => "01100000",31915 => "01110010",31916 => "10111000",31917 => "11101010",31918 => "11110000",31919 => "01001100",31920 => "01011111",31921 => "01010111",31922 => "10011101",31923 => "10011000",31924 => "11001000",31925 => "01001010",31926 => "11100011",31927 => "11111100",31928 => "10101011",31929 => "11101111",31930 => "10001111",31931 => "00000011",31932 => "01011011",31933 => "11110010",31934 => "11111100",31935 => "10111000",31936 => "01000101",31937 => "00010100",31938 => "11001111",31939 => "01011001",31940 => "00111100",31941 => "10111111",31942 => "00100000",31943 => "00111000",31944 => "10000010",31945 => "00110100",31946 => "11001110",31947 => "01000010",31948 => "10111000",31949 => "10010000",31950 => "00011110",31951 => "11101100",31952 => "11100110",31953 => "00001011",31954 => "11000100",31955 => "01111111",31956 => "10011001",31957 => "00010110",31958 => "10100011",31959 => "00101000",31960 => "01101001",31961 => "11010010",31962 => "10010111",31963 => "00010000",31964 => "00010101",31965 => "11011001",31966 => "11111011",31967 => "00001110",31968 => "00110111",31969 => "00110011",31970 => "11001110",31971 => "11101100",31972 => "00001101",31973 => "10010001",31974 => "01000001",31975 => "11110000",31976 => "10010101",31977 => "11000000",31978 => "10000000",31979 => "01000101",31980 => "00101001",31981 => "11110110",31982 => "00001001",31983 => "11011001",31984 => "10011000",31985 => "01010101",31986 => "00111101",31987 => "01000000",31988 => "10111110",31989 => "10100010",31990 => "00010111",31991 => "10011111",31992 => "00101001",31993 => "10100011",31994 => "00111110",31995 => "11011100",31996 => "10100100",31997 => "11110011",31998 => "00000101",31999 => "00000101",32000 => "00011000",32001 => "10101101",32002 => "01010000",32003 => "11101001",32004 => "10000011",32005 => "10111111",32006 => "01011101",32007 => "10010011",32008 => "00111111",32009 => "10011000",32010 => "10011011",32011 => "10010101",32012 => "11100100",32013 => "11001110",32014 => "00011001",32015 => "11011111",32016 => "10000110",32017 => "11110101",32018 => "00001100",32019 => "11001010",32020 => "10100000",32021 => "11010010",32022 => "11101111",32023 => "01100011",32024 => "00010001",32025 => "01000000",32026 => "10101110",32027 => "01000011",32028 => "00100101",32029 => "10011100",32030 => "01000011",32031 => "01010010",32032 => "11111101",32033 => "01011011",32034 => "10010010",32035 => "01011111",32036 => "01101001",32037 => "11011100",32038 => "00110011",32039 => "10110101",32040 => "01000111",32041 => "10111000",32042 => "00011010",32043 => "00001001",32044 => "11000101",32045 => "10111110",32046 => "01111111",32047 => "10100010",32048 => "01110001",32049 => "11110001",32050 => "11100111",32051 => "00100010",32052 => "00101100",32053 => "10110010",32054 => "10000001",32055 => "01010100",32056 => "10111100",32057 => "01110000",32058 => "10110101",32059 => "10110011",32060 => "10001001",32061 => "01110100",32062 => "11111000",32063 => "10110101",32064 => "10010011",32065 => "01010111",32066 => "10111000",32067 => "00000000",32068 => "00101001",32069 => "11001100",32070 => "10101010",32071 => "10000110",32072 => "00010110",32073 => "11111001",32074 => "01111001",32075 => "01110111",32076 => "00010001",32077 => "11101010",32078 => "11010110",32079 => "01111011",32080 => "00100110",32081 => "01100111",32082 => "10011111",32083 => "00010101",32084 => "11001101",32085 => "10110101",32086 => "11001110",32087 => "01101111",32088 => "00111000",32089 => "10100001",32090 => "10100011",32091 => "01010100",32092 => "00100100",32093 => "10100110",32094 => "01000010",32095 => "10011010",32096 => "10001101",32097 => "10111000",32098 => "10011101",32099 => "10101001",32100 => "11011010",32101 => "10010110",32102 => "00010000",32103 => "10010100",32104 => "10101100",32105 => "00001100",32106 => "10001011",32107 => "10110000",32108 => "10101100",32109 => "01110000",32110 => "11010000",32111 => "10101111",32112 => "11010000",32113 => "00110000",32114 => "00011100",32115 => "00111000",32116 => "10010101",32117 => "01010111",32118 => "00111110",32119 => "10110101",32120 => "01110001",32121 => "00110110",32122 => "10000101",32123 => "01001101",32124 => "10010010",32125 => "11111010",32126 => "01010101",32127 => "00101001",32128 => "10001111",32129 => "10111110",32130 => "01011101",32131 => "10110010",32132 => "10110100",32133 => "01011101",32134 => "00101101",32135 => "00001100",32136 => "01001100",32137 => "11110110",32138 => "00001000",32139 => "00001100",32140 => "11000100",32141 => "00001000",32142 => "11111111",32143 => "01100001",32144 => "00011100",32145 => "11011011",32146 => "01111000",32147 => "11101000",32148 => "10101001",32149 => "11100101",32150 => "11010111",32151 => "01011010",32152 => "00010101",32153 => "01011100",32154 => "01100111",32155 => "00011001",32156 => "10100001",32157 => "10100110",32158 => "11110001",32159 => "10101111",32160 => "10101011",32161 => "01101111",32162 => "00111011",32163 => "01000011",32164 => "11110010",32165 => "10101100",32166 => "11001101",32167 => "11111100",32168 => "10001100",32169 => "01001111",32170 => "00001111",32171 => "11011010",32172 => "10011010",32173 => "10010011",32174 => "11110101",32175 => "01011111",32176 => "01110110",32177 => "10111011",32178 => "10011110",32179 => "10010000",32180 => "01001100",32181 => "11011100",32182 => "10101010",32183 => "10001011",32184 => "11010110",32185 => "01101111",32186 => "11011110",32187 => "00010110",32188 => "01011000",32189 => "01110010",32190 => "10010101",32191 => "00011111",32192 => "01111011",32193 => "10110100",32194 => "11000001",32195 => "11110110",32196 => "11110010",32197 => "01110001",32198 => "01010101",32199 => "01010011",32200 => "11101010",32201 => "10001111",32202 => "00000101",32203 => "10110011",32204 => "11000101",32205 => "00100000",32206 => "01001110",32207 => "01100001",32208 => "11101011",32209 => "11110110",32210 => "11101101",32211 => "01001000",32212 => "01111001",32213 => "01110001",32214 => "10101100",32215 => "11010100",32216 => "00101010",32217 => "01101111",32218 => "00010001",32219 => "11111101",32220 => "00010000",32221 => "00111011",32222 => "01110100",32223 => "10101001",32224 => "11010011",32225 => "10011101",32226 => "01001010",32227 => "01001110",32228 => "10100010",32229 => "10101101",32230 => "10111011",32231 => "11111001",32232 => "10000100",32233 => "00101010",32234 => "00100001",32235 => "11000111",32236 => "11101111",32237 => "01111000",32238 => "00100101",32239 => "01100101",32240 => "10110010",32241 => "00001100",32242 => "01101011",32243 => "10100001",32244 => "11100001",32245 => "00110000",32246 => "10110100",32247 => "01101001",32248 => "00000100",32249 => "00110001",32250 => "01000100",32251 => "01101000",32252 => "01011100",32253 => "01000001",32254 => "00011000",32255 => "10010001",32256 => "01011111",32257 => "00111000",32258 => "11010101",32259 => "11100000",32260 => "00011100",32261 => "00111010",32262 => "01111000",32263 => "00101100",32264 => "00000000",32265 => "11001011",32266 => "00000110",32267 => "01101111",32268 => "11011101",32269 => "10011101",32270 => "11000011",32271 => "01101100",32272 => "01001101",32273 => "11011110",32274 => "00111100",32275 => "01100000",32276 => "00011001",32277 => "11011011",32278 => "11010111",32279 => "01101001",32280 => "00000100",32281 => "10010011",32282 => "00010111",32283 => "11010110",32284 => "10110010",32285 => "01111001",32286 => "01001010",32287 => "01010010",32288 => "11010111",32289 => "00100011",32290 => "10000001",32291 => "10001001",32292 => "11011101",32293 => "11001010",32294 => "11100110",32295 => "00001001",32296 => "00000000",32297 => "01100000",32298 => "10101010",32299 => "11000110",32300 => "01010111",32301 => "00110100",32302 => "01100100",32303 => "00101110",32304 => "10001010",32305 => "00001010",32306 => "11101100",32307 => "01101100",32308 => "11000111",32309 => "00100001",32310 => "00111000",32311 => "01001010",32312 => "01101110",32313 => "01000000",32314 => "11110011",32315 => "01100000",32316 => "10011111",32317 => "10110101",32318 => "00110111",32319 => "01111010",32320 => "10100111",32321 => "11101000",32322 => "11001101",32323 => "00011111",32324 => "00110000",32325 => "00100111",32326 => "01100111",32327 => "10101011",32328 => "00100001",32329 => "00010100",32330 => "10100101",32331 => "10000010",32332 => "01010111",32333 => "00111111",32334 => "00111100",32335 => "11111110",32336 => "10010100",32337 => "11000011",32338 => "00111011",32339 => "00100101",32340 => "01010100",32341 => "01110110",32342 => "11110000",32343 => "00110011",32344 => "10001100",32345 => "01100000",32346 => "10000001",32347 => "10000001",32348 => "00110001",32349 => "00111011",32350 => "01111010",32351 => "01111111",32352 => "10010100",32353 => "10010010",32354 => "01011010",32355 => "01000011",32356 => "11011001",32357 => "00001101",32358 => "00001110",32359 => "00100010",32360 => "01110110",32361 => "11000111",32362 => "11110101",32363 => "10001111",32364 => "10010111",32365 => "11011011",32366 => "11100001",32367 => "11011011",32368 => "10000001",32369 => "00110101",32370 => "01001000",32371 => "10001110",32372 => "01111011",32373 => "11000110",32374 => "01001010",32375 => "00101001",32376 => "01111100",32377 => "00110110",32378 => "10000010",32379 => "11010111",32380 => "10110000",32381 => "01011101",32382 => "01001101",32383 => "01101000",32384 => "11110011",32385 => "11110101",32386 => "11110111",32387 => "00010011",32388 => "01100011",32389 => "11101011",32390 => "10011111",32391 => "10000101",32392 => "11011001",32393 => "00101010",32394 => "10110100",32395 => "11010001",32396 => "11101110",32397 => "01000010",32398 => "10001100",32399 => "10010101",32400 => "00110100",32401 => "10100011",32402 => "00011000",32403 => "01111100",32404 => "01001100",32405 => "11011011",32406 => "10101100",32407 => "10100010",32408 => "01010111",32409 => "11111010",32410 => "01100110",32411 => "11111101",32412 => "00011110",32413 => "10001000",32414 => "00011001",32415 => "01110000",32416 => "11011010",32417 => "01011010",32418 => "01101111",32419 => "10001011",32420 => "01011001",32421 => "10011101",32422 => "10000001",32423 => "01011101",32424 => "00000011",32425 => "10011111",32426 => "10101000",32427 => "10000101",32428 => "00011110",32429 => "00100110",32430 => "10101100",32431 => "11101011",32432 => "00000000",32433 => "01111001",32434 => "10111000",32435 => "00010101",32436 => "00000001",32437 => "10110101",32438 => "00000111",32439 => "00000100",32440 => "00101110",32441 => "11110100",32442 => "01111111",32443 => "10011111",32444 => "01011011",32445 => "01011111",32446 => "11000001",32447 => "11100000",32448 => "10011010",32449 => "11111000",32450 => "00100000",32451 => "00111110",32452 => "01000011",32453 => "11100101",32454 => "11010100",32455 => "00111000",32456 => "01101001",32457 => "01010001",32458 => "00011010",32459 => "10000101",32460 => "01010000",32461 => "01110000",32462 => "11110110",32463 => "01011100",32464 => "01011100",32465 => "10111001",32466 => "10101001",32467 => "01010000",32468 => "00111001",32469 => "11001000",32470 => "00010111",32471 => "11111011",32472 => "11001101",32473 => "01110100",32474 => "11100110",32475 => "11100101",32476 => "00001110",32477 => "00111001",32478 => "10100111",32479 => "01000000",32480 => "01100000",32481 => "10101111",32482 => "10001111",32483 => "00001001",32484 => "01001011",32485 => "00000011",32486 => "00111101",32487 => "00011001",32488 => "11101100",32489 => "00101111",32490 => "01011110",32491 => "10110100",32492 => "11110011",32493 => "10010010",32494 => "01101010",32495 => "00010100",32496 => "01101011",32497 => "10011111",32498 => "01001101",32499 => "10111101",32500 => "11001111",32501 => "11001000",32502 => "10111011",32503 => "10011011",32504 => "11101010",32505 => "10011101",32506 => "00001011",32507 => "10000011",32508 => "10110011",32509 => "10000100",32510 => "10011000",32511 => "10110010",32512 => "00101001",32513 => "01010000",32514 => "11100011",32515 => "11000010",32516 => "11001010",32517 => "10010000",32518 => "01100111",32519 => "11100111",32520 => "10111110",32521 => "00100000",32522 => "01000001",32523 => "01011110",32524 => "01010000",32525 => "01101011",32526 => "11000011",32527 => "00111100",32528 => "01001111",32529 => "00000100",32530 => "10100101",32531 => "11100011",32532 => "00011001",32533 => "11000001",32534 => "10000001",32535 => "01101011",32536 => "00010101",32537 => "11010111",32538 => "00000001",32539 => "10111110",32540 => "01110010",32541 => "01100110",32542 => "10101100",32543 => "01110100",32544 => "11010011",32545 => "10100111",32546 => "00010100",32547 => "01011011",32548 => "00001010",32549 => "00010100",32550 => "01110011",32551 => "01101111",32552 => "00110101",32553 => "01000011",32554 => "00100101",32555 => "00100100",32556 => "11111011",32557 => "10010110",32558 => "00101111",32559 => "01100001",32560 => "10010111",32561 => "11100000",32562 => "00001100",32563 => "00110100",32564 => "00111111",32565 => "00111101",32566 => "01111001",32567 => "00100010",32568 => "11001101",32569 => "00110110",32570 => "10000110",32571 => "01110111",32572 => "00010011",32573 => "10001001",32574 => "01101110",32575 => "10111001",32576 => "01001001",32577 => "01000101",32578 => "00010001",32579 => "10110100",32580 => "10011100",32581 => "00101011",32582 => "10101011",32583 => "00010011",32584 => "11011011",32585 => "10001001",32586 => "01000101",32587 => "00100111",32588 => "01000011",32589 => "00001001",32590 => "11011010",32591 => "11101100",32592 => "01100110",32593 => "00101101",32594 => "01101110",32595 => "01111110",32596 => "01010100",32597 => "11111110",32598 => "10001001",32599 => "11010100",32600 => "01001001",32601 => "01011000",32602 => "10010000",32603 => "01001000",32604 => "01110100",32605 => "01100100",32606 => "00010110",32607 => "00111111",32608 => "01000000",32609 => "00110000",32610 => "01110010",32611 => "11101001",32612 => "00000011",32613 => "10011001",32614 => "00000110",32615 => "11000110",32616 => "00000010",32617 => "01111110",32618 => "00010100",32619 => "01100010",32620 => "10010000",32621 => "01011000",32622 => "10001111",32623 => "00000100",32624 => "01000101",32625 => "00101110",32626 => "10010011",32627 => "10000100",32628 => "11110100",32629 => "11111011",32630 => "10011010",32631 => "01000000",32632 => "00001010",32633 => "01101110",32634 => "11001100",32635 => "01101011",32636 => "10100101",32637 => "10001111",32638 => "00001001",32639 => "01111001",32640 => "10010101",32641 => "01101100",32642 => "00000011",32643 => "01001110",32644 => "01101101",32645 => "01100000",32646 => "00100001",32647 => "10000011",32648 => "01000110",32649 => "01011101",32650 => "00111101",32651 => "01101100",32652 => "11011011",32653 => "11010111",32654 => "00111000",32655 => "00010001",32656 => "01110011",32657 => "11111010",32658 => "00011110",32659 => "01011100",32660 => "10101101",32661 => "01101100",32662 => "10000111",32663 => "00010010",32664 => "01000000",32665 => "01110010",32666 => "10011101",32667 => "00110110",32668 => "11100010",32669 => "01011000",32670 => "10010010",32671 => "11010000",32672 => "00111110",32673 => "00101101",32674 => "11010000",32675 => "00010110",32676 => "11011010",32677 => "01011101",32678 => "10110000",32679 => "01010111",32680 => "11001010",32681 => "00011011",32682 => "01011011",32683 => "10000001",32684 => "00001101",32685 => "11010000",32686 => "00010100",32687 => "00001000",32688 => "00100110",32689 => "00011010",32690 => "10000100",32691 => "00011010",32692 => "01000000",32693 => "01011100",32694 => "00000001",32695 => "00111111",32696 => "01011011",32697 => "00011100",32698 => "01010101",32699 => "00000011",32700 => "11000111",32701 => "11011111",32702 => "01011000",32703 => "11111110",32704 => "00101110",32705 => "01101111",32706 => "01110101",32707 => "01100100",32708 => "11000001",32709 => "10101011",32710 => "11101010",32711 => "00100010",32712 => "10110001",32713 => "01100101",32714 => "10101010",32715 => "10010001",32716 => "01110010",32717 => "01110111",32718 => "10110010",32719 => "10011111",32720 => "11111011",32721 => "01111110",32722 => "01000001",32723 => "11111000",32724 => "11011111",32725 => "11010000",32726 => "00101101",32727 => "10010110",32728 => "01001011",32729 => "01011011",32730 => "10101001",32731 => "11001011",32732 => "00111100",32733 => "11000001",32734 => "11111101",32735 => "00010011",32736 => "10110100",32737 => "00001010",32738 => "00010011",32739 => "01010010",32740 => "01101001",32741 => "01010100",32742 => "11111010",32743 => "10001101",32744 => "00011001",32745 => "00001101",32746 => "01001100",32747 => "10111000",32748 => "00101011",32749 => "10110101",32750 => "01001101",32751 => "00100110",32752 => "10010001",32753 => "01110010",32754 => "11000111",32755 => "10100110",32756 => "10110010",32757 => "00001010",32758 => "00010000",32759 => "01000001",32760 => "01000011",32761 => "11100001",32762 => "11101101",32763 => "00101111",32764 => "00111110",32765 => "01110111",32766 => "11001001",32767 => "10110011",32768 => "00100100",32769 => "11011000",32770 => "10010011",32771 => "10010101",32772 => "11100000",32773 => "01100111",32774 => "01110111",32775 => "01001100",32776 => "00001100",32777 => "01001011",32778 => "00111010",32779 => "10100000",32780 => "10101001",32781 => "11001100",32782 => "10011011",32783 => "11110110",32784 => "01010000",32785 => "11100100",32786 => "01010100",32787 => "00011001",32788 => "11101011",32789 => "00100011",32790 => "00101011",32791 => "11011101",32792 => "00011001",32793 => "11000011",32794 => "01110011",32795 => "11000011",32796 => "00011100",32797 => "00111011",32798 => "11000111",32799 => "10011011",32800 => "10111000",32801 => "10010101",32802 => "11000000",32803 => "01010010",32804 => "10110111",32805 => "01111001",32806 => "10100010",32807 => "01000111",32808 => "00001110",32809 => "10011110",32810 => "00110011",32811 => "00001110",32812 => "01001000",32813 => "00010001",32814 => "11100000",32815 => "00010111",32816 => "01001011",32817 => "11110100",32818 => "10110010",32819 => "10010001",32820 => "01111000",32821 => "11100110",32822 => "01111101",32823 => "10000000",32824 => "01010000",32825 => "11011111",32826 => "00001110",32827 => "01011100",32828 => "00100110",32829 => "00000100",32830 => "01110000",32831 => "10100001",32832 => "01111101",32833 => "10000000",32834 => "01111110",32835 => "00011100",32836 => "00100110",32837 => "01101110",32838 => "11111001",32839 => "11101010",32840 => "11010000",32841 => "10101101",32842 => "11110100",32843 => "11000000",32844 => "11001111",32845 => "01110100",32846 => "10010011",32847 => "11011100",32848 => "01001000",32849 => "01100001",32850 => "10011011",32851 => "01101001",32852 => "10000010",32853 => "10100011",32854 => "00110010",32855 => "10110011",32856 => "10000011",32857 => "00011100",32858 => "11010110",32859 => "00000101",32860 => "01010001",32861 => "01001110",32862 => "00010111",32863 => "11011101",32864 => "00001001",32865 => "10010101",32866 => "00111010",32867 => "01111010",32868 => "01111100",32869 => "01111000",32870 => "10011110",32871 => "10110001",32872 => "11111101",32873 => "00111010",32874 => "11100000",32875 => "00011100",32876 => "00101010",32877 => "01000100",32878 => "01111100",32879 => "10000011",32880 => "01111101",32881 => "11000011",32882 => "01111111",32883 => "00100110",32884 => "01011010",32885 => "01001011",32886 => "11001000",32887 => "10011011",32888 => "01001110",32889 => "10000011",32890 => "00111010",32891 => "11101100",32892 => "11000001",32893 => "00100110",32894 => "11100101",32895 => "00100101",32896 => "00001101",32897 => "01000101",32898 => "01110100",32899 => "00100101",32900 => "01110100",32901 => "11100011",32902 => "11101010",32903 => "11010010",32904 => "11110110",32905 => "01110101",32906 => "10111000",32907 => "10010110",32908 => "11010010",32909 => "00001010",32910 => "00111100",32911 => "11100010",32912 => "11100010",32913 => "01110111",32914 => "11011111",32915 => "01111111",32916 => "10011110",32917 => "00101111",32918 => "10111111",32919 => "11001100",32920 => "00100110",32921 => "00100010",32922 => "10000000",32923 => "00000011",32924 => "01001011",32925 => "00001001",32926 => "00100001",32927 => "01100101",32928 => "11111001",32929 => "10101111",32930 => "00001000",32931 => "00110011",32932 => "01110010",32933 => "00011100",32934 => "01010110",32935 => "00111100",32936 => "10011101",32937 => "01110100",32938 => "00010111",32939 => "11100101",32940 => "00110110",32941 => "11101110",32942 => "01100110",32943 => "10101100",32944 => "10100000",32945 => "10101010",32946 => "00110000",32947 => "00001101",32948 => "00011011",32949 => "01010111",32950 => "00101000",32951 => "11000111",32952 => "00101101",32953 => "01010110",32954 => "00110110",32955 => "11001101",32956 => "11111110",32957 => "10101001",32958 => "11111111",32959 => "10100000",32960 => "11010011",32961 => "10101001",32962 => "01001000",32963 => "01010100",32964 => "10110110",32965 => "01110101",32966 => "11011011",32967 => "01111101",32968 => "01100101",32969 => "10000000",32970 => "00111100",32971 => "01011011",32972 => "10101111",32973 => "01110010",32974 => "01110111",32975 => "01000011",32976 => "00101010",32977 => "11101000",32978 => "01110000",32979 => "11101001",32980 => "00100000",32981 => "11101111",32982 => "01101100",32983 => "00110111",32984 => "01111001",32985 => "11001110",32986 => "10111011",32987 => "01001110",32988 => "00101011",32989 => "00010100",32990 => "11111001",32991 => "10010011",32992 => "10011010",32993 => "11100101",32994 => "10100011",32995 => "01010000",32996 => "10111010",32997 => "11000110",32998 => "01000101",32999 => "10101010",33000 => "00011001",33001 => "11111101",33002 => "11010001",33003 => "01100011",33004 => "10000001",33005 => "01101101",33006 => "10100110",33007 => "10010001",33008 => "10110110",33009 => "00010110",33010 => "00000011",33011 => "00110000",33012 => "00011100",33013 => "01100010",33014 => "11001110",33015 => "11000100",33016 => "01110110",33017 => "11000110",33018 => "10100110",33019 => "01110011",33020 => "10001010",33021 => "11110010",33022 => "10100111",33023 => "10100110",33024 => "10001100",33025 => "11110000",33026 => "11001001",33027 => "11000101",33028 => "11101001",33029 => "11000001",33030 => "11001010",33031 => "01101111",33032 => "01010000",33033 => "01110100",33034 => "00000101",33035 => "11100010",33036 => "10100110",33037 => "01000110",33038 => "00000100",33039 => "01111110",33040 => "01101101",33041 => "01010010",33042 => "11110001",33043 => "00001001",33044 => "00010000",33045 => "10011010",33046 => "01101010",33047 => "10101001",33048 => "11101111",33049 => "10110111",33050 => "01011111",33051 => "00011000",33052 => "10100010",33053 => "01101110",33054 => "10010100",33055 => "01011100",33056 => "01111100",33057 => "00101010",33058 => "10101100",33059 => "10100001",33060 => "10100011",33061 => "10100001",33062 => "10000000",33063 => "00010110",33064 => "10000101",33065 => "10111001",33066 => "10111000",33067 => "11111111",33068 => "00101111",33069 => "10000000",33070 => "11000011",33071 => "11000111",33072 => "11111010",33073 => "10001011",33074 => "11001110",33075 => "11111001",33076 => "10101101",33077 => "11110001",33078 => "01001100",33079 => "11000110",33080 => "00111011",33081 => "11001011",33082 => "01011011",33083 => "10011011",33084 => "10000101",33085 => "11110100",33086 => "11011000",33087 => "11011110",33088 => "10010110",33089 => "10011100",33090 => "11001111",33091 => "00000110",33092 => "00101110",33093 => "01010010",33094 => "11101011",33095 => "00100001",33096 => "00100000",33097 => "10110111",33098 => "11110111",33099 => "01100011",33100 => "11010111",33101 => "10001101",33102 => "10010010",33103 => "11110101",33104 => "11111010",33105 => "01100101",33106 => "11110110",33107 => "01011101",33108 => "00111101",33109 => "01001101",33110 => "10001000",33111 => "01110010",33112 => "10001101",33113 => "00100101",33114 => "10000010",33115 => "11010111",33116 => "10010000",33117 => "01000100",33118 => "11000110",33119 => "11010011",33120 => "01000110",33121 => "10000011",33122 => "10011010",33123 => "00010010",33124 => "00010100",33125 => "10101110",33126 => "10111010",33127 => "11010010",33128 => "11011010",33129 => "01101011",33130 => "10101010",33131 => "10000111",33132 => "10011000",33133 => "01011011",33134 => "10101100",33135 => "00011011",33136 => "11010000",33137 => "00000010",33138 => "10010000",33139 => "11101111",33140 => "11011100",33141 => "11001111",33142 => "00101010",33143 => "00000111",33144 => "11010100",33145 => "11011100",33146 => "11001000",33147 => "00100011",33148 => "10001011",33149 => "01101010",33150 => "10001101",33151 => "01010000",33152 => "00010111",33153 => "10111110",33154 => "11010110",33155 => "01101100",33156 => "01000001",33157 => "10100110",33158 => "11010100",33159 => "11001001",33160 => "10010111",33161 => "00110010",33162 => "00000101",33163 => "11011011",33164 => "00100100",33165 => "11101001",33166 => "11101101",33167 => "11110011",33168 => "10000011",33169 => "01001111",33170 => "10100011",33171 => "01010110",33172 => "01001111",33173 => "10010011",33174 => "00110110",33175 => "11010100",33176 => "11010101",33177 => "11111000",33178 => "11011100",33179 => "10111111",33180 => "00111110",33181 => "01101110",33182 => "01010001",33183 => "10110101",33184 => "10011011",33185 => "10001010",33186 => "00001110",33187 => "01010001",33188 => "11101110",33189 => "01011010",33190 => "00011100",33191 => "11101111",33192 => "01110011",33193 => "11010111",33194 => "11011100",33195 => "01100010",33196 => "01100000",33197 => "01000000",33198 => "11101100",33199 => "00001001",33200 => "01110010",33201 => "00111000",33202 => "11111111",33203 => "00010110",33204 => "01101011",33205 => "11000101",33206 => "10011101",33207 => "01000110",33208 => "11100001",33209 => "00110001",33210 => "00001101",33211 => "00011001",33212 => "10101001",33213 => "01010101",33214 => "00110000",33215 => "11010001",33216 => "00110001",33217 => "11000011",33218 => "01001110",33219 => "00111101",33220 => "11101101",33221 => "00000101",33222 => "01111111",33223 => "00010111",33224 => "10101101",33225 => "10110001",33226 => "01001110",33227 => "10010100",33228 => "01010110",33229 => "00000101",33230 => "10011000",33231 => "11010001",33232 => "10100111",33233 => "01010000",33234 => "00100010",33235 => "00100101",33236 => "11010001",33237 => "01010110",33238 => "01010110",33239 => "01001101",33240 => "01011001",33241 => "00100001",33242 => "00111101",33243 => "10100100",33244 => "11001000",33245 => "11111000",33246 => "11011111",33247 => "10100100",33248 => "00010011",33249 => "01001011",33250 => "00111101",33251 => "11110000",33252 => "00010100",33253 => "10110100",33254 => "11110111",33255 => "10110100",33256 => "01101000",33257 => "01110001",33258 => "00101010",33259 => "10111010",33260 => "11011100",33261 => "00000001",33262 => "01000010",33263 => "01000111",33264 => "10000111",33265 => "11011011",33266 => "01010111",33267 => "01110010",33268 => "10001011",33269 => "01111000",33270 => "00110110",33271 => "11011001",33272 => "00001011",33273 => "00001101",33274 => "01001100",33275 => "00000110",33276 => "10001000",33277 => "01011000",33278 => "10110101",33279 => "01000001",33280 => "10011011",33281 => "10001000",33282 => "10011001",33283 => "11110010",33284 => "00010101",33285 => "01101100",33286 => "10000010",33287 => "10000101",33288 => "10111001",33289 => "11010110",33290 => "00011001",33291 => "01010101",33292 => "01100001",33293 => "11100011",33294 => "01110111",33295 => "01101011",33296 => "00011000",33297 => "10111101",33298 => "10100110",33299 => "11001011",33300 => "11000110",33301 => "01010010",33302 => "11011100",33303 => "01110000",33304 => "10011101",33305 => "01011100",33306 => "00101110",33307 => "11100010",33308 => "01100110",33309 => "10010111",33310 => "11001101",33311 => "10101010",33312 => "01000010",33313 => "11100000",33314 => "11001110",33315 => "00111100",33316 => "10111110",33317 => "00011111",33318 => "01000110",33319 => "10111110",33320 => "00011110",33321 => "10100010",33322 => "11101111",33323 => "01110000",33324 => "11011010",33325 => "00011011",33326 => "10011011",33327 => "00001100",33328 => "11000111",33329 => "00001011",33330 => "10000001",33331 => "00100001",33332 => "10000111",33333 => "01100010",33334 => "11010110",33335 => "11110001",33336 => "01001001",33337 => "01011111",33338 => "01010100",33339 => "01010011",33340 => "10111011",33341 => "11110011",33342 => "01101111",33343 => "10011000",33344 => "11100110",33345 => "11011110",33346 => "01000101",33347 => "01101000",33348 => "01000111",33349 => "11011011",33350 => "00101001",33351 => "10100001",33352 => "01101011",33353 => "00110011",33354 => "00110001",33355 => "10110101",33356 => "00011010",33357 => "01001001",33358 => "11001110",33359 => "01001001",33360 => "00100101",33361 => "11011010",33362 => "01110111",33363 => "00000101",33364 => "01000100",33365 => "00110101",33366 => "01010110",33367 => "10111111",33368 => "10001011",33369 => "11111100",33370 => "10010100",33371 => "10001110",33372 => "10001111",33373 => "11100111",33374 => "11000101",33375 => "10010101",33376 => "01100100",33377 => "10000101",33378 => "01011110",33379 => "00010000",33380 => "11001000",33381 => "11110000",33382 => "01101110",33383 => "00111000",33384 => "10111101",33385 => "00111110",33386 => "01110110",33387 => "01000100",33388 => "00000100",33389 => "11000000",33390 => "01100001",33391 => "00100000",33392 => "10110111",33393 => "10101101",33394 => "01110000",33395 => "01101101",33396 => "10001100",33397 => "00101010",33398 => "10010010",33399 => "10110011",33400 => "01001000",33401 => "01111001",33402 => "01011010",33403 => "01111000",33404 => "11000110",33405 => "00101011",33406 => "00001011",33407 => "00101110",33408 => "01001100",33409 => "00110010",33410 => "00011100",33411 => "10100100",33412 => "11011001",33413 => "00000110",33414 => "11101000",33415 => "00011101",33416 => "00001111",33417 => "10110111",33418 => "10101010",33419 => "00101110",33420 => "00101100",33421 => "01111101",33422 => "00010110",33423 => "00000011",33424 => "10011000",33425 => "00110000",33426 => "11011100",33427 => "11010111",33428 => "11101111",33429 => "01000010",33430 => "00011101",33431 => "00010110",33432 => "00001111",33433 => "11000000",33434 => "00110101",33435 => "01000110",33436 => "10110000",33437 => "10001000",33438 => "00101001",33439 => "11001101",33440 => "10000001",33441 => "11111001",33442 => "01110110",33443 => "10100010",33444 => "00110011",33445 => "10001110",33446 => "10110111",33447 => "10111011",33448 => "01100100",33449 => "11010010",33450 => "11011001",33451 => "11101001",33452 => "11111000",33453 => "00111101",33454 => "10000001",33455 => "11001110",33456 => "00100010",33457 => "10100010",33458 => "00110100",33459 => "00111001",33460 => "11011011",33461 => "11001110",33462 => "00110001",33463 => "01000011",33464 => "10100010",33465 => "00101101",33466 => "00011011",33467 => "11111101",33468 => "10010110",33469 => "01110000",33470 => "00001001",33471 => "01010000",33472 => "10110001",33473 => "11001100",33474 => "11111011",33475 => "11100100",33476 => "00100010",33477 => "10000010",33478 => "11001001",33479 => "01011011",33480 => "00100100",33481 => "01100011",33482 => "01001001",33483 => "01010111",33484 => "01000001",33485 => "11110101",33486 => "10001001",33487 => "01000001",33488 => "11110101",33489 => "11101011",33490 => "01001100",33491 => "10110010",33492 => "11011111",33493 => "01000001",33494 => "10010000",33495 => "10011001",33496 => "10000011",33497 => "11001100",33498 => "11101001",33499 => "01110101",33500 => "01001110",33501 => "00010000",33502 => "11111011",33503 => "10101011",33504 => "10001110",33505 => "11000011",33506 => "11010001",33507 => "11100101",33508 => "10011000",33509 => "11111000",33510 => "01111100",33511 => "01100011",33512 => "00101010",33513 => "11111000",33514 => "00000111",33515 => "00010111",33516 => "01100100",33517 => "10000000",33518 => "11110010",33519 => "11000111",33520 => "10110110",33521 => "11010001",33522 => "11101000",33523 => "01000100",33524 => "01111111",33525 => "00100100",33526 => "11101010",33527 => "01111101",33528 => "01001110",33529 => "00010110",33530 => "00100100",33531 => "01100001",33532 => "10010011",33533 => "11001101",33534 => "00100110",33535 => "01011001",33536 => "00110110",33537 => "11110001",33538 => "11001101",33539 => "00100111",33540 => "00011111",33541 => "11001001",33542 => "01100000",33543 => "01110101",33544 => "00110111",33545 => "11110001",33546 => "11000101",33547 => "00100101",33548 => "11100011",33549 => "00110111",33550 => "00010100",33551 => "00000110",33552 => "01111100",33553 => "10010000",33554 => "10011001",33555 => "11011001",33556 => "11011000",33557 => "10011101",33558 => "11111010",33559 => "10110010",33560 => "01111001",33561 => "10101010",33562 => "01000111",33563 => "11011110",33564 => "11001010",33565 => "10000110",33566 => "01011000",33567 => "00100001",33568 => "00110011",33569 => "00100101",33570 => "00101111",33571 => "00001011",33572 => "01110111",33573 => "11111000",33574 => "11000001",33575 => "10100001",33576 => "11101010",33577 => "10101110",33578 => "01010010",33579 => "00111101",33580 => "01011010",33581 => "01110011",33582 => "10000111",33583 => "00101100",33584 => "11100001",33585 => "11100001",33586 => "11011101",33587 => "00100101",33588 => "10000110",33589 => "00110111",33590 => "10110110",33591 => "11010001",33592 => "10101000",33593 => "10000101",33594 => "01110001",33595 => "11011010",33596 => "11101101",33597 => "00110010",33598 => "01000000",33599 => "10000111",33600 => "11001111",33601 => "01100010",33602 => "01101000",33603 => "11111011",33604 => "00001110",33605 => "11011001",33606 => "00001110",33607 => "00101110",33608 => "01000010",33609 => "01001000",33610 => "11011101",33611 => "10001110",33612 => "10101010",33613 => "11110100",33614 => "00110011",33615 => "01110011",33616 => "10101011",33617 => "11101110",33618 => "00001010",33619 => "11011111",33620 => "11000100",33621 => "10100000",33622 => "10010111",33623 => "11010101",33624 => "11000011",33625 => "01100111",33626 => "01111011",33627 => "10110101",33628 => "01110000",33629 => "00010110",33630 => "00000000",33631 => "10001010",33632 => "01100001",33633 => "10100000",33634 => "11110100",33635 => "00100000",33636 => "00011100",33637 => "10100011",33638 => "01001010",33639 => "01111111",33640 => "10000101",33641 => "10100000",33642 => "00101101",33643 => "10110110",33644 => "11011011",33645 => "11001000",33646 => "10010100",33647 => "11001011",33648 => "01100011",33649 => "01111010",33650 => "01011111",33651 => "00000001",33652 => "00110011",33653 => "11010101",33654 => "10111101",33655 => "10011111",33656 => "11001100",33657 => "11011000",33658 => "11000001",33659 => "00101101",33660 => "01000100",33661 => "01100100",33662 => "11001101",33663 => "11001100",33664 => "01000111",33665 => "01010111",33666 => "01011111",33667 => "10001010",33668 => "00110101",33669 => "00100101",33670 => "10001111",33671 => "10110111",33672 => "11110011",33673 => "10010010",33674 => "10001001",33675 => "01111011",33676 => "01111010",33677 => "01100101",33678 => "11010110",33679 => "00110000",33680 => "01111101",33681 => "11011101",33682 => "01101111",33683 => "10101001",33684 => "00110110",33685 => "01010101",33686 => "11011110",33687 => "11100101",33688 => "10101011",33689 => "11111000",33690 => "10000010",33691 => "11000000",33692 => "01110111",33693 => "11001010",33694 => "01001010",33695 => "10000101",33696 => "11011101",33697 => "00110110",33698 => "11100110",33699 => "10000100",33700 => "10111000",33701 => "00110010",33702 => "01010111",33703 => "11000000",33704 => "10111000",33705 => "01000011",33706 => "01001011",33707 => "10111001",33708 => "10111000",33709 => "00110101",33710 => "01111111",33711 => "00010101",33712 => "11010000",33713 => "00101011",33714 => "11010010",33715 => "01000000",33716 => "10011001",33717 => "10110110",33718 => "01101111",33719 => "01001000",33720 => "10110010",33721 => "01111000",33722 => "00101010",33723 => "01110101",33724 => "11100111",33725 => "01011111",33726 => "01110100",33727 => "01101011",33728 => "00100100",33729 => "10011100",33730 => "00010111",33731 => "11010110",33732 => "10010101",33733 => "11010111",33734 => "10100000",33735 => "00011111",33736 => "01000001",33737 => "01111011",33738 => "11001101",33739 => "01011100",33740 => "00111010",33741 => "00000110",33742 => "01110000",33743 => "10101110",33744 => "01010011",33745 => "01010000",33746 => "11100111",33747 => "00010110",33748 => "10000110",33749 => "00111100",33750 => "00001010",33751 => "00000110",33752 => "11101101",33753 => "10000110",33754 => "00000010",33755 => "10101100",33756 => "00111111",33757 => "01000010",33758 => "10011101",33759 => "10111001",33760 => "01111001",33761 => "10011101",33762 => "10010000",33763 => "11100100",33764 => "11110100",33765 => "00111110",33766 => "10011100",33767 => "11100010",33768 => "00011011",33769 => "10000001",33770 => "11100011",33771 => "10111101",33772 => "01111110",33773 => "01001011",33774 => "10100111",33775 => "11000111",33776 => "00000101",33777 => "00101000",33778 => "01011101",33779 => "11101110",33780 => "11011000",33781 => "00110001",33782 => "01001100",33783 => "10110011",33784 => "10110001",33785 => "10000000",33786 => "00000101",33787 => "00001100",33788 => "11000000",33789 => "10000010",33790 => "00000010",33791 => "10011110",33792 => "10011101",33793 => "10000100",33794 => "10001010",33795 => "00110011",33796 => "11110010",33797 => "01100110",33798 => "00110011",33799 => "01101011",33800 => "01110001",33801 => "00110010",33802 => "11101110",33803 => "10000101",33804 => "11010001",33805 => "11100110",33806 => "01001000",33807 => "01000000",33808 => "01010011",33809 => "00111000",33810 => "00000111",33811 => "01101011",33812 => "01101100",33813 => "00000100",33814 => "10101001",33815 => "00001010",33816 => "00110011",33817 => "11111000",33818 => "11101110",33819 => "01110100",33820 => "00110011",33821 => "10101000",33822 => "11010000",33823 => "10110010",33824 => "11011111",33825 => "00101111",33826 => "00101010",33827 => "10000000",33828 => "10111111",33829 => "00101100",33830 => "10011100",33831 => "01011101",33832 => "01001101",33833 => "11000110",33834 => "00001111",33835 => "10110010",33836 => "10111110",33837 => "01001010",33838 => "00111001",33839 => "00010001",33840 => "10011000",33841 => "00111111",33842 => "10111001",33843 => "10100001",33844 => "01101111",33845 => "11001000",33846 => "10110100",33847 => "01100101",33848 => "10000001",33849 => "00000000",33850 => "01110010",33851 => "00001000",33852 => "10111101",33853 => "01001010",33854 => "00001111",33855 => "10100000",33856 => "00010111",33857 => "00101100",33858 => "11110100",33859 => "01010100",33860 => "00110001",33861 => "10101110",33862 => "00101101",33863 => "10101101",33864 => "11111010",33865 => "01111011",33866 => "01010000",33867 => "11011010",33868 => "01000101",33869 => "10111000",33870 => "11110000",33871 => "11010011",33872 => "01111111",33873 => "00101111",33874 => "10100000",33875 => "11111011",33876 => "10100111",33877 => "11111010",33878 => "10100000",33879 => "11010100",33880 => "00101010",33881 => "10101001",33882 => "01101100",33883 => "11110111",33884 => "10011001",33885 => "00000101",33886 => "11111110",33887 => "00101011",33888 => "01100110",33889 => "10101001",33890 => "01000001",33891 => "00001101",33892 => "01001011",33893 => "01101011",33894 => "11101111",33895 => "00100000",33896 => "10101001",33897 => "10110100",33898 => "11001010",33899 => "01000001",33900 => "00000001",33901 => "10001100",33902 => "11101111",33903 => "00101111",33904 => "01110110",33905 => "10001110",33906 => "00011110",33907 => "01001101",33908 => "11010001",33909 => "10111011",33910 => "11100110",33911 => "11010001",33912 => "10010101",33913 => "00010111",33914 => "00001000",33915 => "01111100",33916 => "00000000",33917 => "00001011",33918 => "01000000",33919 => "00110000",33920 => "00000111",33921 => "11001101",33922 => "00001111",33923 => "11101011",33924 => "10110100",33925 => "10000010",33926 => "01001011",33927 => "01010100",33928 => "00000101",33929 => "01110111",33930 => "00100001",33931 => "10010000",33932 => "11101101",33933 => "00001100",33934 => "00110101",33935 => "00011010",33936 => "00111011",33937 => "01000101",33938 => "01001110",33939 => "00011100",33940 => "01000011",33941 => "00100011",33942 => "10011010",33943 => "10011011",33944 => "11111010",33945 => "10110011",33946 => "00101111",33947 => "11101111",33948 => "01001110",33949 => "00011001",33950 => "00100011",33951 => "00011011",33952 => "00111111",33953 => "01000111",33954 => "11111100",33955 => "00010101",33956 => "01100010",33957 => "01101111",33958 => "10101110",33959 => "01101001",33960 => "00001001",33961 => "01110101",33962 => "01101011",33963 => "00001101",33964 => "11111110",33965 => "01011010",33966 => "01010100",33967 => "00101111",33968 => "11000111",33969 => "01001110",33970 => "10110000",33971 => "10101101",33972 => "00011010",33973 => "01100001",33974 => "11111110",33975 => "01110011",33976 => "01111110",33977 => "10101010",33978 => "10011110",33979 => "10111000",33980 => "00100001",33981 => "10101111",33982 => "10100110",33983 => "10111010",33984 => "00110000",33985 => "01100000",33986 => "01110011",33987 => "00100100",33988 => "11110100",33989 => "01000101",33990 => "10011101",33991 => "00011101",33992 => "10000001",33993 => "11110101",33994 => "00110110",33995 => "01100101",33996 => "00000011",33997 => "00111001",33998 => "10001000",33999 => "10110100",34000 => "11101000",34001 => "00010110",34002 => "00010101",34003 => "00100011",34004 => "11110010",34005 => "00001011",34006 => "00111011",34007 => "11010100",34008 => "00011011",34009 => "11110010",34010 => "00110011",34011 => "01110111",34012 => "11100110",34013 => "11100000",34014 => "10001111",34015 => "10100100",34016 => "11011010",34017 => "00100111",34018 => "10011001",34019 => "01011011",34020 => "10001100",34021 => "00010101",34022 => "00111100",34023 => "01011101",34024 => "10101010",34025 => "01001110",34026 => "11010001",34027 => "11100111",34028 => "01001110",34029 => "00011110",34030 => "10110000",34031 => "11011110",34032 => "11111001",34033 => "00100011",34034 => "11100100",34035 => "11101111",34036 => "01001000",34037 => "10110101",34038 => "11111010",34039 => "01101011",34040 => "01100101",34041 => "11011101",34042 => "01001101",34043 => "11011010",34044 => "00100000",34045 => "01010100",34046 => "11010011",34047 => "01011101",34048 => "01100110",34049 => "10010100",34050 => "01000110",34051 => "10110101",34052 => "10010001",34053 => "00100111",34054 => "01100101",34055 => "10010100",34056 => "01100111",34057 => "00101111",34058 => "00111011",34059 => "10100111",34060 => "01111011",34061 => "10111010",34062 => "01100100",34063 => "01011111",34064 => "11011101",34065 => "00011000",34066 => "11011110",34067 => "11100000",34068 => "00111010",34069 => "00001000",34070 => "11010010",34071 => "11100000",34072 => "10111010",34073 => "10001001",34074 => "00010000",34075 => "11110100",34076 => "00111011",34077 => "00001010",34078 => "00010110",34079 => "00000100",34080 => "10001100",34081 => "00100100",34082 => "01000110",34083 => "11001101",34084 => "10111110",34085 => "11001110",34086 => "01011110",34087 => "10100110",34088 => "11011110",34089 => "01111011",34090 => "11010101",34091 => "01001100",34092 => "10110110",34093 => "11001011",34094 => "00111100",34095 => "01001101",34096 => "01110000",34097 => "10011000",34098 => "01110000",34099 => "00010111",34100 => "11000101",34101 => "00110100",34102 => "11100010",34103 => "01010001",34104 => "00010001",34105 => "11011001",34106 => "01001010",34107 => "10100111",34108 => "10101100",34109 => "11000111",34110 => "01011011",34111 => "01011010",34112 => "01000101",34113 => "11010001",34114 => "01111000",34115 => "11011010",34116 => "01010010",34117 => "01001110",34118 => "00010010",34119 => "01100101",34120 => "01111100",34121 => "10110001",34122 => "01100110",34123 => "00001011",34124 => "01011001",34125 => "01000110",34126 => "00000001",34127 => "00100000",34128 => "00101011",34129 => "00110111",34130 => "00100001",34131 => "00110000",34132 => "00110110",34133 => "01110101",34134 => "10111011",34135 => "11100111",34136 => "10101000",34137 => "00011100",34138 => "10110001",34139 => "10101111",34140 => "11110001",34141 => "10010110",34142 => "11100111",34143 => "00001010",34144 => "10101010",34145 => "01111011",34146 => "01011000",34147 => "00101111",34148 => "11001011",34149 => "01000010",34150 => "10111000",34151 => "00100011",34152 => "00101111",34153 => "01111000",34154 => "10001100",34155 => "10101000",34156 => "01000101",34157 => "10111111",34158 => "00000110",34159 => "10111011",34160 => "00100010",34161 => "01111010",34162 => "10111100",34163 => "00111111",34164 => "00111100",34165 => "01001001",34166 => "11100011",34167 => "11001011",34168 => "10010110",34169 => "10111011",34170 => "11101001",34171 => "11011110",34172 => "01010111",34173 => "10100000",34174 => "00011101",34175 => "01100111",34176 => "00000101",34177 => "01000001",34178 => "00100111",34179 => "10101000",34180 => "10010101",34181 => "01001100",34182 => "00100000",34183 => "11110001",34184 => "01001111",34185 => "00100011",34186 => "10001110",34187 => "11110000",34188 => "01101001",34189 => "01000111",34190 => "10001011",34191 => "00010001",34192 => "10001010",34193 => "00100100",34194 => "00011110",34195 => "11000011",34196 => "10110100",34197 => "11001011",34198 => "01010010",34199 => "00100000",34200 => "00001010",34201 => "11010010",34202 => "10000011",34203 => "00001101",34204 => "01011110",34205 => "01101101",34206 => "00111010",34207 => "01100010",34208 => "11011101",34209 => "11111110",34210 => "11001100",34211 => "11100111",34212 => "00001111",34213 => "11011000",34214 => "01110111",34215 => "00100001",34216 => "01101011",34217 => "11010010",34218 => "11011011",34219 => "11010010",34220 => "01100000",34221 => "01111110",34222 => "11110111",34223 => "11101100",34224 => "01111111",34225 => "01000011",34226 => "10011111",34227 => "11100100",34228 => "01111110",34229 => "10110110",34230 => "11111011",34231 => "00010101",34232 => "11011010",34233 => "10100100",34234 => "10111010",34235 => "01101111",34236 => "00101000",34237 => "10001111",34238 => "11111100",34239 => "00010000",34240 => "11111110",34241 => "11111000",34242 => "00110000",34243 => "01101100",34244 => "11110101",34245 => "10101101",34246 => "01111010",34247 => "00001010",34248 => "10001000",34249 => "01011001",34250 => "00100011",34251 => "01000100",34252 => "00010001",34253 => "10110111",34254 => "11110010",34255 => "10001101",34256 => "01101101",34257 => "11000110",34258 => "11110011",34259 => "10000011",34260 => "10111100",34261 => "10000011",34262 => "01111001",34263 => "11100100",34264 => "00011000",34265 => "11110101",34266 => "11011010",34267 => "01001111",34268 => "10011100",34269 => "01101100",34270 => "01000000",34271 => "01100111",34272 => "01010100",34273 => "00010010",34274 => "11010111",34275 => "00011000",34276 => "10000111",34277 => "11001011",34278 => "11010111",34279 => "10100001",34280 => "10111110",34281 => "00000011",34282 => "10010111",34283 => "11001010",34284 => "01011111",34285 => "10010110",34286 => "00010110",34287 => "10011000",34288 => "10011000",34289 => "01101000",34290 => "10001000",34291 => "10111100",34292 => "10000010",34293 => "00000001",34294 => "11010100",34295 => "10011010",34296 => "10010101",34297 => "00011110",34298 => "10010111",34299 => "00110010",34300 => "00110010",34301 => "01011110",34302 => "10111110",34303 => "11010100",34304 => "11001000",34305 => "10011111",34306 => "01111111",34307 => "11111110",34308 => "10101110",34309 => "11011011",34310 => "11110110",34311 => "01001111",34312 => "00111101",34313 => "00001110",34314 => "01001111",34315 => "10101000",34316 => "11011101",34317 => "11011011",34318 => "10010110",34319 => "00010011",34320 => "10101110",34321 => "00110010",34322 => "01101010",34323 => "11010011",34324 => "10110100",34325 => "10111111",34326 => "10110011",34327 => "01101101",34328 => "01011000",34329 => "10000111",34330 => "01000000",34331 => "11100100",34332 => "00100010",34333 => "00010001",34334 => "00100010",34335 => "11101111",34336 => "10100001",34337 => "10111000",34338 => "01000000",34339 => "11010101",34340 => "10101110",34341 => "11111110",34342 => "00000010",34343 => "10011110",34344 => "10001110",34345 => "00111011",34346 => "00110100",34347 => "10111010",34348 => "01111110",34349 => "01010000",34350 => "10011100",34351 => "11100011",34352 => "00010101",34353 => "01000000",34354 => "00100001",34355 => "01001111",34356 => "10001100",34357 => "11101111",34358 => "00010010",34359 => "11010101",34360 => "10110010",34361 => "01111011",34362 => "00111001",34363 => "10001001",34364 => "00100110",34365 => "00000100",34366 => "11111111",34367 => "01011000",34368 => "11010101",34369 => "00100101",34370 => "01101011",34371 => "00100101",34372 => "10111101",34373 => "11100010",34374 => "11100111",34375 => "10111000",34376 => "01000001",34377 => "00101011",34378 => "11011100",34379 => "10101000",34380 => "11011000",34381 => "10010010",34382 => "10110011",34383 => "11101100",34384 => "11001000",34385 => "00001011",34386 => "01100010",34387 => "01101100",34388 => "10011111",34389 => "11110111",34390 => "00111010",34391 => "01011100",34392 => "11011011",34393 => "01001101",34394 => "10110010",34395 => "01111001",34396 => "10101010",34397 => "11010101",34398 => "00101000",34399 => "10110111",34400 => "00001111",34401 => "11010100",34402 => "00110000",34403 => "11011000",34404 => "10011001",34405 => "00011010",34406 => "01010000",34407 => "01010111",34408 => "01011110",34409 => "01000111",34410 => "01111110",34411 => "11101110",34412 => "10011001",34413 => "01101100",34414 => "01010110",34415 => "00000110",34416 => "01001001",34417 => "11100100",34418 => "00000010",34419 => "10100111",34420 => "11111000",34421 => "11111010",34422 => "10001101",34423 => "01001011",34424 => "01000110",34425 => "00010000",34426 => "01111100",34427 => "01001010",34428 => "10100101",34429 => "01000100",34430 => "01110111",34431 => "00001000",34432 => "10101001",34433 => "01111000",34434 => "10100101",34435 => "10010110",34436 => "00011010",34437 => "11000000",34438 => "11111000",34439 => "00000100",34440 => "01010110",34441 => "11110100",34442 => "01100001",34443 => "10100011",34444 => "10111111",34445 => "01111000",34446 => "11011111",34447 => "01001110",34448 => "10001000",34449 => "01101111",34450 => "01010001",34451 => "11110111",34452 => "10111010",34453 => "10000111",34454 => "11010111",34455 => "00111000",34456 => "01010100",34457 => "00101101",34458 => "10110001",34459 => "00100000",34460 => "01011100",34461 => "00011101",34462 => "10100100",34463 => "01010000",34464 => "00001001",34465 => "00101010",34466 => "01100011",34467 => "00110011",34468 => "10010001",34469 => "10000111",34470 => "00111101",34471 => "01000101",34472 => "00001100",34473 => "11111100",34474 => "00001111",34475 => "01001000",34476 => "10011000",34477 => "00010011",34478 => "11110110",34479 => "10000011",34480 => "00001000",34481 => "10100010",34482 => "00001111",34483 => "10111010",34484 => "11001001",34485 => "11100000",34486 => "10111011",34487 => "11000001",34488 => "10100110",34489 => "10111011",34490 => "00010000",34491 => "00101111",34492 => "01101110",34493 => "11001011",34494 => "01000111",34495 => "10011011",34496 => "11101001",34497 => "01110011",34498 => "00101100",34499 => "11101100",34500 => "11011100",34501 => "11001110",34502 => "10000001",34503 => "10000100",34504 => "00101010",34505 => "01110010",34506 => "10011110",34507 => "10110110",34508 => "11110011",34509 => "11000011",34510 => "01110101",34511 => "01010001",34512 => "10011010",34513 => "01110011",34514 => "00100001",34515 => "11110101",34516 => "11001111",34517 => "00101011",34518 => "01100000",34519 => "01010000",34520 => "11001101",34521 => "00001010",34522 => "00111001",34523 => "11011111",34524 => "00011001",34525 => "10100011",34526 => "11010101",34527 => "10110101",34528 => "11000111",34529 => "10100100",34530 => "10001011",34531 => "00101101",34532 => "11010010",34533 => "00011001",34534 => "10011101",34535 => "10101010",34536 => "00000000",34537 => "01111000",34538 => "11011100",34539 => "10000110",34540 => "00000100",34541 => "10000011",34542 => "01101011",34543 => "11101010",34544 => "01100000",34545 => "00001110",34546 => "11010111",34547 => "00011101",34548 => "00001101",34549 => "00000101",34550 => "01110011",34551 => "10100000",34552 => "10011011",34553 => "00010111",34554 => "11010100",34555 => "01100100",34556 => "01011100",34557 => "01010000",34558 => "00010110",34559 => "11000010",34560 => "00000011",34561 => "10001010",34562 => "10001011",34563 => "10111111",34564 => "10001100",34565 => "11011000",34566 => "00011000",34567 => "01101101",34568 => "00101011",34569 => "10110110",34570 => "11000000",34571 => "01111011",34572 => "10110011",34573 => "00001111",34574 => "11110110",34575 => "01000110",34576 => "01010111",34577 => "00010110",34578 => "11111000",34579 => "10011011",34580 => "11100001",34581 => "01111111",34582 => "10100001",34583 => "11000000",34584 => "00010001",34585 => "11010100",34586 => "01111010",34587 => "11010010",34588 => "01110110",34589 => "10101111",34590 => "00100101",34591 => "10010001",34592 => "11101011",34593 => "00111100",34594 => "01001111",34595 => "01011011",34596 => "01011101",34597 => "01110100",34598 => "11111000",34599 => "01110110",34600 => "10110000",34601 => "11110001",34602 => "11101001",34603 => "11111000",34604 => "10000110",34605 => "00010110",34606 => "11010001",34607 => "01001010",34608 => "01101001",34609 => "01111001",34610 => "11110101",34611 => "10011110",34612 => "00001110",34613 => "01110110",34614 => "10100101",34615 => "11000101",34616 => "00000110",34617 => "10111110",34618 => "01111000",34619 => "10100110",34620 => "10000101",34621 => "10100111",34622 => "11011110",34623 => "00001110",34624 => "10101110",34625 => "11011000",34626 => "00000011",34627 => "11111011",34628 => "00100000",34629 => "00000101",34630 => "00111010",34631 => "01011001",34632 => "00110100",34633 => "00111111",34634 => "11100001",34635 => "11101110",34636 => "01101100",34637 => "10111010",34638 => "00101000",34639 => "00000011",34640 => "11111100",34641 => "10100111",34642 => "10101000",34643 => "11101001",34644 => "11000001",34645 => "00111110",34646 => "11000000",34647 => "01101010",34648 => "01110100",34649 => "01101110",34650 => "11010111",34651 => "00010101",34652 => "10101110",34653 => "00100100",34654 => "10101100",34655 => "10010110",34656 => "11110101",34657 => "00111101",34658 => "00010111",34659 => "01110000",34660 => "01101100",34661 => "01111110",34662 => "11001010",34663 => "11000000",34664 => "00111011",34665 => "11110111",34666 => "11100101",34667 => "10011101",34668 => "01110100",34669 => "11011000",34670 => "10100000",34671 => "10101111",34672 => "11111010",34673 => "01111010",34674 => "10110101",34675 => "00100000",34676 => "00011101",34677 => "00010100",34678 => "11110011",34679 => "01011101",34680 => "11010000",34681 => "01110100",34682 => "00110011",34683 => "01011100",34684 => "00110110",34685 => "00111011",34686 => "00110001",34687 => "10101001",34688 => "01101000",34689 => "10011011",34690 => "11101101",34691 => "10111110",34692 => "11010011",34693 => "01010011",34694 => "11000010",34695 => "11100001",34696 => "00000010",34697 => "11011110",34698 => "01010110",34699 => "10000011",34700 => "11101100",34701 => "10011011",34702 => "00100010",34703 => "00011101",34704 => "11101011",34705 => "10111001",34706 => "00001100",34707 => "00001110",34708 => "10011000",34709 => "01111100",34710 => "01001110",34711 => "11001011",34712 => "00110010",34713 => "00000101",34714 => "11011100",34715 => "10000100",34716 => "01001010",34717 => "00100000",34718 => "11100001",34719 => "00001010",34720 => "11010000",34721 => "11101100",34722 => "01000011",34723 => "00111110",34724 => "10100100",34725 => "01011111",34726 => "11101011",34727 => "11000011",34728 => "00110010",34729 => "00010011",34730 => "11011000",34731 => "01101111",34732 => "10100011",34733 => "01011000",34734 => "10101001",34735 => "01111101",34736 => "00001010",34737 => "01001000",34738 => "10111000",34739 => "01111000",34740 => "11101100",34741 => "10000101",34742 => "00101011",34743 => "01111101",34744 => "00001000",34745 => "01001110",34746 => "01011101",34747 => "01101110",34748 => "01100000",34749 => "01100100",34750 => "10110000",34751 => "00111000",34752 => "00001110",34753 => "01100100",34754 => "01100111",34755 => "01111111",34756 => "00111101",34757 => "10110100",34758 => "00000111",34759 => "11010100",34760 => "11010011",34761 => "01010010",34762 => "00111100",34763 => "11000100",34764 => "01010100",34765 => "00000010",34766 => "01101010",34767 => "10011011",34768 => "10110000",34769 => "00000101",34770 => "11100110",34771 => "11100000",34772 => "00011100",34773 => "10110011",34774 => "00011101",34775 => "00100001",34776 => "10111100",34777 => "10000110",34778 => "01011100",34779 => "01100011",34780 => "11011100",34781 => "10100111",34782 => "01001110",34783 => "01000000",34784 => "01111001",34785 => "11011001",34786 => "10111000",34787 => "00111001",34788 => "10110011",34789 => "01110001",34790 => "11001001",34791 => "00010001",34792 => "11010001",34793 => "01011010",34794 => "01010010",34795 => "00100000",34796 => "00000111",34797 => "11100110",34798 => "00011011",34799 => "11000111",34800 => "10011010",34801 => "11000100",34802 => "01110110",34803 => "00000100",34804 => "11110011",34805 => "10110011",34806 => "00000111",34807 => "10011111",34808 => "00001001",34809 => "00001111",34810 => "01001001",34811 => "00100111",34812 => "00000100",34813 => "10010001",34814 => "10111101",34815 => "00000000",34816 => "00110100",34817 => "10101010",34818 => "10011101",34819 => "10010001",34820 => "00110100",34821 => "10100101",34822 => "11110111",34823 => "11010011",34824 => "11010011",34825 => "00010000",34826 => "10010001",34827 => "11110111",34828 => "01010011",34829 => "10100110",34830 => "11011011",34831 => "01001000",34832 => "10101110",34833 => "10110111",34834 => "10000100",34835 => "00001101",34836 => "01110010",34837 => "00111101",34838 => "01001000",34839 => "10011010",34840 => "00111011",34841 => "11111000",34842 => "11100000",34843 => "00010011",34844 => "11100001",34845 => "00001110",34846 => "00111000",34847 => "00011101",34848 => "01110111",34849 => "00010111",34850 => "01001111",34851 => "01001011",34852 => "01011000",34853 => "10000011",34854 => "11011000",34855 => "00001111",34856 => "01100011",34857 => "11110010",34858 => "11101010",34859 => "00000000",34860 => "00100100",34861 => "01000111",34862 => "00011000",34863 => "01001000",34864 => "11100101",34865 => "01100101",34866 => "01101001",34867 => "11110111",34868 => "01110001",34869 => "10101000",34870 => "11011111",34871 => "00000000",34872 => "11101010",34873 => "11001010",34874 => "10000100",34875 => "11011010",34876 => "01000001",34877 => "10101101",34878 => "11001000",34879 => "11100100",34880 => "00010101",34881 => "01100110",34882 => "10110010",34883 => "00100010",34884 => "11001010",34885 => "11001100",34886 => "01010100",34887 => "00000111",34888 => "00100010",34889 => "10010110",34890 => "01101011",34891 => "01111001",34892 => "11011001",34893 => "01111100",34894 => "00011001",34895 => "00010011",34896 => "10110011",34897 => "10111100",34898 => "10101000",34899 => "01010000",34900 => "01111000",34901 => "11001101",34902 => "11000100",34903 => "11100101",34904 => "00111001",34905 => "00001011",34906 => "01000111",34907 => "11101000",34908 => "11011000",34909 => "10101101",34910 => "10101011",34911 => "00010111",34912 => "11011010",34913 => "01110000",34914 => "00010001",34915 => "00110010",34916 => "10001000",34917 => "01010111",34918 => "11001001",34919 => "01101111",34920 => "11011110",34921 => "00001101",34922 => "00101000",34923 => "00010011",34924 => "01011010",34925 => "01011111",34926 => "00011110",34927 => "10000001",34928 => "10101110",34929 => "00100101",34930 => "11000011",34931 => "00110010",34932 => "11111100",34933 => "00100101",34934 => "00111110",34935 => "00110011",34936 => "01110011",34937 => "00011101",34938 => "11100011",34939 => "11000001",34940 => "01101010",34941 => "11011011",34942 => "11011110",34943 => "01010011",34944 => "10001101",34945 => "01111110",34946 => "00000100",34947 => "00110100",34948 => "11001000",34949 => "10111010",34950 => "11110001",34951 => "10011011",34952 => "10000011",34953 => "01111001",34954 => "01101001",34955 => "11100100",34956 => "01101010",34957 => "10111011",34958 => "11011111",34959 => "10110101",34960 => "11001010",34961 => "01011001",34962 => "01100010",34963 => "11010100",34964 => "10100111",34965 => "11010000",34966 => "00010001",34967 => "11110101",34968 => "10010111",34969 => "10110100",34970 => "11111111",34971 => "11001111",34972 => "01110001",34973 => "10010001",34974 => "11111010",34975 => "11011110",34976 => "01010111",34977 => "10010100",34978 => "11101010",34979 => "11001100",34980 => "11010111",34981 => "01000001",34982 => "00001101",34983 => "10011100",34984 => "01101101",34985 => "10101011",34986 => "10000000",34987 => "01111111",34988 => "00010001",34989 => "01110010",34990 => "10000100",34991 => "11011110",34992 => "10110001",34993 => "00100000",34994 => "11100110",34995 => "11010101",34996 => "10001011",34997 => "11010011",34998 => "01111010",34999 => "00000011",35000 => "11011010",35001 => "10000111",35002 => "11111110",35003 => "10111101",35004 => "10010101",35005 => "11110110",35006 => "01110100",35007 => "11101011",35008 => "00001000",35009 => "10101100",35010 => "01011101",35011 => "10010111",35012 => "11000110",35013 => "01101010",35014 => "11001010",35015 => "01110001",35016 => "11101000",35017 => "01111101",35018 => "01001000",35019 => "11100101",35020 => "11111101",35021 => "10001111",35022 => "11010111",35023 => "00000010",35024 => "01101010",35025 => "10011100",35026 => "00001001",35027 => "10100001",35028 => "01111100",35029 => "10101111",35030 => "10001110",35031 => "11001011",35032 => "00010011",35033 => "10000001",35034 => "11000010",35035 => "10001110",35036 => "10000010",35037 => "01111000",35038 => "11111101",35039 => "00101101",35040 => "11000000",35041 => "00001010",35042 => "11010101",35043 => "00001101",35044 => "11100001",35045 => "11110111",35046 => "11100110",35047 => "11100011",35048 => "01011000",35049 => "00001010",35050 => "01000101",35051 => "01000001",35052 => "10110100",35053 => "00000010",35054 => "01110001",35055 => "10011111",35056 => "11011011",35057 => "01010001",35058 => "11010101",35059 => "00110010",35060 => "10101001",35061 => "11000101",35062 => "10011000",35063 => "01101100",35064 => "01100000",35065 => "01101010",35066 => "00000001",35067 => "10010100",35068 => "00011110",35069 => "01010110",35070 => "10100101",35071 => "10001111",35072 => "01011011",35073 => "10011010",35074 => "10011010",35075 => "11111001",35076 => "10011010",35077 => "00100101",35078 => "00101000",35079 => "01000001",35080 => "00010011",35081 => "10011101",35082 => "00110001",35083 => "00110100",35084 => "11011000",35085 => "00110100",35086 => "10001011",35087 => "00110010",35088 => "00111110",35089 => "10100001",35090 => "11001100",35091 => "01000110",35092 => "10110110",35093 => "10101100",35094 => "10111101",35095 => "10101000",35096 => "10010111",35097 => "10000001",35098 => "01011110",35099 => "00100011",35100 => "00111001",35101 => "11000101",35102 => "11111100",35103 => "01010001",35104 => "11100000",35105 => "00100110",35106 => "10010101",35107 => "00101001",35108 => "00110010",35109 => "01101011",35110 => "11010001",35111 => "01000010",35112 => "11010000",35113 => "01010000",35114 => "01101100",35115 => "11110011",35116 => "00111011",35117 => "10100101",35118 => "11011000",35119 => "11000110",35120 => "00100100",35121 => "00000101",35122 => "11000110",35123 => "10000001",35124 => "01010010",35125 => "10001110",35126 => "00010000",35127 => "01011010",35128 => "10000111",35129 => "01110011",35130 => "01011000",35131 => "10111001",35132 => "10110101",35133 => "11110000",35134 => "10011010",35135 => "11010100",35136 => "11110010",35137 => "10111000",35138 => "11110001",35139 => "11001101",35140 => "01101101",35141 => "11011100",35142 => "00010011",35143 => "11011100",35144 => "10110000",35145 => "01100111",35146 => "00001100",35147 => "01110010",35148 => "10001101",35149 => "10010000",35150 => "01101000",35151 => "11100011",35152 => "01011111",35153 => "01100000",35154 => "00111111",35155 => "00110101",35156 => "10100110",35157 => "01001001",35158 => "10011010",35159 => "00001100",35160 => "01000111",35161 => "01110000",35162 => "11001000",35163 => "11110110",35164 => "11001001",35165 => "01101110",35166 => "01100110",35167 => "00000100",35168 => "01100001",35169 => "11001001",35170 => "01000011",35171 => "01110011",35172 => "01011010",35173 => "00010010",35174 => "00110000",35175 => "01000100",35176 => "01101101",35177 => "01010110",35178 => "11101001",35179 => "11011100",35180 => "10000010",35181 => "00011101",35182 => "10011010",35183 => "11000001",35184 => "11110001",35185 => "00100111",35186 => "00000001",35187 => "10010010",35188 => "01001101",35189 => "11101010",35190 => "01101000",35191 => "00001110",35192 => "00011000",35193 => "00011001",35194 => "01001110",35195 => "11110010",35196 => "01110111",35197 => "10110111",35198 => "01101110",35199 => "10100000",35200 => "01001111",35201 => "10011100",35202 => "10000010",35203 => "11111010",35204 => "10010001",35205 => "00001101",35206 => "01001101",35207 => "00100101",35208 => "11110110",35209 => "01111110",35210 => "00111000",35211 => "00011000",35212 => "01100011",35213 => "00101111",35214 => "01100000",35215 => "11010101",35216 => "01000111",35217 => "10100010",35218 => "11001111",35219 => "01101110",35220 => "00101101",35221 => "00000101",35222 => "11111111",35223 => "10111000",35224 => "10111001",35225 => "01111010",35226 => "01100101",35227 => "10101011",35228 => "01101000",35229 => "00000000",35230 => "01011101",35231 => "00101011",35232 => "01001000",35233 => "00100101",35234 => "01101001",35235 => "01101100",35236 => "01011011",35237 => "01110010",35238 => "00110000",35239 => "10111111",35240 => "10110110",35241 => "10010100",35242 => "00100111",35243 => "00011000",35244 => "10001000",35245 => "11101000",35246 => "10010100",35247 => "00010000",35248 => "10010100",35249 => "01101000",35250 => "01001001",35251 => "00010111",35252 => "11111101",35253 => "01111100",35254 => "00110011",35255 => "10010101",35256 => "01001101",35257 => "00100100",35258 => "11111011",35259 => "10000001",35260 => "10001010",35261 => "01100111",35262 => "00101010",35263 => "01001000",35264 => "00011010",35265 => "10001001",35266 => "10011001",35267 => "00111001",35268 => "00011100",35269 => "10111110",35270 => "01010001",35271 => "11001100",35272 => "00010000",35273 => "10111101",35274 => "00100011",35275 => "00101110",35276 => "10010100",35277 => "01010111",35278 => "10111000",35279 => "10101010",35280 => "11000110",35281 => "10000011",35282 => "10001001",35283 => "11101100",35284 => "11011010",35285 => "11111110",35286 => "10100000",35287 => "01000011",35288 => "11110011",35289 => "00110011",35290 => "01111100",35291 => "00101010",35292 => "11110010",35293 => "00110001",35294 => "00101011",35295 => "10111101",35296 => "11100101",35297 => "00111101",35298 => "10111110",35299 => "01011111",35300 => "10001000",35301 => "00101100",35302 => "00110010",35303 => "10001011",35304 => "10001000",35305 => "00110010",35306 => "11111000",35307 => "00001001",35308 => "00111010",35309 => "01101110",35310 => "11100100",35311 => "11010101",35312 => "01111001",35313 => "01001100",35314 => "11010010",35315 => "00110011",35316 => "11110111",35317 => "00010011",35318 => "10100100",35319 => "11000011",35320 => "10001110",35321 => "11000101",35322 => "01010110",35323 => "01001110",35324 => "11111000",35325 => "00011001",35326 => "01100111",35327 => "10100110",35328 => "10110111",35329 => "00101110",35330 => "11100011",35331 => "11010001",35332 => "11111110",35333 => "11100100",35334 => "11000001",35335 => "11111111",35336 => "01001101",35337 => "00011000",35338 => "11001110",35339 => "11000011",35340 => "01111011",35341 => "10111100",35342 => "11001100",35343 => "01001010",35344 => "10000111",35345 => "01111110",35346 => "00101110",35347 => "00000110",35348 => "01010111",35349 => "00101010",35350 => "10010100",35351 => "11101011",35352 => "11011110",35353 => "10101001",35354 => "11110010",35355 => "11000001",35356 => "10110010",35357 => "10001010",35358 => "00000110",35359 => "00000000",35360 => "00011011",35361 => "00100101",35362 => "00010111",35363 => "11111101",35364 => "10000101",35365 => "11010101",35366 => "10000111",35367 => "11001011",35368 => "11000111",35369 => "00101100",35370 => "01100010",35371 => "01001010",35372 => "01001110",35373 => "11010000",35374 => "10100000",35375 => "10111100",35376 => "00001101",35377 => "00001011",35378 => "01110000",35379 => "00001111",35380 => "11111001",35381 => "10111010",35382 => "01000000",35383 => "11111010",35384 => "10000111",35385 => "00110100",35386 => "00001001",35387 => "11011000",35388 => "10101101",35389 => "10010110",35390 => "01011011",35391 => "10000010",35392 => "10001001",35393 => "11100010",35394 => "11110001",35395 => "11011000",35396 => "10110100",35397 => "01011101",35398 => "10001100",35399 => "10110110",35400 => "01101110",35401 => "00111111",35402 => "10000011",35403 => "11001000",35404 => "11111110",35405 => "11100111",35406 => "00111000",35407 => "10100111",35408 => "10000111",35409 => "00010111",35410 => "11100000",35411 => "11101011",35412 => "00110111",35413 => "10100011",35414 => "01111100",35415 => "10011111",35416 => "10100111",35417 => "10110100",35418 => "00101111",35419 => "00010101",35420 => "00000110",35421 => "01000011",35422 => "01100011",35423 => "10101100",35424 => "10001000",35425 => "11011101",35426 => "01101100",35427 => "10111010",35428 => "00110001",35429 => "01011101",35430 => "01000110",35431 => "11100101",35432 => "01101101",35433 => "10110110",35434 => "00110000",35435 => "00110001",35436 => "00100101",35437 => "01011011",35438 => "10000010",35439 => "00101000",35440 => "11000111",35441 => "10001001",35442 => "11110100",35443 => "11000111",35444 => "01100001",35445 => "11101101",35446 => "01110111",35447 => "01110000",35448 => "00011100",35449 => "00010011",35450 => "01110001",35451 => "10001001",35452 => "01011000",35453 => "00001100",35454 => "01000101",35455 => "01100000",35456 => "11010011",35457 => "00100110",35458 => "10011110",35459 => "01100110",35460 => "11000111",35461 => "01010101",35462 => "11100011",35463 => "11100100",35464 => "00101011",35465 => "00000011",35466 => "01101010",35467 => "10000010",35468 => "00001001",35469 => "11111011",35470 => "11100001",35471 => "01001111",35472 => "10110001",35473 => "01000101",35474 => "10111000",35475 => "00011101",35476 => "10000010",35477 => "01010100",35478 => "10000000",35479 => "01101011",35480 => "01100001",35481 => "00100011",35482 => "10111100",35483 => "10110100",35484 => "11101111",35485 => "11000011",35486 => "10011100",35487 => "00110100",35488 => "01101011",35489 => "10101010",35490 => "10010111",35491 => "01110101",35492 => "10111011",35493 => "00111101",35494 => "10010011",35495 => "01010100",35496 => "10000010",35497 => "11100110",35498 => "10101110",35499 => "11111100",35500 => "01011001",35501 => "01000101",35502 => "00011010",35503 => "10101000",35504 => "01000110",35505 => "01000000",35506 => "01111100",35507 => "00111010",35508 => "00011001",35509 => "00110100",35510 => "10110110",35511 => "00000000",35512 => "00010101",35513 => "10100001",35514 => "11011011",35515 => "00110111",35516 => "10011001",35517 => "10100101",35518 => "01111010",35519 => "11101001",35520 => "11001001",35521 => "10010010",35522 => "11101100",35523 => "10000011",35524 => "00101101",35525 => "01001010",35526 => "01101101",35527 => "00101100",35528 => "00101011",35529 => "00101100",35530 => "00101000",35531 => "01011111",35532 => "00011000",35533 => "00111000",35534 => "11110010",35535 => "01110000",35536 => "10110101",35537 => "11010010",35538 => "01000111",35539 => "10100101",35540 => "11000100",35541 => "10010010",35542 => "11110101",35543 => "00100100",35544 => "11010101",35545 => "10111111",35546 => "00110110",35547 => "01101101",35548 => "11111101",35549 => "00101100",35550 => "01001000",35551 => "00111001",35552 => "01010001",35553 => "01101111",35554 => "00111010",35555 => "01011011",35556 => "10110110",35557 => "10101101",35558 => "00010100",35559 => "10011011",35560 => "01100111",35561 => "01011011",35562 => "00011101",35563 => "00010010",35564 => "01101001",35565 => "11111111",35566 => "00011111",35567 => "10100101",35568 => "01101110",35569 => "11110010",35570 => "10101110",35571 => "10111011",35572 => "00000011",35573 => "10000001",35574 => "00111010",35575 => "00111101",35576 => "10110101",35577 => "00001101",35578 => "10101111",35579 => "11000000",35580 => "10101111",35581 => "10101101",35582 => "11111101",35583 => "10010111",35584 => "10000111",35585 => "01111101",35586 => "11101010",35587 => "10100100",35588 => "10001001",35589 => "01111110",35590 => "00010111",35591 => "01010100",35592 => "10111000",35593 => "10010001",35594 => "00001000",35595 => "00100100",35596 => "01011011",35597 => "11010000",35598 => "01100011",35599 => "00001010",35600 => "10111111",35601 => "10010000",35602 => "11000110",35603 => "10110001",35604 => "00111010",35605 => "11011011",35606 => "01010011",35607 => "11101110",35608 => "01001111",35609 => "00010101",35610 => "10100110",35611 => "10110010",35612 => "00000010",35613 => "01101001",35614 => "00010010",35615 => "01001110",35616 => "01001001",35617 => "00001000",35618 => "10000110",35619 => "11110100",35620 => "01011100",35621 => "00000001",35622 => "01101100",35623 => "01111111",35624 => "10100000",35625 => "01100000",35626 => "00001111",35627 => "00000011",35628 => "01000000",35629 => "00101001",35630 => "00011000",35631 => "00111011",35632 => "00011001",35633 => "00000000",35634 => "10010001",35635 => "01110001",35636 => "10001011",35637 => "11010011",35638 => "00101100",35639 => "00000000",35640 => "00010100",35641 => "10111110",35642 => "11010111",35643 => "01000101",35644 => "01111111",35645 => "01011110",35646 => "01010100",35647 => "11011000",35648 => "10001110",35649 => "10001100",35650 => "01101000",35651 => "01111000",35652 => "01101000",35653 => "11001100",35654 => "11101001",35655 => "11001010",35656 => "00111110",35657 => "11001110",35658 => "10101011",35659 => "11110101",35660 => "00101110",35661 => "11110001",35662 => "00100101",35663 => "00100101",35664 => "00001101",35665 => "01010011",35666 => "11100111",35667 => "11111101",35668 => "11001111",35669 => "00110101",35670 => "00110110",35671 => "01100000",35672 => "11010001",35673 => "00011010",35674 => "10001011",35675 => "00001110",35676 => "10010000",35677 => "00101010",35678 => "11111010",35679 => "10110000",35680 => "01110011",35681 => "01110011",35682 => "00101101",35683 => "00100110",35684 => "01011100",35685 => "10001100",35686 => "00011000",35687 => "00100010",35688 => "11100010",35689 => "10011111",35690 => "11100101",35691 => "11111100",35692 => "11111101",35693 => "01111000",35694 => "10101101",35695 => "00110000",35696 => "11011110",35697 => "10000110",35698 => "01110010",35699 => "11011101",35700 => "11101101",35701 => "10010001",35702 => "11101010",35703 => "11100000",35704 => "11001111",35705 => "10000111",35706 => "10111011",35707 => "11001000",35708 => "11011001",35709 => "11000111",35710 => "10111101",35711 => "10111011",35712 => "00011000",35713 => "10010101",35714 => "00000101",35715 => "11000111",35716 => "11011011",35717 => "01100101",35718 => "00101000",35719 => "11101100",35720 => "00001100",35721 => "10100100",35722 => "00010111",35723 => "11110110",35724 => "00001011",35725 => "00110001",35726 => "00111110",35727 => "11111110",35728 => "00001001",35729 => "10001101",35730 => "10101000",35731 => "00101100",35732 => "00111111",35733 => "00110100",35734 => "01110101",35735 => "11111101",35736 => "00100100",35737 => "11000000",35738 => "11110100",35739 => "10011011",35740 => "11000001",35741 => "10101001",35742 => "11010000",35743 => "01110110",35744 => "11001111",35745 => "00011001",35746 => "10100101",35747 => "00010011",35748 => "11111010",35749 => "11000111",35750 => "10011011",35751 => "11100100",35752 => "11100000",35753 => "11000001",35754 => "10010000",35755 => "01101101",35756 => "11101011",35757 => "00111010",35758 => "00010000",35759 => "11101101",35760 => "11010000",35761 => "11100100",35762 => "10010110",35763 => "10111100",35764 => "01111101",35765 => "11001001",35766 => "11111100",35767 => "11000100",35768 => "10001000",35769 => "11110100",35770 => "01000001",35771 => "11101011",35772 => "11011010",35773 => "01001110",35774 => "11110001",35775 => "11001011",35776 => "11110101",35777 => "01001011",35778 => "10011010",35779 => "11101110",35780 => "11100110",35781 => "11101011",35782 => "01000101",35783 => "01111100",35784 => "11001100",35785 => "01101110",35786 => "00001110",35787 => "10110110",35788 => "01001001",35789 => "01110110",35790 => "10001100",35791 => "01101011",35792 => "00001011",35793 => "00001001",35794 => "01110001",35795 => "10000100",35796 => "00011110",35797 => "01101010",35798 => "00101100",35799 => "10011010",35800 => "01000011",35801 => "11100011",35802 => "01000000",35803 => "00100001",35804 => "01100000",35805 => "00000110",35806 => "00100101",35807 => "10101111",35808 => "01001110",35809 => "01110101",35810 => "11000001",35811 => "11011010",35812 => "11011111",35813 => "11110110",35814 => "10100101",35815 => "10001100",35816 => "10101001",35817 => "01000100",35818 => "10011101",35819 => "01101100",35820 => "01000101",35821 => "10001101",35822 => "11111010",35823 => "11010010",35824 => "00101000",35825 => "01010110",35826 => "10111001",35827 => "10001101",35828 => "10111001",35829 => "11100101",35830 => "00111100",35831 => "00111001",35832 => "11010111",35833 => "10000000",35834 => "01110101",35835 => "10010100",35836 => "11011001",35837 => "00111000",35838 => "10010001",35839 => "10011000",35840 => "11011011",35841 => "00110001",35842 => "01000010",35843 => "10111100",35844 => "00010010",35845 => "00110011",35846 => "11010110",35847 => "10100011",35848 => "10110001",35849 => "00111110",35850 => "11000100",35851 => "00010010",35852 => "11111000",35853 => "11110010",35854 => "10100111",35855 => "00101000",35856 => "00001011",35857 => "01101001",35858 => "00010101",35859 => "10000100",35860 => "00001100",35861 => "10111010",35862 => "01111001",35863 => "11110110",35864 => "11000100",35865 => "11001100",35866 => "11000111",35867 => "10010101",35868 => "00111000",35869 => "10100100",35870 => "01001100",35871 => "00110110",35872 => "00101101",35873 => "00110011",35874 => "00100000",35875 => "10011110",35876 => "00110011",35877 => "11100100",35878 => "00111001",35879 => "01010110",35880 => "10100100",35881 => "01000001",35882 => "11110110",35883 => "10011111",35884 => "01000001",35885 => "01000100",35886 => "10101011",35887 => "10100011",35888 => "10011110",35889 => "00110101",35890 => "10110001",35891 => "11111101",35892 => "10111011",35893 => "11000001",35894 => "00110000",35895 => "00111111",35896 => "00110110",35897 => "10001110",35898 => "01110101",35899 => "11111110",35900 => "01010111",35901 => "11010010",35902 => "10000010",35903 => "11110011",35904 => "10111010",35905 => "00010101",35906 => "01001110",35907 => "10111110",35908 => "11101010",35909 => "11001100",35910 => "00111101",35911 => "00000100",35912 => "01011111",35913 => "01000000",35914 => "01001000",35915 => "11000101",35916 => "00011100",35917 => "10001101",35918 => "11010101",35919 => "01010001",35920 => "01000100",35921 => "00000110",35922 => "00111000",35923 => "00000100",35924 => "00111111",35925 => "00001111",35926 => "01100001",35927 => "11110001",35928 => "00000110",35929 => "00110111",35930 => "11100011",35931 => "10111011",35932 => "01110011",35933 => "11100111",35934 => "10010111",35935 => "10110001",35936 => "10011100",35937 => "11111010",35938 => "01001100",35939 => "11011001",35940 => "00100100",35941 => "00111111",35942 => "11101100",35943 => "01101110",35944 => "00111011",35945 => "00100000",35946 => "01100011",35947 => "00011100",35948 => "10110100",35949 => "11100110",35950 => "00110100",35951 => "10011110",35952 => "01111100",35953 => "10110001",35954 => "00011101",35955 => "00110000",35956 => "10111010",35957 => "01110011",35958 => "10011101",35959 => "01111000",35960 => "10010001",35961 => "01001000",35962 => "01001001",35963 => "00011010",35964 => "00111100",35965 => "11001001",35966 => "01100110",35967 => "11101010",35968 => "11011011",35969 => "00000011",35970 => "11100101",35971 => "10010111",35972 => "01010100",35973 => "11110111",35974 => "10100100",35975 => "01110111",35976 => "10111010",35977 => "01010011",35978 => "00001100",35979 => "01111011",35980 => "01101111",35981 => "01111110",35982 => "01101001",35983 => "11001011",35984 => "11010101",35985 => "00111100",35986 => "11101001",35987 => "00110101",35988 => "11100010",35989 => "11011011",35990 => "10111001",35991 => "11101110",35992 => "10110010",35993 => "01111100",35994 => "01010111",35995 => "11010110",35996 => "11011011",35997 => "00011010",35998 => "00101011",35999 => "01101001",36000 => "10000111",36001 => "01100111",36002 => "00100110",36003 => "11000001",36004 => "00110100",36005 => "00001110",36006 => "01101101",36007 => "11111001",36008 => "10011111",36009 => "01011100",36010 => "01010111",36011 => "01100100",36012 => "11010011",36013 => "00100000",36014 => "10111000",36015 => "01011110",36016 => "10111000",36017 => "11001111",36018 => "01011110",36019 => "11010110",36020 => "11000000",36021 => "00011010",36022 => "01110011",36023 => "01101001",36024 => "00100100",36025 => "00101111",36026 => "00111001",36027 => "00110100",36028 => "01111001",36029 => "10111000",36030 => "01000001",36031 => "00011101",36032 => "01111111",36033 => "10111111",36034 => "01111100",36035 => "10101100",36036 => "00000000",36037 => "01010010",36038 => "11111111",36039 => "10101011",36040 => "10101001",36041 => "10001001",36042 => "11101010",36043 => "11001111",36044 => "11110011",36045 => "00001101",36046 => "01000101",36047 => "01010111",36048 => "10101110",36049 => "01000100",36050 => "10011010",36051 => "10001000",36052 => "10111000",36053 => "11100110",36054 => "01011110",36055 => "00011010",36056 => "01000001",36057 => "10000101",36058 => "01101110",36059 => "00110100",36060 => "11001010",36061 => "01000010",36062 => "10011010",36063 => "00111011",36064 => "10000001",36065 => "00111011",36066 => "01011000",36067 => "00011100",36068 => "11010011",36069 => "00111010",36070 => "10000110",36071 => "01000110",36072 => "00101110",36073 => "01010110",36074 => "10000000",36075 => "00101100",36076 => "00001111",36077 => "00111010",36078 => "01110011",36079 => "11111111",36080 => "01110011",36081 => "11101110",36082 => "11110010",36083 => "10010001",36084 => "01000010",36085 => "01011010",36086 => "00111011",36087 => "11010001",36088 => "01000101",36089 => "00001010",36090 => "10011111",36091 => "01111111",36092 => "01111000",36093 => "10110110",36094 => "01001000",36095 => "11000001",36096 => "01010001",36097 => "10001101",36098 => "00111010",36099 => "11010001",36100 => "11100000",36101 => "01111101",36102 => "00101101",36103 => "10101000",36104 => "00111111",36105 => "01011111",36106 => "01001011",36107 => "00101011",36108 => "00000111",36109 => "10010100",36110 => "00111111",36111 => "11011001",36112 => "10101010",36113 => "00100110",36114 => "00000011",36115 => "11011110",36116 => "01111111",36117 => "01100100",36118 => "00010111",36119 => "11100011",36120 => "00000010",36121 => "01010111",36122 => "11011100",36123 => "11011000",36124 => "10111000",36125 => "01101111",36126 => "01000010",36127 => "00001110",36128 => "10001010",36129 => "01011100",36130 => "01100011",36131 => "00010011",36132 => "11111010",36133 => "10000010",36134 => "10111110",36135 => "01011101",36136 => "00011001",36137 => "00000101",36138 => "01110010",36139 => "10101111",36140 => "10011000",36141 => "10011011",36142 => "01111101",36143 => "11100111",36144 => "10000100",36145 => "01010100",36146 => "00010111",36147 => "00011000",36148 => "01100110",36149 => "11100011",36150 => "01001101",36151 => "10110101",36152 => "11000010",36153 => "11001100",36154 => "11111010",36155 => "00111000",36156 => "11010101",36157 => "01001101",36158 => "11001011",36159 => "10100011",36160 => "11110000",36161 => "10110001",36162 => "00001010",36163 => "11100000",36164 => "00110111",36165 => "00000000",36166 => "11000011",36167 => "00100010",36168 => "11101101",36169 => "01011101",36170 => "00111001",36171 => "11110111",36172 => "00010101",36173 => "11110010",36174 => "10101110",36175 => "01001011",36176 => "00011101",36177 => "00011110",36178 => "11000001",36179 => "11101111",36180 => "11001110",36181 => "11011111",36182 => "00110000",36183 => "01100100",36184 => "01101000",36185 => "01111111",36186 => "00100011",36187 => "01001101",36188 => "11101001",36189 => "11000110",36190 => "10000101",36191 => "00100100",36192 => "01010101",36193 => "10101000",36194 => "11000100",36195 => "01110100",36196 => "01110100",36197 => "01101110",36198 => "10101000",36199 => "10111010",36200 => "00000011",36201 => "11010010",36202 => "10000000",36203 => "00111011",36204 => "01011100",36205 => "01101000",36206 => "01010111",36207 => "11010011",36208 => "01101110",36209 => "00110110",36210 => "00110001",36211 => "11011101",36212 => "01110011",36213 => "11001010",36214 => "11010111",36215 => "00111011",36216 => "11101001",36217 => "10000100",36218 => "10011001",36219 => "10110110",36220 => "00110010",36221 => "00000010",36222 => "01111101",36223 => "10011010",36224 => "11011000",36225 => "11100011",36226 => "00100001",36227 => "11010011",36228 => "11010110",36229 => "01000000",36230 => "00101100",36231 => "00010000",36232 => "10110011",36233 => "11101101",36234 => "10110010",36235 => "11111011",36236 => "10001100",36237 => "11100010",36238 => "11110011",36239 => "10001101",36240 => "01000001",36241 => "10101011",36242 => "11100101",36243 => "01001110",36244 => "11111110",36245 => "11001101",36246 => "11010101",36247 => "01001001",36248 => "10110011",36249 => "00010001",36250 => "00001101",36251 => "01001000",36252 => "00100110",36253 => "01110110",36254 => "10101011",36255 => "00011110",36256 => "10010100",36257 => "10010011",36258 => "00110010",36259 => "11110001",36260 => "01101010",36261 => "10100010",36262 => "01001101",36263 => "01101111",36264 => "00000010",36265 => "00101100",36266 => "01110011",36267 => "10111100",36268 => "01011000",36269 => "01001111",36270 => "00011110",36271 => "10101000",36272 => "10110010",36273 => "11111001",36274 => "01111100",36275 => "11100111",36276 => "11101001",36277 => "01001000",36278 => "11001011",36279 => "11011101",36280 => "01011000",36281 => "11110101",36282 => "00001111",36283 => "01100100",36284 => "11111110",36285 => "01101110",36286 => "00100101",36287 => "00011000",36288 => "10101110",36289 => "01011010",36290 => "11101001",36291 => "00000110",36292 => "11110000",36293 => "10111101",36294 => "10100101",36295 => "01101000",36296 => "01000111",36297 => "10111111",36298 => "10000111",36299 => "00011111",36300 => "11110101",36301 => "11110010",36302 => "00110000",36303 => "11111111",36304 => "10011101",36305 => "00111010",36306 => "00001110",36307 => "01001101",36308 => "10110110",36309 => "11011011",36310 => "00001001",36311 => "01100001",36312 => "00110101",36313 => "00000111",36314 => "00111111",36315 => "01111000",36316 => "01100001",36317 => "11001100",36318 => "01111010",36319 => "00010001",36320 => "11000010",36321 => "00000110",36322 => "11010101",36323 => "00101110",36324 => "00111011",36325 => "11111101",36326 => "00110010",36327 => "01100110",36328 => "10100001",36329 => "00110101",36330 => "11100110",36331 => "00111001",36332 => "01110010",36333 => "00110111",36334 => "00101010",36335 => "01000100",36336 => "00001001",36337 => "00000101",36338 => "10111011",36339 => "01100110",36340 => "00010101",36341 => "10001010",36342 => "11010110",36343 => "01110101",36344 => "11111101",36345 => "10110001",36346 => "11001010",36347 => "10101000",36348 => "11001100",36349 => "11011101",36350 => "01011100",36351 => "00100001",36352 => "00110110",36353 => "10101010",36354 => "00011100",36355 => "11101000",36356 => "11110100",36357 => "10001101",36358 => "01011001",36359 => "00101001",36360 => "11100000",36361 => "11000111",36362 => "01001110",36363 => "01010111",36364 => "10100101",36365 => "11110011",36366 => "11011001",36367 => "01111010",36368 => "01101011",36369 => "10011111",36370 => "01100000",36371 => "00111100",36372 => "10011000",36373 => "10000100",36374 => "00100001",36375 => "11010010",36376 => "11000001",36377 => "01001111",36378 => "10001010",36379 => "10001010",36380 => "10011010",36381 => "11110111",36382 => "10101010",36383 => "00000110",36384 => "01100111",36385 => "11000001",36386 => "00001111",36387 => "00110111",36388 => "00100101",36389 => "11011010",36390 => "11010010",36391 => "10000011",36392 => "11110011",36393 => "11110010",36394 => "00001010",36395 => "00111110",36396 => "10000100",36397 => "01110101",36398 => "00111100",36399 => "01000011",36400 => "01110111",36401 => "11011100",36402 => "01101001",36403 => "00000110",36404 => "10111101",36405 => "01001100",36406 => "11010101",36407 => "00000011",36408 => "10100011",36409 => "10001111",36410 => "01110011",36411 => "10111111",36412 => "11011011",36413 => "11111100",36414 => "00111010",36415 => "01101001",36416 => "00011101",36417 => "01001100",36418 => "10001110",36419 => "00111110",36420 => "10101110",36421 => "10100100",36422 => "01100000",36423 => "00101010",36424 => "11000110",36425 => "10101101",36426 => "01100100",36427 => "10111100",36428 => "11101001",36429 => "11000101",36430 => "10011010",36431 => "01100100",36432 => "11001101",36433 => "01000001",36434 => "10100001",36435 => "11111100",36436 => "00110110",36437 => "00100111",36438 => "00000000",36439 => "10111000",36440 => "11110111",36441 => "10000011",36442 => "00010011",36443 => "00100001",36444 => "00100111",36445 => "01011111",36446 => "10010010",36447 => "01011011",36448 => "00101100",36449 => "11010011",36450 => "11101110",36451 => "10100000",36452 => "11101110",36453 => "00010100",36454 => "11000001",36455 => "00011011",36456 => "11101000",36457 => "10101000",36458 => "11101011",36459 => "10010100",36460 => "10011000",36461 => "01000100",36462 => "10011100",36463 => "01100111",36464 => "00001110",36465 => "01110000",36466 => "00011110",36467 => "00000001",36468 => "11000111",36469 => "00001100",36470 => "00101001",36471 => "01111000",36472 => "00111101",36473 => "00001000",36474 => "11001001",36475 => "11011100",36476 => "01100001",36477 => "00100001",36478 => "10111000",36479 => "00101110",36480 => "01000111",36481 => "00100011",36482 => "00001100",36483 => "10101111",36484 => "00000111",36485 => "01010110",36486 => "00010110",36487 => "01110110",36488 => "10001101",36489 => "11001101",36490 => "00010111",36491 => "10101000",36492 => "11000101",36493 => "11111011",36494 => "11010101",36495 => "11100011",36496 => "10000111",36497 => "01001101",36498 => "10011110",36499 => "01011110",36500 => "00000011",36501 => "10010110",36502 => "11001110",36503 => "11100111",36504 => "00111111",36505 => "00110100",36506 => "10010011",36507 => "01010100",36508 => "01011000",36509 => "00001000",36510 => "10001100",36511 => "10011100",36512 => "10001011",36513 => "01110010",36514 => "10010011",36515 => "11011101",36516 => "11111000",36517 => "00001000",36518 => "01001001",36519 => "01111000",36520 => "00000000",36521 => "00101100",36522 => "01100011",36523 => "01110001",36524 => "01010100",36525 => "01111110",36526 => "01100010",36527 => "10101001",36528 => "00011111",36529 => "11011011",36530 => "01111000",36531 => "00011111",36532 => "01100011",36533 => "01000000",36534 => "00111101",36535 => "11000010",36536 => "00000100",36537 => "10000110",36538 => "11011001",36539 => "01010000",36540 => "11001001",36541 => "01000010",36542 => "01111100",36543 => "01010000",36544 => "00100100",36545 => "10111010",36546 => "10100000",36547 => "01110100",36548 => "11111011",36549 => "01110000",36550 => "00110000",36551 => "00010000",36552 => "11010000",36553 => "11011000",36554 => "01011101",36555 => "01111001",36556 => "11111011",36557 => "01011110",36558 => "00111001",36559 => "10101101",36560 => "01101100",36561 => "00001110",36562 => "01010001",36563 => "01000101",36564 => "01011110",36565 => "10011100",36566 => "00100110",36567 => "11100100",36568 => "11010000",36569 => "00111111",36570 => "00010001",36571 => "10011011",36572 => "10000100",36573 => "10110101",36574 => "01111101",36575 => "10010101",36576 => "11001101",36577 => "01111011",36578 => "00100001",36579 => "10011000",36580 => "01111110",36581 => "01100111",36582 => "11001011",36583 => "00010101",36584 => "11111100",36585 => "01110101",36586 => "00011111",36587 => "10010001",36588 => "10100100",36589 => "10001101",36590 => "10011110",36591 => "00111101",36592 => "00010011",36593 => "11011011",36594 => "11111110",36595 => "11001100",36596 => "10010011",36597 => "11100000",36598 => "00000001",36599 => "10110101",36600 => "10110010",36601 => "00010111",36602 => "10011100",36603 => "01110000",36604 => "00100110",36605 => "01110111",36606 => "01000000",36607 => "10100001",36608 => "00010001",36609 => "10100000",36610 => "01011111",36611 => "00000101",36612 => "11111010",36613 => "10110101",36614 => "10011010",36615 => "01111010",36616 => "00100000",36617 => "10100111",36618 => "10111001",36619 => "11101111",36620 => "01110010",36621 => "01100110",36622 => "10101010",36623 => "11110101",36624 => "00110101",36625 => "01001001",36626 => "00101100",36627 => "10110101",36628 => "00011000",36629 => "01001111",36630 => "10110001",36631 => "11111001",36632 => "10001100",36633 => "10110111",36634 => "11000110",36635 => "01101001",36636 => "10110100",36637 => "10000100",36638 => "11110001",36639 => "11011101",36640 => "10000001",36641 => "10111110",36642 => "01011111",36643 => "10100000",36644 => "11001001",36645 => "00111010",36646 => "01101111",36647 => "10101001",36648 => "01110001",36649 => "10010101",36650 => "10111011",36651 => "11000000",36652 => "10110100",36653 => "11000100",36654 => "10100000",36655 => "10100110",36656 => "00110011",36657 => "00010111",36658 => "11111011",36659 => "10001001",36660 => "10000000",36661 => "00110011",36662 => "11101110",36663 => "10101010",36664 => "11111001",36665 => "01101100",36666 => "00101010",36667 => "00100110",36668 => "00001000",36669 => "10010110",36670 => "01100000",36671 => "01010001",36672 => "11100000",36673 => "10111011",36674 => "11100010",36675 => "10011110",36676 => "01111100",36677 => "01101111",36678 => "00110010",36679 => "11110000",36680 => "10100100",36681 => "11110010",36682 => "01111010",36683 => "01000001",36684 => "00100100",36685 => "10101000",36686 => "00010010",36687 => "01001000",36688 => "00010100",36689 => "00011011",36690 => "01001010",36691 => "11101011",36692 => "00000101",36693 => "01000100",36694 => "10101000",36695 => "10000111",36696 => "11100110",36697 => "10110010",36698 => "01100100",36699 => "10011000",36700 => "00110101",36701 => "00011001",36702 => "00101001",36703 => "00100010",36704 => "01110000",36705 => "00011101",36706 => "10010101",36707 => "01001111",36708 => "00011000",36709 => "11111011",36710 => "00111101",36711 => "10001000",36712 => "00110101",36713 => "00000010",36714 => "00111101",36715 => "11111101",36716 => "00110110",36717 => "10101111",36718 => "10001010",36719 => "11001010",36720 => "11010111",36721 => "00101010",36722 => "10000011",36723 => "01001000",36724 => "10111110",36725 => "10010101",36726 => "10001101",36727 => "10011011",36728 => "10110100",36729 => "10101111",36730 => "10111101",36731 => "10101101",36732 => "00010001",36733 => "00011000",36734 => "01010000",36735 => "01010010",36736 => "11101000",36737 => "10000100",36738 => "00110011",36739 => "10111010",36740 => "11111011",36741 => "00111111",36742 => "00110001",36743 => "00001100",36744 => "01001110",36745 => "00110000",36746 => "10100000",36747 => "10001110",36748 => "01110010",36749 => "00100100",36750 => "00010000",36751 => "01010101",36752 => "00010100",36753 => "00110010",36754 => "10101100",36755 => "10000000",36756 => "10010010",36757 => "11010111",36758 => "00000000",36759 => "00000110",36760 => "11000001",36761 => "11111111",36762 => "10100111",36763 => "10010110",36764 => "11001001",36765 => "10001001",36766 => "11010111",36767 => "01110010",36768 => "01110101",36769 => "01010111",36770 => "01100011",36771 => "11011010",36772 => "10101100",36773 => "01001111",36774 => "00101100",36775 => "01110101",36776 => "11101011",36777 => "01011101",36778 => "00111001",36779 => "01001111",36780 => "00010010",36781 => "11010101",36782 => "00011100",36783 => "00001111",36784 => "01100101",36785 => "10111110",36786 => "10100010",36787 => "11010100",36788 => "10011000",36789 => "01101000",36790 => "11011101",36791 => "11010100",36792 => "00111100",36793 => "11000000",36794 => "11001110",36795 => "00111001",36796 => "00011000",36797 => "00111011",36798 => "01011110",36799 => "01011100",36800 => "00000011",36801 => "10010011",36802 => "11000101",36803 => "01001101",36804 => "10000010",36805 => "10000011",36806 => "11111011",36807 => "11001101",36808 => "00010110",36809 => "10101000",36810 => "01000100",36811 => "00010001",36812 => "01111101",36813 => "01001111",36814 => "11010011",36815 => "10000001",36816 => "01100110",36817 => "01110000",36818 => "10100101",36819 => "11111010",36820 => "11000010",36821 => "00100010",36822 => "01011000",36823 => "00110111",36824 => "11000101",36825 => "11110011",36826 => "01111011",36827 => "10000111",36828 => "01000011",36829 => "11110001",36830 => "00011100",36831 => "10100001",36832 => "11101101",36833 => "10111111",36834 => "11110100",36835 => "01101011",36836 => "00010110",36837 => "01001001",36838 => "01110101",36839 => "00011111",36840 => "10000001",36841 => "00000000",36842 => "10010011",36843 => "10110000",36844 => "10000100",36845 => "11101010",36846 => "01011110",36847 => "00111001",36848 => "00000010",36849 => "10110111",36850 => "01100110",36851 => "10011100",36852 => "00111111",36853 => "01101110",36854 => "00010001",36855 => "11111101",36856 => "11110101",36857 => "11011001",36858 => "01101101",36859 => "00100011",36860 => "01010100",36861 => "01110100",36862 => "11110001",36863 => "00001011",36864 => "01001000",36865 => "01100110",36866 => "00110110",36867 => "00011101",36868 => "01010010",36869 => "11010001",36870 => "01111110",36871 => "00101010",36872 => "11100111",36873 => "10000110",36874 => "00101100",36875 => "01010011",36876 => "11111011",36877 => "10011000",36878 => "00100011",36879 => "00110111",36880 => "01100001",36881 => "10101111",36882 => "01100100",36883 => "00101011",36884 => "10101000",36885 => "00110010",36886 => "00101000",36887 => "10010011",36888 => "10000101",36889 => "00111101",36890 => "00101001",36891 => "00100100",36892 => "11011010",36893 => "00011000",36894 => "10111111",36895 => "10111110",36896 => "00100001",36897 => "10101100",36898 => "10001111",36899 => "01101110",36900 => "01010011",36901 => "10100101",36902 => "10101101",36903 => "00100010",36904 => "01111100",36905 => "10001001",36906 => "10010100",36907 => "01101001",36908 => "01011100",36909 => "10011100",36910 => "00111011",36911 => "11101001",36912 => "01100001",36913 => "01001000",36914 => "01101000",36915 => "11011010",36916 => "10100000",36917 => "00110010",36918 => "01100110",36919 => "10010111",36920 => "00110011",36921 => "10100011",36922 => "00011001",36923 => "01100000",36924 => "10110101",36925 => "01111010",36926 => "10011011",36927 => "00000110",36928 => "00110010",36929 => "11010001",36930 => "00100100",36931 => "00001010",36932 => "10010011",36933 => "10100011",36934 => "01101101",36935 => "01000100",36936 => "00001001",36937 => "10011110",36938 => "11100100",36939 => "00010100",36940 => "10101010",36941 => "00110001",36942 => "01111100",36943 => "10100100",36944 => "01111001",36945 => "11101010",36946 => "11000111",36947 => "00010101",36948 => "00111110",36949 => "11001100",36950 => "00010100",36951 => "01110010",36952 => "11111001",36953 => "00100001",36954 => "00000000",36955 => "10111110",36956 => "01010110",36957 => "10011100",36958 => "10010100",36959 => "10101000",36960 => "11010111",36961 => "10011011",36962 => "01010100",36963 => "00001100",36964 => "10010111",36965 => "11111001",36966 => "00001101",36967 => "00111111",36968 => "00010101",36969 => "01000101",36970 => "01010101",36971 => "10000000",36972 => "10111000",36973 => "00010011",36974 => "10101000",36975 => "10010011",36976 => "11011011",36977 => "10101110",36978 => "11100000",36979 => "01110010",36980 => "01000101",36981 => "00110101",36982 => "01101100",36983 => "01100011",36984 => "00000100",36985 => "10000000",36986 => "10101011",36987 => "00011010",36988 => "00001000",36989 => "00110010",36990 => "01001100",36991 => "11101101",36992 => "11010000",36993 => "11000111",36994 => "11000001",36995 => "10101110",36996 => "00001010",36997 => "11101100",36998 => "10010000",36999 => "01011000",37000 => "00010111",37001 => "01011101",37002 => "01001001",37003 => "01010110",37004 => "00000010",37005 => "11111110",37006 => "10000111",37007 => "11100001",37008 => "00001010",37009 => "01101010",37010 => "11101100",37011 => "11000100",37012 => "11001111",37013 => "00010111",37014 => "11110011",37015 => "00001010",37016 => "00001001",37017 => "10001111",37018 => "00111100",37019 => "11001000",37020 => "11100001",37021 => "10000100",37022 => "01101111",37023 => "10100110",37024 => "11111011",37025 => "11000000",37026 => "01000100",37027 => "01001001",37028 => "10111110",37029 => "11111001",37030 => "11111111",37031 => "00111001",37032 => "11111010",37033 => "10110111",37034 => "10001011",37035 => "10100011",37036 => "00011011",37037 => "01100010",37038 => "11101010",37039 => "00001110",37040 => "10000011",37041 => "11111111",37042 => "01001110",37043 => "10101110",37044 => "01000111",37045 => "00110111",37046 => "01011111",37047 => "00000110",37048 => "01001000",37049 => "11111101",37050 => "11010000",37051 => "10111101",37052 => "11110000",37053 => "11101111",37054 => "01101100",37055 => "10011001",37056 => "00001101",37057 => "11111011",37058 => "10010011",37059 => "11010101",37060 => "00010110",37061 => "01100110",37062 => "01101001",37063 => "01111010",37064 => "11010011",37065 => "00110100",37066 => "00010011",37067 => "11011010",37068 => "00000101",37069 => "11101010",37070 => "10110101",37071 => "10101110",37072 => "10010000",37073 => "11000000",37074 => "11010111",37075 => "10010101",37076 => "10101111",37077 => "01011111",37078 => "00111110",37079 => "00100101",37080 => "01001001",37081 => "10001011",37082 => "00101110",37083 => "11100000",37084 => "10110010",37085 => "11000111",37086 => "01110110",37087 => "01101101",37088 => "01000110",37089 => "00101010",37090 => "11100001",37091 => "01000010",37092 => "00000001",37093 => "10110110",37094 => "00000111",37095 => "11011011",37096 => "10111001",37097 => "00100011",37098 => "00011110",37099 => "10110111",37100 => "00001111",37101 => "11100111",37102 => "00101101",37103 => "01010101",37104 => "10001111",37105 => "00011100",37106 => "01100111",37107 => "00000110",37108 => "01111100",37109 => "01110101",37110 => "11001111",37111 => "10000110",37112 => "01001000",37113 => "01000111",37114 => "11101010",37115 => "01100001",37116 => "10010000",37117 => "00110110",37118 => "00010001",37119 => "00111000",37120 => "01010110",37121 => "10100101",37122 => "10011010",37123 => "01110010",37124 => "10100001",37125 => "11001100",37126 => "01100010",37127 => "01100110",37128 => "10110110",37129 => "10010000",37130 => "00110101",37131 => "11010111",37132 => "01100000",37133 => "00001000",37134 => "01000100",37135 => "01100000",37136 => "00110100",37137 => "11001110",37138 => "00101001",37139 => "00101111",37140 => "00101101",37141 => "01001110",37142 => "10011110",37143 => "11111001",37144 => "00110100",37145 => "00110001",37146 => "01011010",37147 => "10110101",37148 => "10101111",37149 => "11011010",37150 => "01000011",37151 => "00010001",37152 => "01011100",37153 => "10001110",37154 => "11011110",37155 => "01011001",37156 => "10000000",37157 => "10101110",37158 => "10011110",37159 => "11000011",37160 => "11110111",37161 => "11001000",37162 => "10001101",37163 => "00000100",37164 => "00001100",37165 => "10111100",37166 => "11110000",37167 => "11001111",37168 => "01001100",37169 => "11001110",37170 => "00010010",37171 => "01001101",37172 => "10100000",37173 => "10011010",37174 => "11101101",37175 => "10101001",37176 => "00001101",37177 => "00101011",37178 => "11010100",37179 => "01001000",37180 => "11101100",37181 => "10110101",37182 => "00010001",37183 => "10110101",37184 => "11101101",37185 => "11010100",37186 => "00101010",37187 => "01000010",37188 => "00000110",37189 => "00011010",37190 => "10111111",37191 => "00100111",37192 => "11100011",37193 => "10110000",37194 => "10000100",37195 => "10001110",37196 => "11111111",37197 => "10110111",37198 => "11111001",37199 => "11000000",37200 => "11010111",37201 => "10000000",37202 => "10010111",37203 => "00101110",37204 => "01001011",37205 => "00100110",37206 => "01101000",37207 => "10000011",37208 => "11110101",37209 => "11101000",37210 => "01110101",37211 => "10010111",37212 => "11101011",37213 => "01101101",37214 => "10000100",37215 => "01010101",37216 => "11111110",37217 => "10101111",37218 => "10011110",37219 => "11111000",37220 => "01011111",37221 => "00000110",37222 => "11101000",37223 => "11000011",37224 => "01101100",37225 => "01000010",37226 => "00101010",37227 => "11110110",37228 => "00001101",37229 => "10101010",37230 => "11111110",37231 => "11111011",37232 => "11100000",37233 => "01001001",37234 => "00000100",37235 => "00011111",37236 => "11100111",37237 => "00011010",37238 => "10001110",37239 => "11111001",37240 => "11111110",37241 => "11100111",37242 => "00100101",37243 => "01101001",37244 => "11101011",37245 => "00001100",37246 => "00000101",37247 => "00111000",37248 => "01110001",37249 => "01001100",37250 => "01000100",37251 => "00001001",37252 => "11110010",37253 => "01010001",37254 => "00110000",37255 => "10001100",37256 => "11111000",37257 => "11011111",37258 => "10000111",37259 => "11010110",37260 => "01010010",37261 => "00100111",37262 => "01100100",37263 => "01000111",37264 => "00000111",37265 => "11000001",37266 => "11011100",37267 => "10111111",37268 => "00000011",37269 => "11011111",37270 => "00001001",37271 => "00111001",37272 => "11000100",37273 => "00010001",37274 => "01100100",37275 => "00011100",37276 => "01000111",37277 => "11101110",37278 => "10110111",37279 => "11110110",37280 => "11010100",37281 => "01111110",37282 => "10111110",37283 => "10010011",37284 => "11001110",37285 => "10011101",37286 => "11011000",37287 => "01011111",37288 => "10010111",37289 => "10000010",37290 => "00101001",37291 => "10011100",37292 => "10011010",37293 => "11010101",37294 => "00110111",37295 => "00100100",37296 => "11101010",37297 => "10101111",37298 => "10101000",37299 => "11000111",37300 => "11011110",37301 => "10010110",37302 => "01010000",37303 => "00101101",37304 => "00110001",37305 => "10110011",37306 => "00101010",37307 => "11111011",37308 => "11110011",37309 => "00111111",37310 => "10100001",37311 => "00010101",37312 => "01010110",37313 => "00110011",37314 => "10010101",37315 => "01100111",37316 => "11000010",37317 => "00010001",37318 => "11111010",37319 => "01111010",37320 => "11101010",37321 => "00000111",37322 => "11111100",37323 => "11001111",37324 => "00010000",37325 => "10101011",37326 => "11100101",37327 => "11111010",37328 => "01110001",37329 => "01010111",37330 => "01111101",37331 => "10110110",37332 => "10101011",37333 => "11110011",37334 => "11011000",37335 => "11111110",37336 => "10111010",37337 => "01100011",37338 => "00110011",37339 => "00011100",37340 => "11111010",37341 => "00011100",37342 => "00101001",37343 => "00011011",37344 => "10111011",37345 => "01011000",37346 => "01101100",37347 => "01101110",37348 => "11110010",37349 => "00100110",37350 => "01111110",37351 => "01101000",37352 => "11111000",37353 => "01011010",37354 => "11001101",37355 => "10101111",37356 => "01001111",37357 => "10110110",37358 => "10100000",37359 => "11001111",37360 => "11101101",37361 => "11110111",37362 => "01111001",37363 => "10000100",37364 => "01100011",37365 => "01011001",37366 => "11100101",37367 => "01010010",37368 => "10010100",37369 => "11110010",37370 => "10011011",37371 => "00101000",37372 => "11000010",37373 => "01101010",37374 => "11100110",37375 => "01110010",37376 => "01101110",37377 => "00101111",37378 => "10010001",37379 => "11011111",37380 => "10010111",37381 => "10100011",37382 => "11011111",37383 => "00100111",37384 => "01010000",37385 => "01110010",37386 => "00100011",37387 => "10101000",37388 => "10100101",37389 => "11100111",37390 => "00100110",37391 => "00001000",37392 => "01111001",37393 => "00000001",37394 => "10101000",37395 => "10100011",37396 => "10111010",37397 => "10101011",37398 => "01000111",37399 => "01011101",37400 => "10101000",37401 => "01000001",37402 => "00001101",37403 => "01010111",37404 => "01110111",37405 => "01110000",37406 => "00010010",37407 => "01101000",37408 => "00111100",37409 => "00100010",37410 => "01000011",37411 => "10111110",37412 => "01000000",37413 => "11100111",37414 => "01111101",37415 => "01011110",37416 => "10001111",37417 => "10010000",37418 => "10001011",37419 => "00111011",37420 => "01101100",37421 => "00101100",37422 => "10111000",37423 => "10111010",37424 => "00110111",37425 => "11010001",37426 => "00010101",37427 => "00100101",37428 => "00000101",37429 => "00100111",37430 => "01111101",37431 => "00011001",37432 => "00010110",37433 => "10100011",37434 => "11000101",37435 => "01110100",37436 => "01011100",37437 => "10110100",37438 => "00101011",37439 => "11000100",37440 => "01010011",37441 => "11001111",37442 => "01111100",37443 => "01110101",37444 => "00101011",37445 => "00011000",37446 => "01100010",37447 => "01101101",37448 => "00001110",37449 => "01000100",37450 => "00110001",37451 => "01011010",37452 => "00001000",37453 => "10001010",37454 => "11110000",37455 => "10101110",37456 => "00000100",37457 => "01111101",37458 => "00011000",37459 => "10111010",37460 => "11000111",37461 => "11100101",37462 => "01001100",37463 => "11011111",37464 => "10100111",37465 => "00101100",37466 => "10010100",37467 => "10111101",37468 => "11110110",37469 => "11111010",37470 => "10111011",37471 => "01111000",37472 => "10101110",37473 => "10010101",37474 => "11000111",37475 => "10100010",37476 => "10000001",37477 => "10010010",37478 => "10001000",37479 => "00110101",37480 => "01011100",37481 => "00000100",37482 => "01101110",37483 => "00011000",37484 => "01001000",37485 => "10101100",37486 => "00100010",37487 => "01000101",37488 => "10010111",37489 => "00001001",37490 => "01011110",37491 => "11001010",37492 => "11111111",37493 => "10111001",37494 => "01111001",37495 => "00110010",37496 => "10001100",37497 => "01111000",37498 => "10101011",37499 => "11100000",37500 => "10000100",37501 => "01001100",37502 => "00010110",37503 => "11111110",37504 => "00010011",37505 => "01101101",37506 => "00000101",37507 => "10011100",37508 => "11010010",37509 => "00100000",37510 => "00110000",37511 => "11101000",37512 => "00111101",37513 => "10000100",37514 => "00110101",37515 => "01111100",37516 => "11110101",37517 => "11101111",37518 => "11010011",37519 => "01100001",37520 => "11000011",37521 => "11000110",37522 => "01000011",37523 => "11011001",37524 => "10101100",37525 => "01111000",37526 => "00001100",37527 => "00001110",37528 => "00111101",37529 => "00111110",37530 => "00001011",37531 => "10001111",37532 => "00011101",37533 => "01100000",37534 => "11111101",37535 => "11101001",37536 => "10010010",37537 => "00111011",37538 => "10000010",37539 => "01100111",37540 => "10111110",37541 => "11111100",37542 => "10011100",37543 => "01111110",37544 => "01011001",37545 => "00110100",37546 => "01010111",37547 => "10101010",37548 => "01011010",37549 => "01001001",37550 => "00010011",37551 => "11110010",37552 => "00010100",37553 => "01101000",37554 => "01011001",37555 => "00011011",37556 => "11110110",37557 => "00100101",37558 => "11111011",37559 => "01111011",37560 => "00111011",37561 => "00111110",37562 => "00001111",37563 => "00101001",37564 => "11010001",37565 => "01100011",37566 => "11101010",37567 => "00011111",37568 => "00011001",37569 => "10010000",37570 => "11100010",37571 => "00011010",37572 => "01110011",37573 => "01011010",37574 => "10101101",37575 => "01111001",37576 => "11110100",37577 => "10011001",37578 => "10000100",37579 => "11011100",37580 => "00101111",37581 => "01001110",37582 => "00101101",37583 => "10000111",37584 => "00111110",37585 => "10100001",37586 => "01000110",37587 => "10101011",37588 => "10100110",37589 => "10101001",37590 => "11010111",37591 => "11010110",37592 => "00111000",37593 => "01100110",37594 => "11000001",37595 => "10111101",37596 => "01000100",37597 => "10000101",37598 => "00000000",37599 => "00110010",37600 => "01111000",37601 => "10111011",37602 => "10000010",37603 => "01101001",37604 => "10111111",37605 => "10010000",37606 => "11000001",37607 => "00111000",37608 => "01011001",37609 => "11101001",37610 => "11011101",37611 => "01011101",37612 => "00101110",37613 => "11100101",37614 => "01010110",37615 => "00100101",37616 => "10000011",37617 => "11001110",37618 => "10011111",37619 => "10101110",37620 => "01100011",37621 => "00001011",37622 => "01000100",37623 => "00101010",37624 => "00101000",37625 => "10001001",37626 => "11101111",37627 => "10101000",37628 => "01111110",37629 => "00111110",37630 => "00111100",37631 => "10010101",37632 => "10100101",37633 => "10000101",37634 => "10000000",37635 => "00111101",37636 => "11000011",37637 => "11011110",37638 => "01111111",37639 => "10110000",37640 => "10011101",37641 => "01110001",37642 => "10000001",37643 => "01001011",37644 => "10110000",37645 => "00100110",37646 => "11111101",37647 => "01001000",37648 => "00101000",37649 => "00000100",37650 => "00010101",37651 => "11010100",37652 => "00100010",37653 => "00110001",37654 => "11100000",37655 => "01100101",37656 => "01010001",37657 => "11110001",37658 => "11100110",37659 => "00111000",37660 => "01011000",37661 => "10110001",37662 => "01011000",37663 => "01001101",37664 => "01110001",37665 => "10001010",37666 => "11011000",37667 => "10001100",37668 => "10110010",37669 => "10000011",37670 => "00110110",37671 => "00010001",37672 => "00001001",37673 => "00111000",37674 => "01011110",37675 => "11101011",37676 => "00111001",37677 => "10110110",37678 => "00110111",37679 => "11101000",37680 => "00100101",37681 => "01010011",37682 => "10100000",37683 => "11011010",37684 => "11000111",37685 => "01110111",37686 => "11001011",37687 => "01110100",37688 => "11110111",37689 => "01100011",37690 => "11101100",37691 => "10011001",37692 => "10000101",37693 => "00100111",37694 => "00000011",37695 => "01111110",37696 => "10001111",37697 => "00110101",37698 => "11010111",37699 => "10110011",37700 => "00110101",37701 => "11110101",37702 => "00000110",37703 => "10001001",37704 => "10100001",37705 => "01001000",37706 => "00011011",37707 => "11110001",37708 => "01000110",37709 => "10011111",37710 => "01001101",37711 => "00010011",37712 => "01111100",37713 => "11110011",37714 => "00110010",37715 => "00111110",37716 => "10111001",37717 => "00100011",37718 => "11110010",37719 => "01010101",37720 => "01100101",37721 => "01001010",37722 => "00001111",37723 => "10001110",37724 => "10111110",37725 => "00110011",37726 => "10000010",37727 => "11101000",37728 => "01010001",37729 => "01001001",37730 => "00001101",37731 => "01111110",37732 => "11110011",37733 => "00100000",37734 => "00111001",37735 => "11111010",37736 => "10011011",37737 => "10010000",37738 => "11001010",37739 => "10111010",37740 => "11011000",37741 => "00000101",37742 => "00000011",37743 => "01111011",37744 => "01000000",37745 => "01001010",37746 => "00111111",37747 => "11100110",37748 => "01111000",37749 => "10101011",37750 => "10111110",37751 => "11000101",37752 => "11011010",37753 => "10010001",37754 => "00001110",37755 => "01100001",37756 => "10011001",37757 => "10001111",37758 => "01001011",37759 => "10011011",37760 => "00010101",37761 => "00101101",37762 => "11111110",37763 => "10110101",37764 => "11101010",37765 => "11001100",37766 => "01110100",37767 => "00001011",37768 => "10110110",37769 => "10101010",37770 => "00001000",37771 => "11111110",37772 => "00100010",37773 => "01111000",37774 => "00000000",37775 => "11000100",37776 => "00111000",37777 => "00011011",37778 => "01000100",37779 => "10011101",37780 => "10100110",37781 => "00011011",37782 => "11001111",37783 => "01010101",37784 => "10011111",37785 => "11011101",37786 => "00101100",37787 => "11010001",37788 => "11101101",37789 => "10110011",37790 => "11100111",37791 => "01111100",37792 => "01000111",37793 => "01010101",37794 => "11100000",37795 => "00100100",37796 => "00010100",37797 => "00101001",37798 => "11110001",37799 => "01011101",37800 => "00100011",37801 => "11100111",37802 => "00010101",37803 => "01001101",37804 => "00110111",37805 => "11111011",37806 => "11001001",37807 => "01011100",37808 => "01111001",37809 => "00000001",37810 => "01011111",37811 => "10001101",37812 => "01010101",37813 => "00101000",37814 => "10010000",37815 => "00110101",37816 => "10110101",37817 => "00011110",37818 => "00101001",37819 => "00011100",37820 => "11001100",37821 => "00111101",37822 => "00101100",37823 => "10010111",37824 => "11010011",37825 => "11000111",37826 => "01110010",37827 => "10101110",37828 => "11011110",37829 => "10111010",37830 => "10011000",37831 => "01110001",37832 => "00010001",37833 => "11101111",37834 => "10011011",37835 => "00100000",37836 => "11110100",37837 => "00011000",37838 => "00111111",37839 => "11110010",37840 => "10111010",37841 => "01111001",37842 => "00111010",37843 => "01111010",37844 => "00011011",37845 => "10011000",37846 => "00100000",37847 => "01111110",37848 => "01110010",37849 => "10001100",37850 => "10010000",37851 => "10111010",37852 => "01110011",37853 => "00100010",37854 => "11010010",37855 => "10101011",37856 => "01000100",37857 => "10011010",37858 => "11111000",37859 => "11101101",37860 => "00000111",37861 => "00001110",37862 => "01000001",37863 => "11110001",37864 => "00101101",37865 => "00100110",37866 => "10110100",37867 => "01011011",37868 => "01111101",37869 => "11111101",37870 => "11110111",37871 => "00110011",37872 => "11010110",37873 => "00101100",37874 => "11010101",37875 => "11101100",37876 => "01100101",37877 => "11110010",37878 => "01010110",37879 => "01110110",37880 => "11110001",37881 => "10100110",37882 => "11000001",37883 => "01011101",37884 => "01010111",37885 => "00010011",37886 => "10011000",37887 => "00010000",37888 => "01000111",37889 => "10101100",37890 => "10101000",37891 => "11110100",37892 => "11010000",37893 => "10000011",37894 => "10010010",37895 => "00111100",37896 => "11010100",37897 => "10111011",37898 => "01101010",37899 => "01000101",37900 => "10100010",37901 => "10110111",37902 => "11001011",37903 => "11100001",37904 => "00110001",37905 => "00000110",37906 => "10100110",37907 => "10100110",37908 => "01100100",37909 => "00100011",37910 => "01010100",37911 => "10001001",37912 => "11101000",37913 => "11000001",37914 => "10010011",37915 => "00000010",37916 => "00101110",37917 => "10011011",37918 => "00011001",37919 => "11101101",37920 => "10111110",37921 => "11011100",37922 => "11001011",37923 => "11111100",37924 => "00100011",37925 => "11011101",37926 => "00000011",37927 => "00011110",37928 => "00011011",37929 => "00101110",37930 => "00000100",37931 => "10110101",37932 => "10101110",37933 => "11100110",37934 => "10110011",37935 => "10101001",37936 => "11011001",37937 => "00001111",37938 => "10010101",37939 => "11100001",37940 => "00000010",37941 => "01111111",37942 => "01100011",37943 => "00111100",37944 => "00101101",37945 => "10001101",37946 => "10010001",37947 => "11011000",37948 => "10011011",37949 => "11001100",37950 => "01011001",37951 => "00010001",37952 => "10111111",37953 => "11001111",37954 => "11011000",37955 => "01000011",37956 => "11010011",37957 => "11011101",37958 => "01100101",37959 => "01000101",37960 => "01101001",37961 => "00110111",37962 => "11011001",37963 => "10010100",37964 => "10001101",37965 => "10110111",37966 => "01000110",37967 => "10110011",37968 => "10001111",37969 => "11001000",37970 => "01110100",37971 => "11010101",37972 => "10100100",37973 => "10111001",37974 => "10010110",37975 => "01101111",37976 => "01111011",37977 => "01110011",37978 => "01111010",37979 => "01010100",37980 => "01110101",37981 => "01010100",37982 => "00110111",37983 => "01001000",37984 => "00111101",37985 => "00011110",37986 => "01001000",37987 => "00010110",37988 => "10101011",37989 => "10010011",37990 => "11100000",37991 => "10010011",37992 => "10101110",37993 => "11001111",37994 => "10001110",37995 => "00100111",37996 => "01010010",37997 => "00000000",37998 => "10110100",37999 => "11111110",38000 => "00101011",38001 => "01110101",38002 => "01001100",38003 => "01011111",38004 => "00001001",38005 => "00111000",38006 => "00001111",38007 => "11110101",38008 => "00101101",38009 => "10000110",38010 => "11111110",38011 => "00001101",38012 => "11010001",38013 => "01110101",38014 => "00101000",38015 => "01101101",38016 => "10110011",38017 => "10010110",38018 => "11111001",38019 => "01010100",38020 => "10110110",38021 => "00011000",38022 => "00101010",38023 => "11100100",38024 => "10110101",38025 => "10101101",38026 => "11111101",38027 => "10010000",38028 => "11110110",38029 => "11010100",38030 => "00001111",38031 => "01010011",38032 => "01101110",38033 => "11111110",38034 => "10100100",38035 => "10110100",38036 => "01111001",38037 => "11111000",38038 => "10000110",38039 => "11100101",38040 => "01001010",38041 => "00111010",38042 => "00111100",38043 => "01001010",38044 => "11010100",38045 => "00010111",38046 => "10110111",38047 => "01001011",38048 => "11100000",38049 => "01010001",38050 => "01110000",38051 => "01010011",38052 => "10001101",38053 => "10111100",38054 => "11010000",38055 => "01100110",38056 => "01010101",38057 => "01010001",38058 => "01001101",38059 => "01011011",38060 => "10111111",38061 => "11010011",38062 => "01110111",38063 => "10001101",38064 => "01010110",38065 => "01100000",38066 => "10100001",38067 => "10010111",38068 => "00101010",38069 => "11101010",38070 => "01101100",38071 => "01110100",38072 => "00111110",38073 => "00000110",38074 => "00000011",38075 => "00000010",38076 => "11011111",38077 => "00010010",38078 => "10010001",38079 => "01011010",38080 => "11110000",38081 => "11110011",38082 => "00101110",38083 => "11001011",38084 => "10100100",38085 => "01111000",38086 => "01011001",38087 => "00000010",38088 => "01101101",38089 => "11010111",38090 => "10001101",38091 => "00010100",38092 => "01001011",38093 => "11001101",38094 => "10110101",38095 => "00000110",38096 => "01100101",38097 => "01111001",38098 => "11011000",38099 => "01001001",38100 => "10001001",38101 => "10100001",38102 => "00111000",38103 => "01000010",38104 => "00001101",38105 => "11011000",38106 => "10000001",38107 => "11111011",38108 => "11110000",38109 => "01000101",38110 => "00110100",38111 => "00100111",38112 => "11010111",38113 => "11100100",38114 => "00000100",38115 => "00100001",38116 => "01110000",38117 => "01101010",38118 => "00111011",38119 => "00010010",38120 => "10001001",38121 => "11010100",38122 => "10010011",38123 => "00101001",38124 => "00001101",38125 => "01000101",38126 => "11100000",38127 => "10001110",38128 => "11011101",38129 => "10001011",38130 => "00110100",38131 => "11101010",38132 => "01111111",38133 => "10010000",38134 => "10111110",38135 => "11101010",38136 => "10100001",38137 => "11000100",38138 => "10010111",38139 => "01001101",38140 => "11100101",38141 => "10000100",38142 => "10111010",38143 => "01101111",38144 => "00111111",38145 => "01100111",38146 => "11010110",38147 => "10000101",38148 => "10010000",38149 => "01001110",38150 => "11100110",38151 => "01100111",38152 => "01110001",38153 => "00100110",38154 => "00010110",38155 => "11110100",38156 => "10111000",38157 => "01011000",38158 => "00000100",38159 => "01101010",38160 => "10011001",38161 => "10110000",38162 => "01101010",38163 => "10011110",38164 => "00101010",38165 => "00101010",38166 => "00011110",38167 => "01010001",38168 => "10000111",38169 => "10000001",38170 => "00100010",38171 => "10010001",38172 => "00010010",38173 => "00001001",38174 => "10100111",38175 => "10110100",38176 => "11110001",38177 => "10101001",38178 => "01001110",38179 => "10001011",38180 => "00111111",38181 => "00011000",38182 => "10100111",38183 => "11001111",38184 => "11010011",38185 => "01011110",38186 => "00111110",38187 => "00001101",38188 => "01101110",38189 => "11010111",38190 => "01110001",38191 => "00010011",38192 => "11111100",38193 => "00011010",38194 => "11110111",38195 => "11110100",38196 => "10000010",38197 => "11010101",38198 => "10101010",38199 => "11000011",38200 => "01000000",38201 => "11010111",38202 => "10111111",38203 => "00101111",38204 => "01100010",38205 => "01000110",38206 => "10000110",38207 => "01000000",38208 => "11011010",38209 => "01111101",38210 => "10001001",38211 => "01110111",38212 => "11101001",38213 => "11000110",38214 => "11001010",38215 => "00111111",38216 => "10011001",38217 => "01000111",38218 => "10100011",38219 => "00110011",38220 => "00110111",38221 => "11000000",38222 => "01100100",38223 => "01000001",38224 => "00011111",38225 => "00011101",38226 => "10000000",38227 => "00001111",38228 => "10011110",38229 => "00111010",38230 => "11111111",38231 => "10001010",38232 => "00110101",38233 => "10111111",38234 => "01110110",38235 => "00100001",38236 => "10000000",38237 => "00101101",38238 => "10100110",38239 => "01001100",38240 => "00110111",38241 => "00100011",38242 => "11010010",38243 => "01111011",38244 => "11111001",38245 => "00010101",38246 => "01010111",38247 => "01001000",38248 => "00110110",38249 => "00110010",38250 => "10110000",38251 => "10100101",38252 => "01111110",38253 => "10110010",38254 => "10100010",38255 => "10111010",38256 => "00100011",38257 => "00101000",38258 => "11011101",38259 => "01100000",38260 => "11110011",38261 => "10101101",38262 => "11011001",38263 => "01100110",38264 => "11101111",38265 => "10111010",38266 => "01100111",38267 => "01100100",38268 => "10101111",38269 => "00101110",38270 => "00110010",38271 => "10011011",38272 => "11001111",38273 => "00010100",38274 => "10010011",38275 => "11000001",38276 => "01110000",38277 => "01011001",38278 => "01101010",38279 => "01111001",38280 => "00101101",38281 => "11000011",38282 => "01011010",38283 => "00001111",38284 => "11101010",38285 => "00001110",38286 => "00110101",38287 => "00101010",38288 => "11011111",38289 => "11110110",38290 => "11100101",38291 => "11100100",38292 => "00011000",38293 => "00110010",38294 => "01111100",38295 => "01101111",38296 => "00011000",38297 => "11011011",38298 => "10100110",38299 => "11110010",38300 => "11110010",38301 => "10101001",38302 => "01001110",38303 => "01011101",38304 => "00011100",38305 => "00111111",38306 => "10000100",38307 => "01110010",38308 => "10111111",38309 => "01000110",38310 => "10101101",38311 => "01001100",38312 => "11010011",38313 => "01001101",38314 => "00010110",38315 => "11011110",38316 => "11000001",38317 => "01110010",38318 => "00100101",38319 => "10011110",38320 => "01010010",38321 => "10000111",38322 => "11011011",38323 => "01100010",38324 => "11010001",38325 => "00001001",38326 => "01001010",38327 => "10001010",38328 => "11001100",38329 => "00000101",38330 => "00001111",38331 => "10011101",38332 => "10000100",38333 => "10010010",38334 => "10100101",38335 => "11000000",38336 => "11100010",38337 => "10111101",38338 => "11100111",38339 => "01011110",38340 => "00110100",38341 => "10010011",38342 => "10110110",38343 => "10010011",38344 => "11100001",38345 => "10101010",38346 => "11110010",38347 => "01010101",38348 => "10110011",38349 => "10110001",38350 => "00110111",38351 => "10011001",38352 => "00111000",38353 => "11100110",38354 => "00011110",38355 => "10110110",38356 => "00111101",38357 => "00110001",38358 => "01110101",38359 => "10001110",38360 => "00011101",38361 => "01110011",38362 => "01000100",38363 => "01000110",38364 => "10001100",38365 => "11000101",38366 => "10110101",38367 => "01011010",38368 => "11000011",38369 => "01001111",38370 => "10100001",38371 => "01011101",38372 => "10100110",38373 => "00101100",38374 => "10001000",38375 => "10101000",38376 => "00011110",38377 => "11111011",38378 => "10001111",38379 => "10110001",38380 => "00010111",38381 => "11111010",38382 => "00101000",38383 => "11011100",38384 => "01100000",38385 => "11101010",38386 => "11111111",38387 => "00101001",38388 => "11011111",38389 => "10011011",38390 => "01101010",38391 => "10000100",38392 => "00011000",38393 => "01000001",38394 => "10111110",38395 => "00011111",38396 => "00100011",38397 => "10100010",38398 => "11001100",38399 => "00000101",38400 => "01110100",38401 => "11101011",38402 => "11010100",38403 => "10101001",38404 => "10011011",38405 => "00011000",38406 => "11101110",38407 => "00000111",38408 => "01010011",38409 => "00010011",38410 => "00000111",38411 => "00001101",38412 => "11100010",38413 => "01101000",38414 => "10011101",38415 => "00111110",38416 => "00010101",38417 => "11001000",38418 => "00001100",38419 => "10011010",38420 => "00001000",38421 => "00000010",38422 => "01001110",38423 => "10100000",38424 => "11110010",38425 => "11100010",38426 => "00100001",38427 => "00100001",38428 => "01010110",38429 => "01100000",38430 => "10001000",38431 => "10001010",38432 => "01101111",38433 => "11110011",38434 => "01000000",38435 => "01100010",38436 => "11000001",38437 => "00111100",38438 => "01011101",38439 => "01101110",38440 => "10111010",38441 => "11100000",38442 => "00110001",38443 => "00001011",38444 => "10010011",38445 => "11100111",38446 => "10011101",38447 => "00111111",38448 => "00000110",38449 => "11111000",38450 => "01101011",38451 => "10010001",38452 => "11011110",38453 => "00000111",38454 => "10111011",38455 => "00000001",38456 => "00011011",38457 => "10110110",38458 => "10111000",38459 => "00101011",38460 => "10011000",38461 => "00010100",38462 => "11100010",38463 => "10100100",38464 => "11001101",38465 => "11110001",38466 => "10100110",38467 => "00010000",38468 => "10011110",38469 => "11101100",38470 => "11101110",38471 => "00111010",38472 => "01001110",38473 => "10111010",38474 => "10000001",38475 => "10010100",38476 => "00100001",38477 => "11011001",38478 => "01110010",38479 => "11111011",38480 => "11100100",38481 => "11000000",38482 => "10011001",38483 => "01111101",38484 => "00101100",38485 => "10011011",38486 => "11001101",38487 => "10001100",38488 => "01011000",38489 => "01110111",38490 => "01100110",38491 => "01011101",38492 => "11101010",38493 => "10101000",38494 => "11111010",38495 => "01001101",38496 => "10110101",38497 => "01011110",38498 => "11100001",38499 => "00001110",38500 => "11111110",38501 => "10010110",38502 => "01100010",38503 => "10101010",38504 => "01000100",38505 => "01000001",38506 => "00000111",38507 => "11100000",38508 => "10011010",38509 => "01010011",38510 => "00101011",38511 => "10101101",38512 => "10001010",38513 => "00001100",38514 => "01011011",38515 => "00101011",38516 => "10000001",38517 => "11001011",38518 => "00100000",38519 => "00101001",38520 => "10111001",38521 => "00011011",38522 => "11011110",38523 => "00100101",38524 => "00001110",38525 => "00111010",38526 => "11001101",38527 => "11000100",38528 => "10010000",38529 => "01000010",38530 => "01110011",38531 => "01000010",38532 => "11001101",38533 => "01110100",38534 => "01000101",38535 => "10011100",38536 => "11011110",38537 => "01001000",38538 => "00000010",38539 => "11101000",38540 => "01101100",38541 => "11011111",38542 => "10001111",38543 => "01100111",38544 => "11011101",38545 => "00000101",38546 => "10101001",38547 => "01010000",38548 => "11010001",38549 => "00100111",38550 => "01000000",38551 => "10000101",38552 => "01110111",38553 => "00111011",38554 => "01001001",38555 => "00111100",38556 => "00011110",38557 => "11101001",38558 => "10010111",38559 => "00001010",38560 => "11000111",38561 => "10001100",38562 => "00001001",38563 => "10001101",38564 => "01110011",38565 => "00101111",38566 => "01000101",38567 => "10101100",38568 => "00010100",38569 => "10100001",38570 => "10101111",38571 => "01010011",38572 => "00001111",38573 => "00001011",38574 => "00111011",38575 => "10110100",38576 => "10101010",38577 => "00110100",38578 => "11111001",38579 => "10101001",38580 => "01100110",38581 => "00000011",38582 => "00011010",38583 => "11100010",38584 => "01110011",38585 => "01001111",38586 => "00110011",38587 => "11111111",38588 => "01100010",38589 => "01010110",38590 => "00110101",38591 => "01111101",38592 => "10111000",38593 => "00100100",38594 => "00101011",38595 => "00101011",38596 => "11111100",38597 => "10100010",38598 => "01100011",38599 => "10101101",38600 => "11010000",38601 => "00111111",38602 => "11110111",38603 => "11100100",38604 => "11000010",38605 => "01000110",38606 => "11110100",38607 => "01011101",38608 => "11101111",38609 => "10101111",38610 => "01010010",38611 => "00000010",38612 => "10001100",38613 => "01111011",38614 => "11110100",38615 => "11110110",38616 => "11110110",38617 => "11001110",38618 => "10101101",38619 => "10111101",38620 => "00111110",38621 => "00101110",38622 => "10110111",38623 => "11010001",38624 => "00110101",38625 => "10100100",38626 => "01110010",38627 => "00001000",38628 => "00110111",38629 => "00010011",38630 => "01100011",38631 => "00100100",38632 => "00101100",38633 => "10001100",38634 => "01010101",38635 => "01010011",38636 => "10011101",38637 => "00001110",38638 => "11101000",38639 => "11010110",38640 => "10101100",38641 => "10000011",38642 => "00100001",38643 => "11001001",38644 => "11100111",38645 => "10010000",38646 => "00011110",38647 => "11010000",38648 => "01000001",38649 => "11001010",38650 => "01001110",38651 => "11100110",38652 => "10111001",38653 => "11010001",38654 => "00100101",38655 => "01010001",38656 => "11011100",38657 => "01101100",38658 => "00110111",38659 => "11011100",38660 => "01100001",38661 => "11100011",38662 => "00011000",38663 => "01001011",38664 => "10101010",38665 => "00110010",38666 => "11101110",38667 => "10110000",38668 => "10010000",38669 => "01110100",38670 => "11001011",38671 => "00000101",38672 => "00010000",38673 => "01100011",38674 => "11011000",38675 => "10011101",38676 => "11011101",38677 => "11011000",38678 => "00101000",38679 => "10101010",38680 => "10101001",38681 => "00000100",38682 => "00001001",38683 => "10010101",38684 => "11001110",38685 => "01011011",38686 => "01100101",38687 => "00111001",38688 => "01100101",38689 => "11111011",38690 => "10011001",38691 => "10001110",38692 => "01011000",38693 => "11010011",38694 => "11110001",38695 => "11010100",38696 => "10111011",38697 => "10111101",38698 => "01010011",38699 => "00100110",38700 => "10001010",38701 => "11110000",38702 => "11110111",38703 => "10110000",38704 => "10101111",38705 => "01100011",38706 => "10101111",38707 => "11111011",38708 => "10101011",38709 => "11101100",38710 => "10010001",38711 => "10111111",38712 => "11110100",38713 => "10110001",38714 => "11001000",38715 => "01111000",38716 => "11101010",38717 => "00010100",38718 => "00100110",38719 => "00110110",38720 => "10000000",38721 => "11000011",38722 => "11101010",38723 => "01111111",38724 => "00111011",38725 => "01011011",38726 => "11100011",38727 => "00111000",38728 => "01011111",38729 => "10110001",38730 => "01001110",38731 => "11101110",38732 => "00001011",38733 => "11110111",38734 => "11100010",38735 => "01000110",38736 => "01001101",38737 => "11011101",38738 => "00011101",38739 => "10100101",38740 => "11100100",38741 => "11111100",38742 => "00101101",38743 => "01101111",38744 => "00111111",38745 => "11011010",38746 => "11000001",38747 => "00011011",38748 => "00101010",38749 => "00111001",38750 => "11111000",38751 => "01010101",38752 => "10100000",38753 => "00101100",38754 => "11000011",38755 => "10100000",38756 => "00110010",38757 => "01001001",38758 => "00110001",38759 => "01110010",38760 => "00111100",38761 => "00000111",38762 => "11011000",38763 => "10010100",38764 => "00000110",38765 => "01100111",38766 => "10111000",38767 => "11001001",38768 => "10010101",38769 => "10000011",38770 => "11110100",38771 => "00100101",38772 => "01000001",38773 => "01110110",38774 => "01111111",38775 => "00001110",38776 => "11111001",38777 => "00011110",38778 => "11100011",38779 => "10100011",38780 => "11100100",38781 => "10101000",38782 => "11101111",38783 => "11011111",38784 => "11110000",38785 => "10001001",38786 => "10001011",38787 => "11110110",38788 => "11101100",38789 => "10100101",38790 => "00101001",38791 => "10100101",38792 => "10100011",38793 => "11101010",38794 => "10010000",38795 => "00110011",38796 => "11100000",38797 => "10011100",38798 => "01101111",38799 => "00011101",38800 => "00010010",38801 => "00110110",38802 => "10100111",38803 => "00001000",38804 => "10111010",38805 => "01100010",38806 => "10101011",38807 => "11001101",38808 => "01011001",38809 => "11001011",38810 => "11100011",38811 => "11011001",38812 => "10001011",38813 => "01001111",38814 => "00110110",38815 => "00011011",38816 => "10110111",38817 => "01010011",38818 => "01000111",38819 => "01001110",38820 => "00000111",38821 => "01111000",38822 => "11001111",38823 => "11000111",38824 => "11011000",38825 => "00000101",38826 => "01111011",38827 => "11110001",38828 => "01001110",38829 => "10011100",38830 => "11000001",38831 => "11010111",38832 => "00110000",38833 => "01111101",38834 => "01110111",38835 => "10101111",38836 => "01000010",38837 => "01111110",38838 => "01010001",38839 => "00110011",38840 => "11101001",38841 => "00011001",38842 => "10100011",38843 => "11110010",38844 => "11011011",38845 => "01111011",38846 => "00101111",38847 => "11010010",38848 => "10010101",38849 => "00101010",38850 => "01011111",38851 => "00101010",38852 => "00011110",38853 => "01111011",38854 => "11011101",38855 => "11100011",38856 => "00001110",38857 => "01111101",38858 => "10001100",38859 => "00001001",38860 => "10111100",38861 => "11101001",38862 => "00000110",38863 => "00010110",38864 => "11000101",38865 => "10000110",38866 => "10011110",38867 => "10001111",38868 => "10001110",38869 => "11000101",38870 => "01101011",38871 => "10110100",38872 => "11001010",38873 => "00101001",38874 => "00011101",38875 => "11000111",38876 => "11000111",38877 => "10011001",38878 => "00111110",38879 => "10110010",38880 => "10100111",38881 => "11011100",38882 => "11010101",38883 => "01111001",38884 => "10101011",38885 => "10000101",38886 => "11010111",38887 => "11011111",38888 => "00011101",38889 => "00001111",38890 => "00011000",38891 => "01110001",38892 => "11101010",38893 => "00111111",38894 => "00101100",38895 => "01101010",38896 => "01010001",38897 => "00001000",38898 => "10111110",38899 => "11100010",38900 => "00001011",38901 => "01001001",38902 => "10111000",38903 => "11111010",38904 => "10100000",38905 => "00101000",38906 => "11101010",38907 => "10111000",38908 => "11111101",38909 => "01101010",38910 => "11100111",38911 => "11101010",38912 => "11001110",38913 => "01000011",38914 => "10110011",38915 => "01111000",38916 => "10000010",38917 => "10011010",38918 => "10110101",38919 => "10000000",38920 => "10101000",38921 => "01110111",38922 => "00000000",38923 => "00001001",38924 => "01001101",38925 => "00110111",38926 => "01001110",38927 => "00101111",38928 => "10110100",38929 => "10111110",38930 => "01010101",38931 => "00110010",38932 => "01000001",38933 => "10100111",38934 => "10000000",38935 => "00000110",38936 => "11100011",38937 => "10011111",38938 => "10100011",38939 => "01011010",38940 => "11001110",38941 => "10011000",38942 => "00010110",38943 => "00011101",38944 => "01101110",38945 => "10010010",38946 => "11000010",38947 => "01101101",38948 => "01010111",38949 => "11100101",38950 => "11101110",38951 => "00100111",38952 => "10010001",38953 => "01001111",38954 => "11011010",38955 => "01111010",38956 => "00110111",38957 => "00010110",38958 => "01011100",38959 => "10001010",38960 => "10100011",38961 => "11011101",38962 => "10001010",38963 => "11011010",38964 => "01000010",38965 => "01101101",38966 => "11011000",38967 => "11100101",38968 => "00110001",38969 => "00101010",38970 => "01111000",38971 => "10110110",38972 => "11000000",38973 => "10001100",38974 => "10001001",38975 => "10001001",38976 => "11100111",38977 => "01111100",38978 => "11001001",38979 => "01100101",38980 => "00100010",38981 => "01001110",38982 => "01011111",38983 => "11010001",38984 => "00100110",38985 => "11000011",38986 => "11001001",38987 => "01000101",38988 => "10100010",38989 => "11111100",38990 => "01010011",38991 => "00111101",38992 => "01100011",38993 => "11111110",38994 => "00001111",38995 => "11110101",38996 => "00111001",38997 => "00001110",38998 => "11001111",38999 => "01111000",39000 => "10111111",39001 => "00100000",39002 => "10110011",39003 => "00001011",39004 => "10001111",39005 => "10001100",39006 => "01001110",39007 => "10101000",39008 => "10011100",39009 => "11010000",39010 => "11111010",39011 => "00010000",39012 => "01111111",39013 => "10110001",39014 => "01110101",39015 => "10110110",39016 => "10111101",39017 => "00101001",39018 => "00111011",39019 => "11010111",39020 => "10001011",39021 => "00111011",39022 => "01001000",39023 => "01110101",39024 => "00100111",39025 => "00110000",39026 => "00010100",39027 => "00110000",39028 => "01001110",39029 => "11101110",39030 => "00101001",39031 => "00000111",39032 => "11000010",39033 => "01001100",39034 => "01010100",39035 => "00110011",39036 => "00000101",39037 => "00011000",39038 => "00101010",39039 => "01101100",39040 => "00011111",39041 => "10001100",39042 => "11001011",39043 => "01110100",39044 => "00100100",39045 => "11110100",39046 => "10101100",39047 => "11110101",39048 => "01001001",39049 => "10101001",39050 => "01000110",39051 => "01011100",39052 => "01000100",39053 => "11000000",39054 => "00000011",39055 => "10111011",39056 => "00100000",39057 => "10000011",39058 => "10011001",39059 => "01010001",39060 => "11100001",39061 => "00010101",39062 => "11011101",39063 => "00001010",39064 => "01111001",39065 => "00111110",39066 => "00101111",39067 => "00000100",39068 => "11101001",39069 => "10010111",39070 => "11000010",39071 => "00011111",39072 => "01011100",39073 => "01110011",39074 => "00111111",39075 => "10011000",39076 => "10100101",39077 => "11110101",39078 => "01100110",39079 => "10110110",39080 => "00000001",39081 => "01100111",39082 => "01110011",39083 => "11001011",39084 => "10101111",39085 => "11000000",39086 => "01000000",39087 => "01110011",39088 => "00001111",39089 => "11100100",39090 => "10101010",39091 => "01110010",39092 => "01100001",39093 => "00000000",39094 => "10011000",39095 => "01011100",39096 => "11000111",39097 => "01000100",39098 => "00011000",39099 => "11010101",39100 => "10110011",39101 => "11001110",39102 => "10100100",39103 => "01101110",39104 => "11001101",39105 => "00100111",39106 => "11010011",39107 => "11100101",39108 => "11000001",39109 => "11101011",39110 => "11011011",39111 => "11111110",39112 => "00100101",39113 => "01000011",39114 => "10001111",39115 => "00000110",39116 => "10101011",39117 => "11111100",39118 => "00100111",39119 => "11010011",39120 => "11111010",39121 => "10011110",39122 => "01001110",39123 => "11111101",39124 => "00000110",39125 => "10001100",39126 => "11100000",39127 => "10011010",39128 => "11010110",39129 => "11100011",39130 => "11101110",39131 => "00010011",39132 => "01001100",39133 => "10100100",39134 => "11101000",39135 => "00011111",39136 => "00001111",39137 => "00111100",39138 => "00001001",39139 => "01100101",39140 => "00001101",39141 => "11001010",39142 => "01011101",39143 => "11100010",39144 => "11110110",39145 => "10100000",39146 => "00111101",39147 => "11011111",39148 => "11000101",39149 => "01000000",39150 => "10110001",39151 => "11101110",39152 => "00110010",39153 => "01110101",39154 => "10111111",39155 => "10010111",39156 => "00110001",39157 => "01010001",39158 => "01101100",39159 => "01011110",39160 => "00010101",39161 => "00000010",39162 => "10101101",39163 => "01011101",39164 => "00011010",39165 => "01010010",39166 => "00100010",39167 => "10101110",39168 => "10111001",39169 => "00011011",39170 => "00111010",39171 => "11101010",39172 => "11110110",39173 => "11000111",39174 => "10110010",39175 => "10001111",39176 => "11000100",39177 => "11101101",39178 => "00100101",39179 => "11001100",39180 => "00101111",39181 => "00010001",39182 => "11000111",39183 => "01111110",39184 => "11000101",39185 => "11101000",39186 => "00100110",39187 => "01001011",39188 => "11001100",39189 => "11010000",39190 => "10010010",39191 => "10111000",39192 => "11010011",39193 => "11000110",39194 => "00011011",39195 => "10111101",39196 => "00001000",39197 => "00110000",39198 => "00000010",39199 => "00111001",39200 => "01111101",39201 => "01011101",39202 => "00100101",39203 => "11010100",39204 => "11111110",39205 => "00011001",39206 => "01111000",39207 => "10100100",39208 => "01100110",39209 => "00111111",39210 => "00000111",39211 => "00011000",39212 => "00010100",39213 => "11010100",39214 => "11001000",39215 => "00011010",39216 => "11100111",39217 => "01001011",39218 => "10001101",39219 => "01110011",39220 => "01100011",39221 => "11101010",39222 => "00111100",39223 => "11010000",39224 => "10101010",39225 => "11110110",39226 => "11110011",39227 => "11100100",39228 => "01001011",39229 => "00111101",39230 => "00101100",39231 => "11001000",39232 => "10010010",39233 => "00011001",39234 => "01000001",39235 => "01110001",39236 => "00111011",39237 => "01101111",39238 => "00011001",39239 => "00111011",39240 => "11110111",39241 => "10100111",39242 => "11001010",39243 => "10110000",39244 => "11111001",39245 => "11000011",39246 => "11101100",39247 => "11100010",39248 => "00100111",39249 => "00011110",39250 => "11111011",39251 => "00011000",39252 => "10011000",39253 => "10110111",39254 => "10011100",39255 => "11011010",39256 => "01011111",39257 => "10000101",39258 => "11101001",39259 => "00001000",39260 => "11111011",39261 => "11001111",39262 => "00000100",39263 => "00100111",39264 => "11101010",39265 => "01011000",39266 => "11110110",39267 => "11101111",39268 => "11100001",39269 => "10011011",39270 => "11010110",39271 => "11110010",39272 => "00011010",39273 => "11010111",39274 => "11100110",39275 => "01101000",39276 => "00011011",39277 => "10011000",39278 => "11000000",39279 => "01111001",39280 => "01011111",39281 => "10001011",39282 => "10010000",39283 => "01011100",39284 => "10011100",39285 => "01110101",39286 => "01111101",39287 => "10011001",39288 => "11111011",39289 => "11101100",39290 => "00100000",39291 => "10001110",39292 => "11100010",39293 => "01000000",39294 => "01111010",39295 => "10011110",39296 => "11010010",39297 => "01001110",39298 => "11001110",39299 => "01000101",39300 => "10000111",39301 => "10101100",39302 => "01001100",39303 => "01111011",39304 => "11110101",39305 => "01011011",39306 => "00001010",39307 => "10000000",39308 => "11000001",39309 => "00001010",39310 => "01101001",39311 => "00000010",39312 => "11101100",39313 => "01000110",39314 => "10110100",39315 => "11100100",39316 => "10101000",39317 => "01010110",39318 => "10011001",39319 => "11101100",39320 => "00110011",39321 => "01101011",39322 => "00011000",39323 => "10101100",39324 => "11011010",39325 => "01000011",39326 => "10001010",39327 => "01110010",39328 => "10011000",39329 => "11110000",39330 => "01111110",39331 => "01101111",39332 => "00010010",39333 => "01000110",39334 => "01100110",39335 => "00000010",39336 => "01010100",39337 => "00001100",39338 => "11100011",39339 => "10000111",39340 => "11000001",39341 => "11111010",39342 => "10111100",39343 => "00010000",39344 => "00011110",39345 => "10100000",39346 => "10110010",39347 => "10100110",39348 => "11110101",39349 => "01110111",39350 => "01111000",39351 => "01011101",39352 => "10100110",39353 => "10101100",39354 => "10001011",39355 => "10010011",39356 => "01111000",39357 => "10110111",39358 => "00111000",39359 => "00110001",39360 => "01111010",39361 => "01111111",39362 => "01110000",39363 => "00000010",39364 => "10111000",39365 => "01011011",39366 => "11101001",39367 => "01111010",39368 => "00011011",39369 => "00000101",39370 => "00011000",39371 => "01001110",39372 => "11001110",39373 => "01011100",39374 => "01010001",39375 => "10111010",39376 => "00110110",39377 => "11100010",39378 => "11101010",39379 => "10011111",39380 => "10011100",39381 => "11100111",39382 => "01000111",39383 => "11101110",39384 => "10000010",39385 => "11000100",39386 => "00100100",39387 => "10010000",39388 => "11001110",39389 => "01101101",39390 => "01100100",39391 => "00111001",39392 => "11100010",39393 => "00111110",39394 => "01000111",39395 => "01110010",39396 => "00001111",39397 => "00111110",39398 => "10111111",39399 => "00110001",39400 => "00111001",39401 => "01111000",39402 => "01000001",39403 => "10110110",39404 => "10011100",39405 => "00100010",39406 => "10101100",39407 => "01001010",39408 => "10001011",39409 => "11100010",39410 => "01100011",39411 => "11010010",39412 => "00010010",39413 => "01010001",39414 => "11101100",39415 => "11000001",39416 => "00101000",39417 => "10010000",39418 => "11011011",39419 => "11000100",39420 => "10010110",39421 => "00111000",39422 => "01101111",39423 => "10101010",39424 => "10000001",39425 => "00010010",39426 => "10011010",39427 => "01011001",39428 => "11010101",39429 => "11111010",39430 => "11010111",39431 => "00111010",39432 => "11110010",39433 => "10101010",39434 => "01101000",39435 => "11010011",39436 => "00101001",39437 => "10101010",39438 => "11010001",39439 => "11000011",39440 => "10111111",39441 => "10011111",39442 => "00011001",39443 => "01110001",39444 => "01000011",39445 => "00101001",39446 => "11011011",39447 => "00110111",39448 => "11001011",39449 => "01010010",39450 => "00000000",39451 => "10101011",39452 => "00011110",39453 => "11101110",39454 => "00001011",39455 => "11111110",39456 => "11111011",39457 => "01110101",39458 => "11000100",39459 => "11000011",39460 => "01110011",39461 => "00100111",39462 => "01011111",39463 => "10101000",39464 => "11000010",39465 => "11001110",39466 => "10111100",39467 => "00101110",39468 => "10111010",39469 => "10001010",39470 => "11001001",39471 => "01011110",39472 => "10111000",39473 => "00011101",39474 => "10011111",39475 => "01000100",39476 => "01100011",39477 => "11110101",39478 => "10000101",39479 => "00000100",39480 => "01110000",39481 => "11011100",39482 => "10001001",39483 => "01001101",39484 => "10010011",39485 => "11001000",39486 => "01110101",39487 => "01001001",39488 => "10100000",39489 => "11000010",39490 => "10011110",39491 => "11100110",39492 => "01111101",39493 => "10100010",39494 => "10001111",39495 => "00110011",39496 => "01010100",39497 => "10000101",39498 => "10101000",39499 => "10000010",39500 => "01001111",39501 => "00010011",39502 => "01101001",39503 => "10010110",39504 => "11011101",39505 => "11111010",39506 => "11000000",39507 => "00011011",39508 => "10001101",39509 => "11001100",39510 => "11010011",39511 => "10010000",39512 => "10011111",39513 => "10010001",39514 => "01111100",39515 => "01000001",39516 => "01101111",39517 => "00010010",39518 => "10001101",39519 => "01110111",39520 => "11110011",39521 => "01111001",39522 => "01011100",39523 => "11010101",39524 => "00001010",39525 => "01000111",39526 => "10000100",39527 => "01010000",39528 => "01010100",39529 => "11111110",39530 => "11010010",39531 => "01010100",39532 => "11101101",39533 => "01001101",39534 => "11000100",39535 => "00100101",39536 => "00110101",39537 => "11000000",39538 => "00111110",39539 => "00000011",39540 => "01111011",39541 => "00010010",39542 => "01100110",39543 => "00011100",39544 => "11000011",39545 => "00111010",39546 => "00101101",39547 => "00110101",39548 => "11110011",39549 => "11011100",39550 => "10001000",39551 => "10000100",39552 => "11111000",39553 => "10001011",39554 => "00110000",39555 => "10011110",39556 => "11101000",39557 => "01011111",39558 => "00100101",39559 => "10001011",39560 => "00011110",39561 => "00010101",39562 => "00000001",39563 => "01010010",39564 => "01010010",39565 => "11110011",39566 => "01011001",39567 => "10111100",39568 => "10110000",39569 => "10011110",39570 => "00100111",39571 => "10000101",39572 => "01011001",39573 => "00001110",39574 => "00000111",39575 => "10010110",39576 => "10101101",39577 => "10110110",39578 => "01111110",39579 => "00111000",39580 => "10110011",39581 => "00011001",39582 => "11110111",39583 => "11000101",39584 => "11101111",39585 => "11110100",39586 => "10011000",39587 => "10011010",39588 => "01101010",39589 => "10111111",39590 => "11111100",39591 => "10010101",39592 => "00011110",39593 => "10110010",39594 => "01101001",39595 => "11111001",39596 => "10001011",39597 => "11101100",39598 => "00010110",39599 => "11011100",39600 => "10110100",39601 => "11011010",39602 => "00000000",39603 => "11111101",39604 => "10110110",39605 => "01000110",39606 => "10110010",39607 => "10010110",39608 => "00000101",39609 => "10101110",39610 => "10010000",39611 => "10001010",39612 => "01110110",39613 => "00101101",39614 => "11111000",39615 => "10110010",39616 => "00110010",39617 => "11011101",39618 => "01011110",39619 => "01111111",39620 => "00011100",39621 => "01110101",39622 => "00000001",39623 => "10000101",39624 => "01111010",39625 => "01010011",39626 => "00011010",39627 => "10110001",39628 => "11100010",39629 => "10110000",39630 => "01110111",39631 => "11001100",39632 => "11111010",39633 => "01110010",39634 => "00101011",39635 => "00110111",39636 => "01010011",39637 => "10011100",39638 => "11101010",39639 => "01110100",39640 => "01000000",39641 => "00101010",39642 => "10101010",39643 => "11110000",39644 => "00110011",39645 => "01101001",39646 => "00100010",39647 => "10110100",39648 => "00010000",39649 => "10110110",39650 => "01001000",39651 => "10011011",39652 => "11000001",39653 => "00111110",39654 => "01110011",39655 => "10010011",39656 => "10110000",39657 => "00000011",39658 => "00011101",39659 => "10001110",39660 => "00000110",39661 => "00111000",39662 => "00101011",39663 => "00001110",39664 => "11001010",39665 => "00110111",39666 => "10100100",39667 => "00101110",39668 => "11010010",39669 => "10111111",39670 => "00010011",39671 => "01010110",39672 => "11110111",39673 => "11111011",39674 => "01001010",39675 => "10001101",39676 => "11100101",39677 => "00111110",39678 => "01111010",39679 => "11011111",39680 => "01000110",39681 => "01101100",39682 => "11010011",39683 => "10010000",39684 => "01011000",39685 => "01101110",39686 => "11100100",39687 => "10010000",39688 => "00110111",39689 => "00111110",39690 => "01100001",39691 => "10100010",39692 => "10000111",39693 => "11001001",39694 => "10001001",39695 => "11011000",39696 => "10000100",39697 => "01000000",39698 => "00100011",39699 => "10011110",39700 => "10000110",39701 => "01001010",39702 => "11101011",39703 => "10010100",39704 => "11010010",39705 => "11001100",39706 => "01101000",39707 => "10110110",39708 => "10100001",39709 => "00001000",39710 => "00110101",39711 => "01101110",39712 => "01111101",39713 => "11101010",39714 => "10001000",39715 => "10111100",39716 => "10000001",39717 => "11100000",39718 => "00011000",39719 => "01000111",39720 => "00111001",39721 => "11100110",39722 => "01010111",39723 => "11000101",39724 => "00001100",39725 => "10111010",39726 => "00000010",39727 => "11110110",39728 => "11011110",39729 => "00111101",39730 => "01001001",39731 => "11001011",39732 => "01011011",39733 => "10100001",39734 => "10101110",39735 => "00001110",39736 => "00111001",39737 => "11010001",39738 => "01000011",39739 => "10111100",39740 => "00101111",39741 => "00101001",39742 => "00010011",39743 => "11001001",39744 => "10100011",39745 => "01001001",39746 => "11100011",39747 => "01101100",39748 => "11100010",39749 => "00000001",39750 => "11110110",39751 => "01101101",39752 => "00100101",39753 => "10000000",39754 => "10100010",39755 => "11011101",39756 => "10111010",39757 => "00100000",39758 => "00101100",39759 => "10110001",39760 => "11111000",39761 => "11001010",39762 => "00001011",39763 => "00111011",39764 => "00111010",39765 => "01101110",39766 => "00101010",39767 => "01100011",39768 => "11100110",39769 => "00111111",39770 => "01011100",39771 => "00011111",39772 => "00000000",39773 => "10110111",39774 => "00011011",39775 => "01100111",39776 => "00110010",39777 => "01111110",39778 => "01010101",39779 => "10100001",39780 => "00110001",39781 => "11000100",39782 => "11011101",39783 => "01111110",39784 => "11100011",39785 => "00111011",39786 => "11100101",39787 => "00001010",39788 => "01111111",39789 => "01000111",39790 => "00011100",39791 => "10001101",39792 => "00100101",39793 => "01000110",39794 => "11101000",39795 => "01101101",39796 => "00001000",39797 => "10001110",39798 => "00100110",39799 => "10101000",39800 => "10111000",39801 => "00000101",39802 => "01100000",39803 => "00011111",39804 => "00000101",39805 => "10000100",39806 => "00111011",39807 => "01110110",39808 => "10011001",39809 => "01001110",39810 => "11001111",39811 => "10101010",39812 => "00001001",39813 => "11000010",39814 => "11110011",39815 => "11011011",39816 => "00000100",39817 => "11111101",39818 => "11101001",39819 => "01100011",39820 => "00000000",39821 => "00101010",39822 => "11010111",39823 => "11001010",39824 => "00101000",39825 => "11111001",39826 => "01011011",39827 => "00001111",39828 => "00100001",39829 => "11010011",39830 => "10001101",39831 => "11101010",39832 => "11000101",39833 => "10111001",39834 => "10101010",39835 => "00001111",39836 => "10011101",39837 => "00111011",39838 => "00110010",39839 => "00100110",39840 => "00010011",39841 => "00110111",39842 => "01011110",39843 => "01100011",39844 => "10101011",39845 => "00011001",39846 => "01100011",39847 => "00101000",39848 => "11011011",39849 => "11011110",39850 => "00111000",39851 => "01000111",39852 => "00010011",39853 => "11110100",39854 => "00111000",39855 => "00001110",39856 => "11100001",39857 => "00110001",39858 => "10011010",39859 => "01101111",39860 => "00011011",39861 => "01001100",39862 => "10010110",39863 => "01001011",39864 => "10000000",39865 => "01000001",39866 => "00100001",39867 => "00111000",39868 => "00100111",39869 => "01100101",39870 => "00110000",39871 => "00001001",39872 => "00000100",39873 => "10110001",39874 => "01101001",39875 => "00111111",39876 => "11111110",39877 => "11100000",39878 => "11001010",39879 => "11110011",39880 => "10100001",39881 => "10000101",39882 => "10110111",39883 => "11000111",39884 => "11110111",39885 => "01101101",39886 => "10110010",39887 => "11011111",39888 => "00011001",39889 => "10110101",39890 => "10010100",39891 => "00101001",39892 => "10101100",39893 => "11100101",39894 => "01111101",39895 => "10011100",39896 => "10110011",39897 => "10100010",39898 => "00110101",39899 => "10000000",39900 => "01101110",39901 => "10011000",39902 => "01001010",39903 => "00000111",39904 => "10101100",39905 => "01111110",39906 => "00001101",39907 => "01110111",39908 => "01010011",39909 => "00111010",39910 => "11100100",39911 => "01100110",39912 => "01101000",39913 => "11000100",39914 => "01101110",39915 => "01111001",39916 => "10111011",39917 => "01001011",39918 => "11100011",39919 => "00011001",39920 => "10000111",39921 => "11110010",39922 => "01000010",39923 => "10101010",39924 => "01100110",39925 => "00100111",39926 => "00111010",39927 => "00101101",39928 => "01010001",39929 => "01111110",39930 => "11100001",39931 => "00001001",39932 => "11000011",39933 => "11001011",39934 => "11100101",39935 => "00101001",39936 => "11101101",39937 => "01000010",39938 => "01000010",39939 => "01010001",39940 => "10111101",39941 => "10011111",39942 => "11000101",39943 => "11010110",39944 => "11110111",39945 => "10010101",39946 => "01110101",39947 => "11011000",39948 => "00101111",39949 => "10111101",39950 => "00010010",39951 => "00000000",39952 => "01110110",39953 => "11001000",39954 => "10000000",39955 => "01100010",39956 => "11000011",39957 => "10000011",39958 => "00111101",39959 => "11011111",39960 => "10000100",39961 => "10101110",39962 => "10101000",39963 => "11011001",39964 => "10011110",39965 => "11001011",39966 => "00111101",39967 => "11110010",39968 => "00100100",39969 => "00100111",39970 => "10010111",39971 => "11111111",39972 => "11000110",39973 => "10101100",39974 => "01001100",39975 => "11011001",39976 => "11111010",39977 => "10000100",39978 => "11100011",39979 => "10111000",39980 => "11001001",39981 => "10000101",39982 => "11100010",39983 => "10110110",39984 => "11101010",39985 => "11101100",39986 => "11101100",39987 => "01111110",39988 => "11000011",39989 => "11001001",39990 => "00111011",39991 => "11010110",39992 => "11011011",39993 => "01111000",39994 => "01110101",39995 => "00111101",39996 => "01101111",39997 => "01010101",39998 => "10100100",39999 => "10101010",40000 => "10110000",40001 => "01100001",40002 => "00100101",40003 => "01101111",40004 => "11001100",40005 => "11111000",40006 => "11010101",40007 => "10101110",40008 => "10000010",40009 => "01101100",40010 => "00011011",40011 => "10000001",40012 => "10110110",40013 => "11100100",40014 => "11110101",40015 => "11100110",40016 => "01101111",40017 => "11000110",40018 => "10011001",40019 => "11011111",40020 => "01111111",40021 => "11111001",40022 => "00111101",40023 => "11111111",40024 => "10011011",40025 => "00001001",40026 => "10011001",40027 => "10010110",40028 => "00000110",40029 => "01110011",40030 => "11010100",40031 => "11100011",40032 => "01111111",40033 => "11010010",40034 => "00011010",40035 => "00010101",40036 => "10110010",40037 => "10111110",40038 => "01100011",40039 => "10101000",40040 => "00111101",40041 => "10000100",40042 => "01001110",40043 => "00011011",40044 => "01111101",40045 => "10101010",40046 => "10010100",40047 => "00010000",40048 => "11010011",40049 => "01011111",40050 => "10100100",40051 => "11111110",40052 => "10000100",40053 => "10110101",40054 => "10100010",40055 => "00100101",40056 => "10101100",40057 => "11100100",40058 => "10100101",40059 => "00011100",40060 => "00010010",40061 => "11111100",40062 => "01101101",40063 => "01001110",40064 => "01010101",40065 => "10010110",40066 => "10010110",40067 => "00011001",40068 => "11010010",40069 => "10001010",40070 => "10001110",40071 => "00110110",40072 => "10101110",40073 => "11010101",40074 => "10010100",40075 => "01101101",40076 => "10111011",40077 => "11110100",40078 => "11010010",40079 => "01111001",40080 => "11000010",40081 => "11010101",40082 => "01101010",40083 => "01000110",40084 => "01110111",40085 => "11001000",40086 => "11111001",40087 => "10011011",40088 => "10011111",40089 => "01110001",40090 => "00111010",40091 => "00011101",40092 => "11100010",40093 => "11111110",40094 => "01000110",40095 => "00011000",40096 => "01011000",40097 => "00111010",40098 => "11010101",40099 => "10001101",40100 => "01111100",40101 => "10101001",40102 => "01011001",40103 => "01000001",40104 => "11100010",40105 => "00010110",40106 => "11101000",40107 => "01001011",40108 => "01101101",40109 => "01111001",40110 => "01101110",40111 => "11010001",40112 => "00011010",40113 => "11100000",40114 => "01100111",40115 => "10001001",40116 => "10010110",40117 => "00000110",40118 => "10110100",40119 => "00000000",40120 => "10000000",40121 => "11001000",40122 => "10111000",40123 => "01100110",40124 => "11000001",40125 => "10101101",40126 => "10001010",40127 => "01011110",40128 => "00101111",40129 => "00001001",40130 => "01001011",40131 => "00100000",40132 => "01011011",40133 => "00110110",40134 => "11101000",40135 => "01101010",40136 => "00110001",40137 => "10010110",40138 => "01000010",40139 => "00110100",40140 => "10011010",40141 => "01011100",40142 => "01100101",40143 => "11000111",40144 => "00011101",40145 => "00011101",40146 => "11010001",40147 => "00011000",40148 => "01111101",40149 => "00010101",40150 => "11000100",40151 => "10010010",40152 => "10110001",40153 => "10000011",40154 => "01001001",40155 => "01101111",40156 => "00111111",40157 => "01010100",40158 => "00001001",40159 => "01100110",40160 => "11110101",40161 => "00111011",40162 => "00100110",40163 => "11010100",40164 => "01111001",40165 => "10000010",40166 => "01110111",40167 => "00111010",40168 => "10000100",40169 => "00011100",40170 => "01000110",40171 => "11011111",40172 => "10001010",40173 => "01101010",40174 => "11111111",40175 => "00001101",40176 => "00000001",40177 => "01011010",40178 => "00010110",40179 => "11011100",40180 => "00010110",40181 => "00010000",40182 => "11110011",40183 => "10110011",40184 => "10111111",40185 => "01010111",40186 => "01111101",40187 => "01010001",40188 => "11010111",40189 => "10011001",40190 => "10010110",40191 => "10000010",40192 => "10001011",40193 => "11010100",40194 => "11100001",40195 => "11111111",40196 => "01100100",40197 => "11001011",40198 => "11000101",40199 => "01000110",40200 => "10110100",40201 => "10000100",40202 => "11101010",40203 => "10000001",40204 => "00100110",40205 => "01001001",40206 => "10111000",40207 => "11111011",40208 => "01011000",40209 => "00011111",40210 => "01000001",40211 => "11111111",40212 => "00011000",40213 => "01011100",40214 => "10001101",40215 => "10000100",40216 => "11101100",40217 => "10010101",40218 => "11000101",40219 => "10011110",40220 => "11011001",40221 => "01100100",40222 => "01100011",40223 => "01001111",40224 => "01011010",40225 => "01101010",40226 => "00000100",40227 => "11100001",40228 => "01010110",40229 => "10110101",40230 => "11111111",40231 => "00101110",40232 => "11111111",40233 => "10001100",40234 => "01000011",40235 => "10010110",40236 => "11001111",40237 => "11010010",40238 => "11100010",40239 => "11100101",40240 => "00111100",40241 => "11101010",40242 => "00000100",40243 => "00010111",40244 => "01100111",40245 => "00101101",40246 => "00110000",40247 => "01100011",40248 => "10111100",40249 => "11010100",40250 => "00101111",40251 => "11110001",40252 => "11100110",40253 => "10100110",40254 => "11100110",40255 => "11101100",40256 => "10111110",40257 => "01000110",40258 => "10111010",40259 => "00100110",40260 => "10001010",40261 => "11000010",40262 => "00010010",40263 => "11001100",40264 => "10110001",40265 => "01100011",40266 => "10110110",40267 => "01110010",40268 => "00010111",40269 => "01111110",40270 => "00110011",40271 => "10001101",40272 => "01111001",40273 => "00110101",40274 => "11101110",40275 => "00000000",40276 => "00010001",40277 => "00011011",40278 => "11101000",40279 => "01011100",40280 => "01011010",40281 => "00001011",40282 => "10101111",40283 => "01001101",40284 => "01001001",40285 => "00110101",40286 => "10100010",40287 => "11110001",40288 => "00101101",40289 => "10011101",40290 => "01001101",40291 => "10001010",40292 => "10111100",40293 => "01011101",40294 => "01100010",40295 => "10101001",40296 => "10111001",40297 => "10100000",40298 => "01000011",40299 => "10000010",40300 => "01010011",40301 => "01110000",40302 => "01111001",40303 => "10000101",40304 => "00010010",40305 => "01100000",40306 => "10001000",40307 => "01111010",40308 => "11100111",40309 => "10000101",40310 => "00010100",40311 => "00101100",40312 => "11010111",40313 => "00110010",40314 => "01100110",40315 => "00000100",40316 => "10010010",40317 => "10110111",40318 => "10010100",40319 => "00110011",40320 => "01000000",40321 => "01001110",40322 => "01101111",40323 => "11010101",40324 => "11110010",40325 => "01110010",40326 => "11101010",40327 => "01101000",40328 => "00010101",40329 => "11000100",40330 => "11000101",40331 => "10000000",40332 => "10110000",40333 => "00000000",40334 => "10101110",40335 => "01011010",40336 => "01110010",40337 => "10001001",40338 => "00111010",40339 => "00111111",40340 => "01011110",40341 => "11101100",40342 => "10010001",40343 => "10010110",40344 => "11101011",40345 => "01000111",40346 => "11000111",40347 => "01010110",40348 => "01101000",40349 => "10000001",40350 => "01111100",40351 => "00010110",40352 => "11010111",40353 => "11001101",40354 => "11100111",40355 => "10011001",40356 => "01100011",40357 => "01001111",40358 => "10001110",40359 => "10011111",40360 => "00110000",40361 => "00011011",40362 => "10010110",40363 => "11100010",40364 => "11111111",40365 => "11101101",40366 => "00110101",40367 => "00011011",40368 => "01101111",40369 => "00100111",40370 => "00001100",40371 => "01100100",40372 => "10100000",40373 => "10100001",40374 => "01001101",40375 => "01101000",40376 => "01111100",40377 => "00011000",40378 => "01000101",40379 => "01001111",40380 => "00111101",40381 => "00111111",40382 => "00111110",40383 => "11011000",40384 => "10110100",40385 => "10000111",40386 => "11100011",40387 => "01001111",40388 => "00111000",40389 => "10000110",40390 => "00010000",40391 => "00010100",40392 => "00011100",40393 => "01111000",40394 => "11111101",40395 => "10100011",40396 => "01001010",40397 => "10010110",40398 => "01101000",40399 => "01101111",40400 => "10100110",40401 => "10101011",40402 => "10000101",40403 => "11111010",40404 => "11110101",40405 => "01101101",40406 => "00100011",40407 => "10011001",40408 => "11101001",40409 => "00001100",40410 => "01101001",40411 => "10100111",40412 => "10101110",40413 => "01001110",40414 => "01001100",40415 => "11100111",40416 => "01110010",40417 => "00001110",40418 => "10110110",40419 => "11110010",40420 => "10101010",40421 => "01010011",40422 => "00001011",40423 => "01001001",40424 => "10100010",40425 => "00010000",40426 => "00111000",40427 => "11101100",40428 => "11010100",40429 => "11010011",40430 => "10000110",40431 => "01010011",40432 => "01111110",40433 => "01011101",40434 => "00111100",40435 => "10110001",40436 => "11101111",40437 => "00100001",40438 => "10011001",40439 => "00001000",40440 => "11001010",40441 => "00111000",40442 => "00001000",40443 => "11010110",40444 => "00110011",40445 => "10001110",40446 => "01011111",40447 => "00110010",40448 => "11101000",40449 => "01010110",40450 => "11000101",40451 => "11100101",40452 => "10101100",40453 => "10001010",40454 => "10001010",40455 => "10111111",40456 => "00010010",40457 => "10011001",40458 => "10011100",40459 => "00010011",40460 => "00011100",40461 => "00000000",40462 => "10011111",40463 => "10101101",40464 => "10100010",40465 => "10011010",40466 => "11011010",40467 => "11110110",40468 => "00111011",40469 => "00100010",40470 => "01010110",40471 => "11000110",40472 => "01101110",40473 => "01001101",40474 => "00001111",40475 => "11000001",40476 => "00011001",40477 => "00100000",40478 => "11111100",40479 => "11001110",40480 => "11000011",40481 => "10100111",40482 => "00001001",40483 => "01110110",40484 => "01111001",40485 => "11100100",40486 => "11111011",40487 => "01000101",40488 => "10100000",40489 => "01001011",40490 => "00101011",40491 => "11101100",40492 => "10001000",40493 => "00011011",40494 => "01101011",40495 => "10110001",40496 => "01001110",40497 => "01111000",40498 => "11010000",40499 => "00011010",40500 => "00001001",40501 => "00101001",40502 => "10111101",40503 => "00001111",40504 => "00011000",40505 => "10000001",40506 => "00101001",40507 => "00100000",40508 => "10101011",40509 => "00111110",40510 => "00101011",40511 => "01101111",40512 => "11110010",40513 => "11111111",40514 => "11001011",40515 => "01000011",40516 => "01010110",40517 => "11101001",40518 => "00001011",40519 => "00110111",40520 => "00000000",40521 => "10010100",40522 => "00000111",40523 => "00011000",40524 => "01000101",40525 => "10010001",40526 => "10011011",40527 => "11100110",40528 => "11110100",40529 => "00111101",40530 => "11101110",40531 => "10011011",40532 => "11110000",40533 => "11001100",40534 => "01000101",40535 => "10101000",40536 => "11001110",40537 => "10001110",40538 => "00001000",40539 => "00111100",40540 => "10111000",40541 => "10010101",40542 => "10101111",40543 => "10011101",40544 => "00011001",40545 => "11111011",40546 => "00111010",40547 => "01110100",40548 => "01001001",40549 => "10011011",40550 => "01000111",40551 => "00111111",40552 => "11010111",40553 => "00100000",40554 => "11011111",40555 => "00011101",40556 => "01101101",40557 => "00110001",40558 => "00000000",40559 => "01100010",40560 => "11110100",40561 => "11001000",40562 => "01101000",40563 => "01111011",40564 => "11110000",40565 => "11110001",40566 => "01110101",40567 => "01101100",40568 => "01111000",40569 => "01100011",40570 => "11011000",40571 => "00101111",40572 => "01001111",40573 => "00110011",40574 => "00011100",40575 => "10110110",40576 => "11011001",40577 => "11101100",40578 => "00001111",40579 => "10001010",40580 => "01000000",40581 => "10110110",40582 => "01010011",40583 => "11100111",40584 => "00111000",40585 => "10010000",40586 => "01010100",40587 => "00100101",40588 => "11001001",40589 => "00101010",40590 => "00101101",40591 => "11101011",40592 => "11111111",40593 => "10000000",40594 => "00101111",40595 => "01010110",40596 => "10110001",40597 => "01111010",40598 => "01100000",40599 => "00010000",40600 => "11100100",40601 => "11101100",40602 => "10100001",40603 => "10110101",40604 => "11011111",40605 => "11110010",40606 => "00000010",40607 => "10111001",40608 => "11111010",40609 => "00010011",40610 => "01010011",40611 => "00001100",40612 => "00101000",40613 => "11000110",40614 => "01110100",40615 => "00100011",40616 => "00101101",40617 => "01101000",40618 => "00001001",40619 => "01100001",40620 => "01000001",40621 => "11000001",40622 => "00101001",40623 => "10100011",40624 => "00110010",40625 => "01100111",40626 => "11000111",40627 => "11001101",40628 => "11010111",40629 => "10110101",40630 => "11011000",40631 => "11011110",40632 => "10011101",40633 => "11110011",40634 => "10000010",40635 => "11001001",40636 => "10010011",40637 => "00010110",40638 => "01000010",40639 => "11001100",40640 => "00011111",40641 => "01011010",40642 => "11010010",40643 => "01111001",40644 => "10101010",40645 => "11101010",40646 => "11010110",40647 => "11001010",40648 => "10100101",40649 => "10100010",40650 => "00001101",40651 => "00000101",40652 => "11010101",40653 => "10100000",40654 => "11110110",40655 => "10110110",40656 => "01111111",40657 => "00110010",40658 => "01010100",40659 => "01001111",40660 => "00101110",40661 => "00111101",40662 => "01000101",40663 => "11111001",40664 => "11010001",40665 => "01110000",40666 => "11111110",40667 => "11000100",40668 => "00110001",40669 => "00101000",40670 => "11110100",40671 => "11010001",40672 => "01000000",40673 => "00010110",40674 => "10011111",40675 => "01101010",40676 => "01100110",40677 => "11111111",40678 => "11111000",40679 => "01011011",40680 => "11101000",40681 => "11010111",40682 => "10110011",40683 => "11010011",40684 => "01000001",40685 => "01000101",40686 => "11101011",40687 => "00111101",40688 => "11100101",40689 => "11000000",40690 => "00001100",40691 => "00101100",40692 => "10110100",40693 => "10001011",40694 => "01110000",40695 => "00011111",40696 => "10011111",40697 => "10110101",40698 => "11100011",40699 => "01100111",40700 => "00111010",40701 => "01101001",40702 => "11110111",40703 => "00011100",40704 => "00010010",40705 => "00110100",40706 => "00001000",40707 => "11010101",40708 => "01110001",40709 => "01010100",40710 => "11110011",40711 => "10111100",40712 => "00101011",40713 => "01001010",40714 => "00100111",40715 => "01111110",40716 => "01000000",40717 => "11110100",40718 => "01010110",40719 => "10101001",40720 => "01001111",40721 => "11110001",40722 => "11001101",40723 => "11000010",40724 => "10010000",40725 => "10100111",40726 => "10010010",40727 => "01001110",40728 => "01011000",40729 => "11001001",40730 => "10001100",40731 => "01101110",40732 => "11110010",40733 => "01111100",40734 => "11010000",40735 => "10010010",40736 => "11101000",40737 => "00010101",40738 => "01010000",40739 => "01001101",40740 => "00011111",40741 => "11011101",40742 => "01001011",40743 => "10010101",40744 => "11101001",40745 => "11001000",40746 => "01100011",40747 => "10000101",40748 => "01001001",40749 => "10111100",40750 => "01111100",40751 => "01001000",40752 => "01111101",40753 => "01101001",40754 => "01000010",40755 => "10101001",40756 => "00111011",40757 => "00100001",40758 => "10011011",40759 => "01011001",40760 => "11011001",40761 => "01000100",40762 => "11011111",40763 => "11100110",40764 => "10110111",40765 => "01101100",40766 => "00011011",40767 => "01101011",40768 => "10110000",40769 => "10011010",40770 => "01110100",40771 => "10001000",40772 => "10010110",40773 => "01001000",40774 => "01010101",40775 => "01110011",40776 => "11011010",40777 => "00010100",40778 => "00010100",40779 => "10010001",40780 => "00001100",40781 => "10001100",40782 => "11100011",40783 => "11001001",40784 => "01111101",40785 => "10110100",40786 => "10100110",40787 => "11100010",40788 => "01010000",40789 => "01100100",40790 => "00101101",40791 => "01010011",40792 => "11110100",40793 => "11000000",40794 => "10010000",40795 => "11010100",40796 => "01100111",40797 => "00010001",40798 => "00110100",40799 => "01010110",40800 => "10001011",40801 => "00110100",40802 => "10100111",40803 => "10011100",40804 => "11110011",40805 => "11101100",40806 => "11101110",40807 => "10001001",40808 => "00110110",40809 => "10000100",40810 => "11011101",40811 => "10110100",40812 => "11110100",40813 => "10000001",40814 => "10100001",40815 => "10010001",40816 => "00000111",40817 => "00110011",40818 => "10001100",40819 => "10110111",40820 => "01110110",40821 => "01000011",40822 => "11001101",40823 => "01100001",40824 => "11010000",40825 => "10010010",40826 => "01001111",40827 => "00111001",40828 => "00011001",40829 => "10100000",40830 => "00000011",40831 => "11001000",40832 => "00110001",40833 => "10010010",40834 => "01101011",40835 => "10101100",40836 => "11111111",40837 => "01000110",40838 => "10000011",40839 => "00001110",40840 => "11100000",40841 => "01011011",40842 => "00000010",40843 => "10110101",40844 => "01100100",40845 => "01100010",40846 => "01001100",40847 => "01110011",40848 => "00010101",40849 => "11000110",40850 => "01001100",40851 => "01111100",40852 => "10000111",40853 => "00110011",40854 => "10111101",40855 => "00100011",40856 => "10010101",40857 => "01000110",40858 => "11111110",40859 => "11010001",40860 => "11000111",40861 => "10111100",40862 => "10001001",40863 => "01101111",40864 => "10011101",40865 => "01010100",40866 => "10100110",40867 => "01100101",40868 => "10101011",40869 => "11111111",40870 => "10010100",40871 => "01010111",40872 => "00001110",40873 => "00111100",40874 => "11011101",40875 => "01011010",40876 => "00111111",40877 => "11101001",40878 => "00101100",40879 => "01000100",40880 => "01011000",40881 => "00100101",40882 => "01000001",40883 => "10100011",40884 => "10000000",40885 => "11111000",40886 => "00100100",40887 => "10100001",40888 => "10111101",40889 => "11100111",40890 => "10000010",40891 => "01110001",40892 => "01000101",40893 => "11110000",40894 => "11000001",40895 => "00011110",40896 => "01100100",40897 => "01000111",40898 => "00011010",40899 => "11010000",40900 => "10110110",40901 => "01000000",40902 => "11100110",40903 => "11110000",40904 => "01010000",40905 => "11101110",40906 => "11110010",40907 => "11110011",40908 => "10000110",40909 => "10111000",40910 => "00010100",40911 => "01111101",40912 => "11011001",40913 => "01011001",40914 => "10101110",40915 => "01110100",40916 => "01110000",40917 => "11100000",40918 => "11100000",40919 => "01001011",40920 => "00010100",40921 => "00101110",40922 => "10111110",40923 => "11101010",40924 => "00100111",40925 => "11001011",40926 => "00100010",40927 => "11001011",40928 => "10000111",40929 => "11011010",40930 => "11110001",40931 => "00000000",40932 => "00100011",40933 => "00001000",40934 => "11101111",40935 => "01011011",40936 => "11101101",40937 => "00100010",40938 => "10111001",40939 => "01011100",40940 => "10011001",40941 => "01100100",40942 => "10000000",40943 => "10110010",40944 => "10111110",40945 => "11101111",40946 => "01010110",40947 => "00110101",40948 => "00001101",40949 => "01110010",40950 => "11001100",40951 => "01100101",40952 => "01010001",40953 => "01100100",40954 => "10000010",40955 => "11100100",40956 => "00011010",40957 => "01010010",40958 => "00011011",40959 => "11101000",40960 => "11111111",40961 => "00001110",40962 => "00100101",40963 => "10010000",40964 => "00110111",40965 => "11111101",40966 => "11100000",40967 => "00111100",40968 => "01100110",40969 => "01011100",40970 => "11110101",40971 => "10101101",40972 => "00101010",40973 => "10100011",40974 => "11111000",40975 => "11100101",40976 => "11101001",40977 => "11101110",40978 => "11101001",40979 => "10010101",40980 => "00100011",40981 => "00001001",40982 => "11010100",40983 => "00110010",40984 => "01010000",40985 => "00001001",40986 => "00111001",40987 => "11000110",40988 => "11001101",40989 => "01111111",40990 => "11110001",40991 => "00000100",40992 => "00101111",40993 => "00011111",40994 => "11111101",40995 => "00110110",40996 => "10101010",40997 => "11010001",40998 => "10101011",40999 => "00011100",41000 => "10100101",41001 => "00101011",41002 => "01000110",41003 => "11110001",41004 => "00000100",41005 => "01000001",41006 => "11101101",41007 => "01101111",41008 => "11010001",41009 => "11001111",41010 => "10000100",41011 => "10011110",41012 => "11101111",41013 => "11110011",41014 => "01011100",41015 => "01000011",41016 => "10010000",41017 => "01000101",41018 => "00111111",41019 => "10101000",41020 => "10011111",41021 => "11010010",41022 => "01111001",41023 => "01100100",41024 => "00010010",41025 => "10010011",41026 => "01001001",41027 => "10000011",41028 => "00010110",41029 => "00110100",41030 => "10000111",41031 => "01011010",41032 => "00001010",41033 => "01010011",41034 => "01110011",41035 => "10100011",41036 => "10010110",41037 => "00100100",41038 => "10010101",41039 => "01111010",41040 => "01100110",41041 => "11011101",41042 => "00001101",41043 => "10110101",41044 => "00011011",41045 => "10101011",41046 => "00001111",41047 => "00101010",41048 => "10101001",41049 => "00010001",41050 => "11010000",41051 => "01100111",41052 => "01100011",41053 => "01001001",41054 => "00011000",41055 => "01010001",41056 => "00001110",41057 => "11110100",41058 => "00011001",41059 => "00001000",41060 => "11000000",41061 => "11101011",41062 => "01111100",41063 => "10001011",41064 => "10001000",41065 => "10000000",41066 => "10010011",41067 => "10111001",41068 => "11001010",41069 => "00011011",41070 => "10011100",41071 => "11010001",41072 => "10001110",41073 => "10111110",41074 => "10001010",41075 => "00011011",41076 => "00010111",41077 => "00001000",41078 => "01111010",41079 => "01110011",41080 => "10111001",41081 => "10100110",41082 => "11000001",41083 => "01011001",41084 => "00011110",41085 => "11000011",41086 => "11011011",41087 => "00011110",41088 => "10000001",41089 => "11000110",41090 => "00111110",41091 => "01101011",41092 => "01010010",41093 => "00000010",41094 => "10111000",41095 => "01101100",41096 => "10001001",41097 => "10010110",41098 => "10111111",41099 => "10000001",41100 => "10111111",41101 => "11000111",41102 => "11011110",41103 => "10001110",41104 => "10101010",41105 => "01011001",41106 => "01100010",41107 => "11001110",41108 => "10101011",41109 => "00001010",41110 => "00011001",41111 => "00000100",41112 => "11110011",41113 => "01101000",41114 => "11110000",41115 => "00111110",41116 => "11100010",41117 => "10111101",41118 => "01011111",41119 => "00111000",41120 => "11101010",41121 => "10000000",41122 => "00110011",41123 => "11100101",41124 => "10101111",41125 => "00010001",41126 => "00001010",41127 => "10110001",41128 => "11001111",41129 => "01000101",41130 => "00110010",41131 => "00001111",41132 => "01110000",41133 => "01110101",41134 => "11100110",41135 => "00110001",41136 => "00000001",41137 => "01101001",41138 => "10100100",41139 => "11000011",41140 => "00100000",41141 => "00100110",41142 => "00101000",41143 => "10101001",41144 => "01001010",41145 => "00111111",41146 => "01010100",41147 => "11110111",41148 => "00010011",41149 => "00110011",41150 => "10011110",41151 => "01001010",41152 => "01010111",41153 => "10000011",41154 => "11100010",41155 => "10110001",41156 => "11101001",41157 => "00000011",41158 => "11110110",41159 => "10111011",41160 => "10001101",41161 => "11011111",41162 => "01000010",41163 => "11001000",41164 => "11011101",41165 => "01010000",41166 => "01000110",41167 => "10111011",41168 => "11101111",41169 => "00011000",41170 => "00111100",41171 => "11010100",41172 => "01101001",41173 => "01110000",41174 => "00100101",41175 => "11000000",41176 => "10111100",41177 => "01000111",41178 => "01011101",41179 => "11010000",41180 => "00111011",41181 => "00111010",41182 => "10001100",41183 => "01101101",41184 => "10010111",41185 => "11111010",41186 => "01000011",41187 => "10010001",41188 => "01000010",41189 => "10000010",41190 => "01111001",41191 => "00001100",41192 => "11101010",41193 => "00100011",41194 => "01011110",41195 => "10001001",41196 => "10000000",41197 => "11100100",41198 => "01110100",41199 => "00111100",41200 => "10000000",41201 => "00110010",41202 => "11010100",41203 => "11111010",41204 => "11010001",41205 => "10110101",41206 => "00101101",41207 => "01110011",41208 => "00110111",41209 => "01101100",41210 => "00001101",41211 => "01000010",41212 => "00011010",41213 => "00101100",41214 => "11001000",41215 => "11001001",41216 => "01011111",41217 => "11010010",41218 => "10101110",41219 => "01111001",41220 => "11100000",41221 => "01010011",41222 => "11110111",41223 => "10010111",41224 => "10011111",41225 => "11011101",41226 => "11010100",41227 => "11001000",41228 => "10111010",41229 => "01000111",41230 => "11010111",41231 => "11110011",41232 => "11111101",41233 => "01000110",41234 => "10000110",41235 => "00111100",41236 => "11111100",41237 => "01101111",41238 => "00100010",41239 => "01010111",41240 => "10010110",41241 => "00010011",41242 => "11111101",41243 => "00100111",41244 => "10111111",41245 => "00001110",41246 => "10010010",41247 => "00100010",41248 => "11111101",41249 => "00011000",41250 => "01101110",41251 => "00000010",41252 => "00110011",41253 => "01001010",41254 => "01011110",41255 => "10110010",41256 => "01001010",41257 => "11110010",41258 => "10011010",41259 => "01000111",41260 => "10101000",41261 => "11000111",41262 => "10111100",41263 => "11000011",41264 => "10000010",41265 => "10111001",41266 => "11011001",41267 => "01101110",41268 => "00110110",41269 => "11011111",41270 => "10110111",41271 => "10101011",41272 => "10010010",41273 => "10010000",41274 => "10000000",41275 => "10100111",41276 => "01101100",41277 => "11111111",41278 => "11111111",41279 => "10111011",41280 => "01001100",41281 => "00101001",41282 => "10101111",41283 => "10111010",41284 => "10001010",41285 => "00011010",41286 => "10000100",41287 => "10011000",41288 => "01000001",41289 => "11000000",41290 => "01001101",41291 => "10000100",41292 => "01000110",41293 => "01011010",41294 => "10111101",41295 => "11100001",41296 => "01110100",41297 => "01101001",41298 => "01100010",41299 => "01110101",41300 => "01110001",41301 => "11010101",41302 => "11101010",41303 => "01100011",41304 => "01001100",41305 => "10110111",41306 => "10111001",41307 => "11001001",41308 => "01100111",41309 => "01011100",41310 => "10000110",41311 => "01010000",41312 => "10001110",41313 => "01001110",41314 => "10000111",41315 => "10101001",41316 => "00011010",41317 => "10001111",41318 => "00011001",41319 => "00111110",41320 => "01001110",41321 => "10111110",41322 => "11011111",41323 => "11110111",41324 => "10101000",41325 => "01011000",41326 => "10101100",41327 => "01001100",41328 => "00101011",41329 => "00100001",41330 => "01101001",41331 => "11110111",41332 => "10000010",41333 => "10110011",41334 => "01100100",41335 => "01001101",41336 => "11111100",41337 => "00001100",41338 => "10110011",41339 => "01010011",41340 => "00001111",41341 => "10000000",41342 => "11101010",41343 => "11110101",41344 => "00111100",41345 => "10110100",41346 => "01001010",41347 => "11000100",41348 => "01000001",41349 => "01100100",41350 => "00010100",41351 => "11001010",41352 => "11110101",41353 => "01111000",41354 => "11111010",41355 => "00011111",41356 => "10001011",41357 => "00111111",41358 => "00000010",41359 => "00100011",41360 => "11100000",41361 => "00111110",41362 => "00110100",41363 => "10110101",41364 => "10100100",41365 => "10111101",41366 => "01000000",41367 => "11000110",41368 => "00100011",41369 => "01011111",41370 => "01110110",41371 => "10001100",41372 => "10011000",41373 => "11110011",41374 => "01111110",41375 => "11001100",41376 => "01110010",41377 => "01001011",41378 => "11101110",41379 => "00001010",41380 => "00111000",41381 => "11101001",41382 => "01110011",41383 => "01010111",41384 => "00011000",41385 => "11110101",41386 => "10100100",41387 => "01111100",41388 => "00101011",41389 => "11011010",41390 => "01100010",41391 => "00110111",41392 => "01011100",41393 => "00001110",41394 => "00111001",41395 => "10001100",41396 => "10100110",41397 => "10000000",41398 => "01111010",41399 => "11000010",41400 => "10001010",41401 => "00101001",41402 => "11101000",41403 => "01001110",41404 => "11011110",41405 => "11111010",41406 => "01100010",41407 => "10101001",41408 => "10000010",41409 => "10111011",41410 => "11001101",41411 => "00100000",41412 => "00110110",41413 => "01100101",41414 => "11011010",41415 => "00110000",41416 => "01110000",41417 => "00000101",41418 => "01101010",41419 => "01001010",41420 => "11100000",41421 => "01100111",41422 => "00000000",41423 => "11110100",41424 => "00001010",41425 => "01111101",41426 => "01011111",41427 => "01111001",41428 => "00110011",41429 => "10101100",41430 => "01111001",41431 => "10001011",41432 => "01000111",41433 => "00010000",41434 => "00001101",41435 => "10100001",41436 => "00111001",41437 => "00011000",41438 => "10001011",41439 => "01110110",41440 => "10101110",41441 => "10100100",41442 => "00010100",41443 => "00110100",41444 => "00010111",41445 => "00101110",41446 => "01111010",41447 => "10001000",41448 => "11011010",41449 => "00110001",41450 => "10010000",41451 => "10101011",41452 => "01100100",41453 => "10011001",41454 => "10111011",41455 => "10001111",41456 => "10011010",41457 => "01000000",41458 => "00101110",41459 => "00111001",41460 => "01101011",41461 => "00101100",41462 => "01110111",41463 => "01000100",41464 => "10100101",41465 => "10010110",41466 => "01010011",41467 => "10001010",41468 => "10010010",41469 => "00100101",41470 => "10000011",41471 => "01000101",41472 => "11000101",41473 => "00101000",41474 => "00111101",41475 => "10011000",41476 => "00101111",41477 => "10100011",41478 => "01110001",41479 => "00111001",41480 => "11001110",41481 => "00111011",41482 => "00111110",41483 => "10000110",41484 => "11010011",41485 => "10000010",41486 => "01111000",41487 => "01011000",41488 => "10101010",41489 => "00101001",41490 => "11100110",41491 => "01000110",41492 => "01110110",41493 => "11111101",41494 => "10110111",41495 => "11100011",41496 => "10101111",41497 => "11010100",41498 => "01000111",41499 => "01010000",41500 => "10001111",41501 => "00010010",41502 => "11010110",41503 => "01111101",41504 => "01010011",41505 => "11111111",41506 => "00001010",41507 => "11100001",41508 => "00100100",41509 => "01111111",41510 => "01111010",41511 => "01010101",41512 => "11100110",41513 => "00110101",41514 => "11100001",41515 => "11010000",41516 => "01010011",41517 => "11000100",41518 => "11110011",41519 => "11000101",41520 => "10110111",41521 => "10100011",41522 => "11011111",41523 => "00001111",41524 => "10110100",41525 => "10100110",41526 => "11110100",41527 => "00111000",41528 => "11011010",41529 => "11101000",41530 => "10110000",41531 => "00110001",41532 => "11111110",41533 => "10001110",41534 => "10110011",41535 => "11110011",41536 => "00010101",41537 => "00100101",41538 => "00110111",41539 => "10010100",41540 => "10010000",41541 => "11011010",41542 => "00111110",41543 => "10011001",41544 => "10001010",41545 => "10101001",41546 => "00011011",41547 => "11000101",41548 => "01001000",41549 => "10010100",41550 => "00100001",41551 => "00011110",41552 => "10101011",41553 => "00111000",41554 => "10010000",41555 => "01111011",41556 => "10001011",41557 => "11010101",41558 => "10101010",41559 => "01110001",41560 => "10101010",41561 => "01011111",41562 => "10111011",41563 => "01111101",41564 => "11101000",41565 => "11001010",41566 => "11011000",41567 => "11110100",41568 => "11101111",41569 => "11011110",41570 => "10011100",41571 => "00001010",41572 => "11010000",41573 => "00001001",41574 => "01110001",41575 => "00010010",41576 => "10110100",41577 => "10010001",41578 => "01101011",41579 => "11100010",41580 => "10000001",41581 => "01111101",41582 => "11100011",41583 => "10101101",41584 => "00111001",41585 => "01100100",41586 => "00110001",41587 => "00011011",41588 => "01010100",41589 => "01010111",41590 => "11101000",41591 => "01001111",41592 => "11001001",41593 => "00001010",41594 => "01000011",41595 => "11010110",41596 => "11110000",41597 => "01111101",41598 => "01000001",41599 => "10111001",41600 => "01010010",41601 => "10000000",41602 => "11100011",41603 => "01111010",41604 => "11001000",41605 => "10001110",41606 => "01011000",41607 => "11011101",41608 => "01100011",41609 => "00011001",41610 => "01100111",41611 => "11001111",41612 => "01100010",41613 => "01010000",41614 => "00110001",41615 => "01010010",41616 => "00110000",41617 => "11110001",41618 => "10111110",41619 => "10011001",41620 => "11101011",41621 => "11011000",41622 => "11010101",41623 => "10011111",41624 => "11000010",41625 => "11111100",41626 => "00011101",41627 => "00010110",41628 => "11111111",41629 => "01010100",41630 => "10110010",41631 => "10011101",41632 => "01011011",41633 => "00000110",41634 => "11110000",41635 => "00001001",41636 => "00100000",41637 => "00110100",41638 => "10111011",41639 => "01101000",41640 => "01010001",41641 => "10100000",41642 => "01010110",41643 => "01010110",41644 => "00110000",41645 => "00100101",41646 => "11001100",41647 => "10011000",41648 => "01011011",41649 => "10001001",41650 => "11111011",41651 => "10101000",41652 => "10001100",41653 => "01010011",41654 => "00001010",41655 => "00111111",41656 => "11011010",41657 => "11011100",41658 => "11110001",41659 => "01001100",41660 => "10110000",41661 => "10011101",41662 => "01011000",41663 => "10000111",41664 => "01110001",41665 => "10110101",41666 => "00110100",41667 => "11000000",41668 => "01011011",41669 => "10100001",41670 => "10011110",41671 => "00110010",41672 => "11110011",41673 => "11111111",41674 => "01000010",41675 => "01011100",41676 => "01001111",41677 => "11110010",41678 => "10111110",41679 => "10011100",41680 => "10101110",41681 => "10101111",41682 => "11001001",41683 => "11101100",41684 => "11101110",41685 => "01101111",41686 => "01001001",41687 => "00000011",41688 => "00010010",41689 => "00101110",41690 => "00101010",41691 => "01111100",41692 => "01010110",41693 => "00000100",41694 => "10001011",41695 => "10001101",41696 => "00001001",41697 => "01111001",41698 => "00001001",41699 => "10001110",41700 => "10000101",41701 => "11010101",41702 => "11011010",41703 => "10110111",41704 => "11111111",41705 => "10000010",41706 => "11011101",41707 => "11011111",41708 => "01000101",41709 => "00011111",41710 => "01001110",41711 => "00110011",41712 => "10100011",41713 => "00001110",41714 => "10110011",41715 => "00111010",41716 => "00010001",41717 => "01100111",41718 => "01010110",41719 => "10010110",41720 => "01010010",41721 => "11010101",41722 => "10001111",41723 => "11000010",41724 => "00101111",41725 => "00101101",41726 => "11011010",41727 => "00100010",41728 => "00010000",41729 => "01001111",41730 => "00110010",41731 => "00101001",41732 => "01011000",41733 => "11110100",41734 => "01011001",41735 => "11011001",41736 => "01011110",41737 => "01101101",41738 => "11110001",41739 => "11111011",41740 => "10111001",41741 => "10100011",41742 => "00100110",41743 => "01111101",41744 => "10111100",41745 => "00101110",41746 => "11100000",41747 => "11110101",41748 => "00111000",41749 => "00110101",41750 => "11001111",41751 => "10011001",41752 => "11000010",41753 => "11000001",41754 => "10010011",41755 => "00101010",41756 => "11010010",41757 => "11111110",41758 => "10001010",41759 => "00110100",41760 => "00110011",41761 => "11110010",41762 => "10001111",41763 => "10101000",41764 => "00100101",41765 => "11011000",41766 => "11001110",41767 => "00100110",41768 => "11011010",41769 => "01110011",41770 => "11001000",41771 => "01101010",41772 => "10010110",41773 => "00111011",41774 => "01001000",41775 => "11101101",41776 => "01111010",41777 => "11010111",41778 => "00010110",41779 => "11100100",41780 => "00100111",41781 => "10000110",41782 => "01010000",41783 => "11010100",41784 => "00011100",41785 => "01101010",41786 => "00001001",41787 => "00011110",41788 => "10111100",41789 => "10010000",41790 => "00110001",41791 => "11101001",41792 => "11100110",41793 => "00000011",41794 => "01011100",41795 => "00110110",41796 => "01100101",41797 => "11101100",41798 => "10100011",41799 => "01110110",41800 => "11011001",41801 => "00100110",41802 => "10100001",41803 => "00100101",41804 => "01010111",41805 => "11110001",41806 => "10100010",41807 => "10011000",41808 => "11100100",41809 => "01101000",41810 => "01100100",41811 => "10100110",41812 => "00111110",41813 => "11111101",41814 => "00110001",41815 => "10000110",41816 => "00001100",41817 => "11101000",41818 => "11111110",41819 => "00100111",41820 => "10011111",41821 => "11100111",41822 => "11000000",41823 => "10111011",41824 => "11010110",41825 => "01111010",41826 => "01111011",41827 => "11110110",41828 => "00111111",41829 => "11111110",41830 => "11101110",41831 => "10110010",41832 => "01011101",41833 => "00011110",41834 => "00100001",41835 => "11001111",41836 => "11001101",41837 => "00101010",41838 => "10110000",41839 => "11110010",41840 => "11001001",41841 => "01101000",41842 => "00101001",41843 => "00100010",41844 => "10000010",41845 => "01001011",41846 => "00000111",41847 => "01011110",41848 => "11001000",41849 => "11011110",41850 => "11101111",41851 => "11100000",41852 => "01101001",41853 => "10100010",41854 => "11111000",41855 => "11111110",41856 => "00010001",41857 => "01100001",41858 => "01011010",41859 => "11110110",41860 => "00100100",41861 => "11001110",41862 => "10011100",41863 => "00100111",41864 => "11110110",41865 => "00111101",41866 => "11001100",41867 => "01000101",41868 => "10010101",41869 => "00011101",41870 => "11111010",41871 => "01111100",41872 => "01010100",41873 => "00010101",41874 => "01001001",41875 => "11111011",41876 => "00011000",41877 => "10110111",41878 => "01001110",41879 => "11101101",41880 => "10100110",41881 => "00101110",41882 => "00110011",41883 => "10010000",41884 => "11010011",41885 => "00010101",41886 => "00001001",41887 => "00101011",41888 => "01110111",41889 => "01111111",41890 => "10000011",41891 => "01101010",41892 => "10000110",41893 => "01000111",41894 => "11111011",41895 => "01000010",41896 => "11001000",41897 => "00011011",41898 => "10101110",41899 => "01011110",41900 => "00111011",41901 => "10100101",41902 => "00100101",41903 => "01011000",41904 => "11011110",41905 => "10011010",41906 => "10101001",41907 => "11100000",41908 => "01110010",41909 => "11010010",41910 => "10010110",41911 => "10001101",41912 => "01010101",41913 => "00010010",41914 => "00110001",41915 => "10100110",41916 => "10000011",41917 => "10011011",41918 => "01110010",41919 => "10011111",41920 => "01001111",41921 => "11101001",41922 => "00011100",41923 => "01010011",41924 => "11110111",41925 => "11000011",41926 => "00110111",41927 => "11110010",41928 => "11111010",41929 => "11100001",41930 => "10001110",41931 => "01001000",41932 => "01010101",41933 => "00110011",41934 => "10111010",41935 => "01010010",41936 => "01000110",41937 => "11111100",41938 => "00101111",41939 => "10110111",41940 => "00000001",41941 => "00110011",41942 => "11000000",41943 => "01010111",41944 => "01110001",41945 => "10010011",41946 => "00001110",41947 => "10110001",41948 => "10001010",41949 => "01110000",41950 => "01011101",41951 => "11011000",41952 => "10001101",41953 => "01101000",41954 => "11000010",41955 => "01001000",41956 => "01000011",41957 => "10110111",41958 => "00110100",41959 => "10000011",41960 => "01001100",41961 => "11101111",41962 => "10101001",41963 => "11101000",41964 => "01011100",41965 => "10101001",41966 => "11111101",41967 => "10100101",41968 => "01101010",41969 => "01001100",41970 => "01110011",41971 => "10001000",41972 => "10101011",41973 => "00010111",41974 => "01011100",41975 => "11101001",41976 => "10011011",41977 => "11100011",41978 => "11100111",41979 => "10011110",41980 => "10011100",41981 => "01001101",41982 => "00001001",41983 => "01000111",41984 => "10000111",41985 => "10011001",41986 => "10111111",41987 => "00001110",41988 => "01100001",41989 => "01011010",41990 => "00001110",41991 => "10110001",41992 => "01001010",41993 => "00000011",41994 => "10011111",41995 => "01101001",41996 => "00100110",41997 => "01110100",41998 => "10111010",41999 => "11100100",42000 => "10001011",42001 => "00101000",42002 => "11111110",42003 => "01110010",42004 => "11101000",42005 => "11100100",42006 => "11011111",42007 => "10011101",42008 => "10001010",42009 => "00001011",42010 => "11101001",42011 => "00110011",42012 => "00110010",42013 => "00110011",42014 => "11101101",42015 => "00000101",42016 => "01010111",42017 => "01100011",42018 => "00100010",42019 => "10001110",42020 => "01000010",42021 => "11000000",42022 => "01010101",42023 => "01000100",42024 => "11010100",42025 => "00100110",42026 => "11111011",42027 => "00011010",42028 => "01110100",42029 => "01101110",42030 => "10110100",42031 => "01100001",42032 => "11111010",42033 => "10101010",42034 => "10000001",42035 => "01010111",42036 => "11000010",42037 => "01011001",42038 => "00000101",42039 => "01100011",42040 => "10000001",42041 => "11000011",42042 => "11010010",42043 => "11111001",42044 => "00100010",42045 => "11111001",42046 => "10111001",42047 => "10101110",42048 => "10010011",42049 => "00111011",42050 => "00110000",42051 => "00011111",42052 => "01001001",42053 => "00011101",42054 => "00100111",42055 => "00011100",42056 => "00001111",42057 => "01111101",42058 => "10110001",42059 => "11010011",42060 => "11111111",42061 => "01101011",42062 => "01111100",42063 => "11111001",42064 => "11101001",42065 => "11100111",42066 => "11011110",42067 => "01110110",42068 => "10111010",42069 => "11010001",42070 => "11110110",42071 => "01111101",42072 => "10100000",42073 => "01010111",42074 => "01000010",42075 => "01110101",42076 => "00100100",42077 => "11001100",42078 => "00101111",42079 => "01111001",42080 => "10101000",42081 => "10101100",42082 => "11101000",42083 => "11010011",42084 => "01011010",42085 => "10011000",42086 => "11010011",42087 => "10010100",42088 => "01110101",42089 => "10011101",42090 => "00001111",42091 => "10100110",42092 => "01000110",42093 => "00110001",42094 => "01000111",42095 => "00110100",42096 => "00101011",42097 => "00010100",42098 => "10110010",42099 => "01100000",42100 => "11100010",42101 => "11001010",42102 => "00001001",42103 => "00011001",42104 => "00111011",42105 => "10001011",42106 => "01001101",42107 => "01011001",42108 => "11011011",42109 => "00001011",42110 => "01001100",42111 => "00101101",42112 => "10100010",42113 => "00111111",42114 => "00011110",42115 => "00001010",42116 => "10000001",42117 => "10000100",42118 => "01001100",42119 => "10101010",42120 => "01110010",42121 => "00000100",42122 => "00000110",42123 => "00000101",42124 => "01001001",42125 => "01001100",42126 => "00001000",42127 => "11000011",42128 => "11001111",42129 => "11001100",42130 => "00001111",42131 => "00010011",42132 => "00101101",42133 => "00001000",42134 => "00000001",42135 => "11010010",42136 => "01010101",42137 => "10111001",42138 => "00001001",42139 => "11111011",42140 => "11001110",42141 => "10000011",42142 => "10001010",42143 => "01000100",42144 => "01110101",42145 => "01110010",42146 => "10000011",42147 => "10011010",42148 => "00000110",42149 => "10110001",42150 => "01000011",42151 => "11000101",42152 => "11110110",42153 => "10110101",42154 => "00100000",42155 => "11101010",42156 => "01111011",42157 => "11010101",42158 => "01001001",42159 => "01011011",42160 => "10100101",42161 => "11110000",42162 => "10011100",42163 => "11001010",42164 => "00101110",42165 => "01100011",42166 => "01010010",42167 => "01001100",42168 => "10100110",42169 => "00011011",42170 => "00011000",42171 => "11100110",42172 => "11100001",42173 => "01101001",42174 => "00010000",42175 => "01100110",42176 => "10001010",42177 => "10111011",42178 => "11101001",42179 => "11011000",42180 => "10000101",42181 => "10111011",42182 => "11101110",42183 => "10010100",42184 => "00000000",42185 => "11000001",42186 => "11110011",42187 => "00110001",42188 => "11111110",42189 => "11011100",42190 => "01010011",42191 => "11011111",42192 => "00101010",42193 => "00010101",42194 => "01101100",42195 => "11000111",42196 => "10111101",42197 => "10100000",42198 => "00110011",42199 => "10111110",42200 => "10011101",42201 => "10000010",42202 => "10000011",42203 => "01001011",42204 => "10111010",42205 => "00111011",42206 => "00101000",42207 => "00110100",42208 => "10101110",42209 => "00001001",42210 => "01110010",42211 => "11111010",42212 => "00001001",42213 => "00000011",42214 => "11110010",42215 => "11100001",42216 => "10100101",42217 => "10110101",42218 => "11001110",42219 => "01111011",42220 => "00110010",42221 => "11000110",42222 => "11000101",42223 => "11100000",42224 => "11101000",42225 => "00010100",42226 => "10101111",42227 => "10000101",42228 => "01111111",42229 => "11011111",42230 => "01110100",42231 => "01000110",42232 => "01010001",42233 => "00101000",42234 => "01111011",42235 => "11100000",42236 => "10110000",42237 => "01011001",42238 => "00011100",42239 => "10010110",42240 => "10100001",42241 => "10100010",42242 => "01111011",42243 => "11110011",42244 => "10100000",42245 => "00110100",42246 => "11011011",42247 => "00011010",42248 => "11011010",42249 => "10100100",42250 => "10011010",42251 => "01100101",42252 => "01010110",42253 => "10001001",42254 => "01010111",42255 => "01110111",42256 => "11110101",42257 => "01100000",42258 => "10011001",42259 => "10111101",42260 => "00001000",42261 => "10001110",42262 => "00001100",42263 => "00010001",42264 => "11110001",42265 => "11011011",42266 => "01010100",42267 => "10100100",42268 => "00101011",42269 => "01110111",42270 => "01111010",42271 => "00101110",42272 => "10010010",42273 => "11100010",42274 => "10100001",42275 => "00111001",42276 => "10011001",42277 => "10001110",42278 => "00001101",42279 => "10010111",42280 => "00000110",42281 => "11101110",42282 => "01010110",42283 => "10000011",42284 => "00100010",42285 => "01011110",42286 => "00100100",42287 => "00100100",42288 => "01101000",42289 => "11110101",42290 => "10000010",42291 => "01001001",42292 => "00111100",42293 => "01101110",42294 => "01101010",42295 => "01010010",42296 => "00000101",42297 => "11100010",42298 => "01011010",42299 => "00101011",42300 => "11001100",42301 => "11011111",42302 => "00110010",42303 => "01101010",42304 => "11000010",42305 => "00100100",42306 => "11010111",42307 => "01011011",42308 => "10100111",42309 => "01011110",42310 => "01000010",42311 => "10000000",42312 => "10111101",42313 => "10010011",42314 => "00000101",42315 => "00011101",42316 => "11000000",42317 => "11101000",42318 => "01010100",42319 => "01110110",42320 => "00101001",42321 => "11011001",42322 => "11110011",42323 => "00000000",42324 => "11011010",42325 => "00110001",42326 => "00011010",42327 => "00001100",42328 => "01100101",42329 => "01000101",42330 => "00110001",42331 => "11110000",42332 => "10100110",42333 => "11001100",42334 => "11110011",42335 => "01001010",42336 => "10100100",42337 => "01000101",42338 => "00011100",42339 => "01110010",42340 => "11100110",42341 => "10010010",42342 => "01000110",42343 => "11011000",42344 => "10100000",42345 => "01111000",42346 => "11010100",42347 => "00011011",42348 => "11111101",42349 => "00110011",42350 => "00000111",42351 => "10101101",42352 => "11001001",42353 => "00010100",42354 => "00110101",42355 => "00001111",42356 => "10101110",42357 => "10100101",42358 => "11000100",42359 => "00100101",42360 => "11101100",42361 => "01011000",42362 => "11011011",42363 => "11111000",42364 => "01010100",42365 => "11001110",42366 => "01101101",42367 => "11000110",42368 => "11001001",42369 => "11111001",42370 => "11001100",42371 => "10001110",42372 => "11000111",42373 => "10011001",42374 => "00111011",42375 => "01101110",42376 => "11100100",42377 => "00000011",42378 => "11001001",42379 => "11101110",42380 => "10100101",42381 => "00010010",42382 => "11100110",42383 => "01101111",42384 => "00010100",42385 => "10111001",42386 => "10101110",42387 => "01001010",42388 => "01100111",42389 => "00100000",42390 => "11010101",42391 => "00011101",42392 => "11100101",42393 => "00111011",42394 => "10011001",42395 => "01111110",42396 => "01101000",42397 => "01100101",42398 => "10001111",42399 => "00111100",42400 => "11000100",42401 => "00110011",42402 => "11010000",42403 => "01110111",42404 => "11011010",42405 => "11111011",42406 => "11011101",42407 => "00101011",42408 => "00100011",42409 => "00000101",42410 => "11111010",42411 => "01000100",42412 => "10011011",42413 => "00000000",42414 => "11011100",42415 => "11110111",42416 => "11000111",42417 => "10001001",42418 => "11111110",42419 => "01111011",42420 => "01110000",42421 => "00100000",42422 => "11100101",42423 => "01110111",42424 => "00001110",42425 => "01010011",42426 => "01100101",42427 => "10101110",42428 => "10000110",42429 => "00101111",42430 => "01111101",42431 => "01110000",42432 => "01111100",42433 => "10001111",42434 => "10001110",42435 => "11000000",42436 => "11100111",42437 => "10001010",42438 => "01111010",42439 => "11110010",42440 => "01100111",42441 => "01110100",42442 => "11000001",42443 => "01010011",42444 => "01110100",42445 => "11000011",42446 => "10011111",42447 => "10000000",42448 => "11000100",42449 => "00110001",42450 => "10001000",42451 => "00000101",42452 => "01110110",42453 => "11000001",42454 => "00000011",42455 => "11100000",42456 => "11011000",42457 => "00101000",42458 => "01101011",42459 => "01100001",42460 => "00010100",42461 => "01110010",42462 => "10101011",42463 => "10000110",42464 => "01100010",42465 => "01010110",42466 => "00011111",42467 => "10001011",42468 => "00111110",42469 => "10110011",42470 => "00100001",42471 => "01100001",42472 => "01001011",42473 => "11011110",42474 => "10111010",42475 => "11101111",42476 => "11001100",42477 => "01000011",42478 => "00110111",42479 => "00010101",42480 => "01011001",42481 => "11001101",42482 => "00011100",42483 => "00101011",42484 => "00111110",42485 => "11111011",42486 => "10001011",42487 => "01001001",42488 => "00001111",42489 => "10111110",42490 => "00010010",42491 => "01011001",42492 => "01111000",42493 => "01101100",42494 => "00101100",42495 => "01110110",42496 => "00010011",42497 => "00011011",42498 => "01001010",42499 => "10001011",42500 => "11000111",42501 => "10010010",42502 => "11100000",42503 => "10111100",42504 => "01110101",42505 => "01000010",42506 => "00001110",42507 => "01111101",42508 => "01111111",42509 => "11010100",42510 => "10111100",42511 => "01111010",42512 => "01010000",42513 => "01010111",42514 => "11111101",42515 => "10011100",42516 => "11111111",42517 => "00000101",42518 => "00011011",42519 => "00000101",42520 => "10111100",42521 => "10000101",42522 => "10010010",42523 => "11100101",42524 => "00011011",42525 => "11010001",42526 => "01010011",42527 => "10110101",42528 => "11100011",42529 => "01110110",42530 => "00000001",42531 => "00001001",42532 => "00101001",42533 => "00000011",42534 => "00010110",42535 => "11100011",42536 => "01011001",42537 => "00111110",42538 => "10011111",42539 => "01100011",42540 => "00100111",42541 => "01010010",42542 => "01100010",42543 => "10010000",42544 => "11100011",42545 => "01000110",42546 => "11010111",42547 => "00111011",42548 => "10100001",42549 => "11001100",42550 => "10011010",42551 => "01110110",42552 => "01101010",42553 => "10011010",42554 => "01001010",42555 => "00010000",42556 => "00011011",42557 => "01001001",42558 => "10101001",42559 => "00110000",42560 => "01111010",42561 => "10001011",42562 => "00101000",42563 => "11010011",42564 => "11001111",42565 => "00001110",42566 => "11101001",42567 => "01101011",42568 => "11111110",42569 => "11100100",42570 => "10001011",42571 => "10100011",42572 => "11100101",42573 => "11000101",42574 => "11010010",42575 => "00011100",42576 => "00111010",42577 => "10110000",42578 => "11100001",42579 => "10111011",42580 => "01010100",42581 => "10010011",42582 => "11001000",42583 => "00010000",42584 => "01010101",42585 => "11010010",42586 => "01110111",42587 => "10001110",42588 => "00101010",42589 => "11001010",42590 => "01011010",42591 => "11100101",42592 => "10001100",42593 => "01110011",42594 => "11111110",42595 => "10000000",42596 => "01111001",42597 => "10111000",42598 => "10011011",42599 => "11101011",42600 => "11111110",42601 => "11101000",42602 => "01101010",42603 => "10100011",42604 => "10011011",42605 => "11110111",42606 => "11111101",42607 => "11010110",42608 => "01011001",42609 => "11101000",42610 => "10111100",42611 => "11010010",42612 => "01110011",42613 => "10101001",42614 => "00111101",42615 => "01110101",42616 => "11010111",42617 => "10011100",42618 => "10101110",42619 => "10010000",42620 => "10111111",42621 => "11000011",42622 => "01101000",42623 => "01110010",42624 => "00100110",42625 => "00111001",42626 => "00010011",42627 => "11000010",42628 => "01110100",42629 => "10100010",42630 => "01110011",42631 => "11101011",42632 => "00101010",42633 => "11001100",42634 => "11101001",42635 => "00001101",42636 => "11110001",42637 => "01011101",42638 => "11010000",42639 => "11111110",42640 => "01000001",42641 => "11101111",42642 => "01100000",42643 => "11010111",42644 => "11110100",42645 => "00010101",42646 => "01000011",42647 => "11100100",42648 => "01100100",42649 => "10010000",42650 => "11011000",42651 => "01011110",42652 => "10011000",42653 => "00110010",42654 => "01010101",42655 => "00010001",42656 => "00110111",42657 => "00101011",42658 => "01000001",42659 => "00110110",42660 => "01111111",42661 => "00110000",42662 => "01010000",42663 => "00101011",42664 => "00101011",42665 => "10000001",42666 => "00000011",42667 => "00111100",42668 => "01101000",42669 => "00100101",42670 => "01010100",42671 => "00100010",42672 => "01011111",42673 => "01000011",42674 => "00000101",42675 => "00001000",42676 => "10110010",42677 => "11100111",42678 => "10100000",42679 => "00010010",42680 => "01111000",42681 => "01110001",42682 => "01111001",42683 => "00010011",42684 => "01110001",42685 => "10011111",42686 => "11000001",42687 => "01010101",42688 => "01000101",42689 => "00000101",42690 => "10010111",42691 => "00001000",42692 => "00011010",42693 => "01011010",42694 => "01101100",42695 => "00010000",42696 => "01111010",42697 => "01100100",42698 => "10010110",42699 => "00111111",42700 => "11010010",42701 => "10011110",42702 => "10101001",42703 => "01011011",42704 => "00100101",42705 => "11101100",42706 => "01001101",42707 => "10101101",42708 => "00111100",42709 => "10110011",42710 => "00001100",42711 => "10001011",42712 => "11011101",42713 => "00000011",42714 => "10100100",42715 => "11110001",42716 => "11110011",42717 => "10110000",42718 => "01000110",42719 => "01010011",42720 => "10111001",42721 => "10101101",42722 => "11111111",42723 => "10011001",42724 => "10111010",42725 => "01100011",42726 => "11110001",42727 => "00110100",42728 => "01001001",42729 => "10111111",42730 => "00011011",42731 => "00110001",42732 => "00111111",42733 => "01111011",42734 => "00010000",42735 => "00001101",42736 => "01000011",42737 => "01101100",42738 => "11111010",42739 => "01011010",42740 => "11100111",42741 => "11110001",42742 => "10100100",42743 => "01001111",42744 => "00100100",42745 => "11100100",42746 => "11010111",42747 => "01010111",42748 => "01010000",42749 => "10001000",42750 => "00010110",42751 => "10101011",42752 => "00101001",42753 => "01111101",42754 => "01101111",42755 => "10111000",42756 => "01011001",42757 => "01010011",42758 => "00011000",42759 => "11111010",42760 => "10010100",42761 => "00011100",42762 => "11011100",42763 => "10101001",42764 => "00100001",42765 => "01101011",42766 => "01011110",42767 => "11000101",42768 => "11100100",42769 => "01111010",42770 => "01100101",42771 => "10101001",42772 => "01001000",42773 => "00111010",42774 => "10001100",42775 => "11011101",42776 => "00001001",42777 => "01001011",42778 => "01001110",42779 => "11111011",42780 => "10111001",42781 => "00101111",42782 => "01010011",42783 => "01101111",42784 => "10000100",42785 => "11010000",42786 => "10100000",42787 => "00110100",42788 => "10011110",42789 => "11000000",42790 => "11010111",42791 => "01001100",42792 => "01010100",42793 => "00000010",42794 => "11111011",42795 => "10101111",42796 => "11100000",42797 => "01111111",42798 => "11010110",42799 => "10011100",42800 => "10001001",42801 => "11010100",42802 => "11110001",42803 => "01101110",42804 => "00001111",42805 => "10111110",42806 => "00011001",42807 => "00100110",42808 => "10111110",42809 => "01001100",42810 => "01011110",42811 => "11110010",42812 => "11111010",42813 => "00111000",42814 => "01110101",42815 => "00101110",42816 => "01001101",42817 => "11100101",42818 => "10100001",42819 => "00011111",42820 => "01111001",42821 => "01100100",42822 => "00110000",42823 => "00010111",42824 => "00101001",42825 => "11000010",42826 => "01011110",42827 => "00001011",42828 => "10101010",42829 => "00110111",42830 => "00000110",42831 => "11011010",42832 => "11110011",42833 => "10101000",42834 => "00001011",42835 => "10111001",42836 => "11001111",42837 => "11000111",42838 => "10101001",42839 => "01010111",42840 => "11101101",42841 => "10011000",42842 => "00000001",42843 => "11010001",42844 => "10100101",42845 => "11111001",42846 => "10001000",42847 => "11011010",42848 => "11010000",42849 => "10010110",42850 => "01001111",42851 => "00001111",42852 => "00000000",42853 => "10011111",42854 => "01010110",42855 => "00111111",42856 => "01101101",42857 => "10001110",42858 => "01101010",42859 => "00010111",42860 => "01100101",42861 => "11011011",42862 => "01101011",42863 => "10101110",42864 => "10011001",42865 => "10001111",42866 => "10011110",42867 => "11100101",42868 => "01110010",42869 => "01000001",42870 => "10011111",42871 => "00000101",42872 => "10010000",42873 => "10000101",42874 => "00101011",42875 => "10001101",42876 => "01110010",42877 => "01110011",42878 => "10101101",42879 => "01001010",42880 => "01010110",42881 => "00001101",42882 => "01100100",42883 => "11110001",42884 => "00001111",42885 => "11110010",42886 => "11110101",42887 => "00100011",42888 => "10001101",42889 => "11001100",42890 => "01100110",42891 => "10101111",42892 => "10100111",42893 => "00111010",42894 => "10011001",42895 => "01110000",42896 => "11110101",42897 => "00011110",42898 => "01101100",42899 => "11010001",42900 => "00110001",42901 => "00000010",42902 => "10100010",42903 => "10101110",42904 => "00111101",42905 => "11001000",42906 => "00111100",42907 => "00010100",42908 => "11010011",42909 => "10100000",42910 => "01111000",42911 => "01000110",42912 => "00100110",42913 => "00011101",42914 => "10101010",42915 => "01100101",42916 => "10010001",42917 => "01110111",42918 => "01110001",42919 => "10100000",42920 => "11000000",42921 => "10101011",42922 => "10100100",42923 => "11011100",42924 => "11011110",42925 => "01000100",42926 => "01110000",42927 => "01100101",42928 => "11110100",42929 => "01111110",42930 => "11100100",42931 => "10111001",42932 => "00111000",42933 => "00010111",42934 => "01011110",42935 => "00101010",42936 => "00010010",42937 => "10010001",42938 => "00011011",42939 => "00101010",42940 => "00000001",42941 => "00111111",42942 => "11101011",42943 => "11001110",42944 => "11000000",42945 => "00101110",42946 => "01001110",42947 => "00011011",42948 => "10010000",42949 => "11111111",42950 => "01100000",42951 => "00001001",42952 => "11011101",42953 => "10001001",42954 => "01111000",42955 => "11000010",42956 => "10101100",42957 => "10011111",42958 => "11000110",42959 => "00100100",42960 => "00010110",42961 => "01100111",42962 => "00000010",42963 => "00001110",42964 => "01110111",42965 => "01010111",42966 => "01110011",42967 => "11010001",42968 => "01010100",42969 => "10000010",42970 => "10100101",42971 => "00010001",42972 => "01101001",42973 => "00110011",42974 => "00101011",42975 => "10101101",42976 => "10111110",42977 => "10000111",42978 => "00010001",42979 => "00111100",42980 => "01000001",42981 => "11000110",42982 => "00010001",42983 => "10011000",42984 => "00100010",42985 => "01110110",42986 => "01001011",42987 => "01001110",42988 => "11111110",42989 => "10000110",42990 => "11110000",42991 => "00111110",42992 => "01001001",42993 => "10000001",42994 => "10001100",42995 => "11101110",42996 => "11101000",42997 => "01000111",42998 => "10010100",42999 => "11100001",43000 => "10010010",43001 => "10100101",43002 => "10001100",43003 => "00000001",43004 => "01111010",43005 => "10001010",43006 => "10000000",43007 => "11011011",43008 => "10111000",43009 => "11011111",43010 => "00000101",43011 => "10111111",43012 => "11101001",43013 => "11111101",43014 => "10011000",43015 => "01010010",43016 => "10010101",43017 => "11011111",43018 => "10011011",43019 => "01010101",43020 => "11110101",43021 => "00111110",43022 => "10100001",43023 => "11100000",43024 => "01100100",43025 => "11100010",43026 => "01000101",43027 => "01010100",43028 => "10111001",43029 => "10110001",43030 => "11001011",43031 => "11111001",43032 => "00000000",43033 => "11011001",43034 => "10111110",43035 => "01010000",43036 => "01010111",43037 => "11000010",43038 => "01011110",43039 => "00101010",43040 => "10110010",43041 => "10001000",43042 => "10000111",43043 => "11011110",43044 => "10011000",43045 => "11100110",43046 => "10110000",43047 => "00011010",43048 => "01000100",43049 => "01010001",43050 => "01011101",43051 => "11011111",43052 => "00100000",43053 => "00111110",43054 => "10100000",43055 => "01010100",43056 => "00100111",43057 => "00111000",43058 => "10010001",43059 => "10010010",43060 => "00110100",43061 => "00101110",43062 => "10100110",43063 => "11010100",43064 => "01010011",43065 => "10010111",43066 => "00001110",43067 => "10100111",43068 => "10110111",43069 => "11000011",43070 => "01101101",43071 => "01011010",43072 => "01011010",43073 => "00110101",43074 => "00100000",43075 => "00101110",43076 => "11100011",43077 => "11101101",43078 => "10111010",43079 => "01011100",43080 => "11000100",43081 => "01111001",43082 => "00010000",43083 => "00110001",43084 => "00111111",43085 => "00000111",43086 => "00101100",43087 => "11110001",43088 => "00001101",43089 => "10111011",43090 => "01101000",43091 => "11011101",43092 => "01101100",43093 => "11111010",43094 => "00001110",43095 => "01100010",43096 => "11111001",43097 => "11100111",43098 => "01100010",43099 => "10000011",43100 => "11100000",43101 => "00100101",43102 => "10011011",43103 => "00000000",43104 => "01011111",43105 => "11101001",43106 => "10011100",43107 => "01100110",43108 => "01011100",43109 => "10000110",43110 => "00110111",43111 => "01111101",43112 => "11011001",43113 => "00010100",43114 => "10100111",43115 => "10011010",43116 => "11110101",43117 => "10100111",43118 => "11011110",43119 => "01010101",43120 => "01100011",43121 => "11110110",43122 => "10000000",43123 => "10011000",43124 => "01111101",43125 => "11111010",43126 => "11110000",43127 => "01111001",43128 => "00101001",43129 => "11000100",43130 => "00101100",43131 => "01011011",43132 => "00101000",43133 => "01000101",43134 => "10110011",43135 => "10011100",43136 => "10011101",43137 => "10110010",43138 => "11010010",43139 => "00011101",43140 => "10001001",43141 => "11011111",43142 => "10001100",43143 => "01011110",43144 => "01101011",43145 => "00000001",43146 => "10110010",43147 => "01100101",43148 => "00011100",43149 => "00101100",43150 => "00111110",43151 => "00000001",43152 => "11100111",43153 => "00011110",43154 => "01011011",43155 => "11011011",43156 => "00101100",43157 => "00101010",43158 => "11110101",43159 => "00101000",43160 => "11101000",43161 => "10011001",43162 => "00101010",43163 => "10100010",43164 => "01010001",43165 => "11001010",43166 => "10000101",43167 => "01110010",43168 => "01111100",43169 => "11110010",43170 => "11110111",43171 => "00000111",43172 => "10001000",43173 => "11110110",43174 => "11000011",43175 => "10100101",43176 => "01010100",43177 => "10000011",43178 => "01001100",43179 => "01000011",43180 => "00111011",43181 => "11111000",43182 => "00100110",43183 => "00010101",43184 => "01010110",43185 => "00010001",43186 => "10001101",43187 => "10101001",43188 => "00100111",43189 => "10110001",43190 => "10111010",43191 => "10110011",43192 => "01111101",43193 => "01101100",43194 => "10110100",43195 => "00100011",43196 => "01011110",43197 => "01011001",43198 => "01110110",43199 => "10111110",43200 => "01101101",43201 => "11100110",43202 => "11001101",43203 => "10000010",43204 => "01011101",43205 => "10000101",43206 => "01111110",43207 => "01100011",43208 => "01011100",43209 => "11000100",43210 => "01101111",43211 => "01100110",43212 => "10101010",43213 => "11000101",43214 => "00100110",43215 => "10000101",43216 => "10101111",43217 => "10001101",43218 => "10001001",43219 => "01000110",43220 => "00100010",43221 => "11010110",43222 => "01000100",43223 => "00100111",43224 => "01011000",43225 => "10011111",43226 => "10011010",43227 => "10010011",43228 => "01010000",43229 => "11101100",43230 => "11110001",43231 => "01011101",43232 => "11011010",43233 => "10100111",43234 => "00101010",43235 => "10100110",43236 => "10000010",43237 => "00000101",43238 => "11110100",43239 => "01101101",43240 => "11000000",43241 => "00101001",43242 => "10011111",43243 => "01010110",43244 => "00111111",43245 => "11011011",43246 => "11010001",43247 => "00101101",43248 => "11101111",43249 => "00100101",43250 => "10010010",43251 => "00110000",43252 => "00010100",43253 => "10100110",43254 => "01010001",43255 => "01001001",43256 => "01010110",43257 => "11111000",43258 => "10010000",43259 => "01100100",43260 => "00111010",43261 => "11110110",43262 => "11101010",43263 => "01011101",43264 => "11111011",43265 => "10010000",43266 => "00110000",43267 => "01100110",43268 => "01001010",43269 => "01110110",43270 => "01110011",43271 => "01100110",43272 => "01111011",43273 => "10101001",43274 => "10111110",43275 => "11000011",43276 => "11101101",43277 => "00011101",43278 => "11111010",43279 => "11111001",43280 => "00110010",43281 => "01111000",43282 => "00000000",43283 => "00000000",43284 => "11000101",43285 => "11000000",43286 => "01100001",43287 => "01000110",43288 => "11010101",43289 => "10000001",43290 => "10010010",43291 => "00011000",43292 => "10010111",43293 => "01010100",43294 => "01101001",43295 => "01110010",43296 => "10110010",43297 => "10111000",43298 => "00001111",43299 => "00011000",43300 => "01011111",43301 => "01001011",43302 => "01010001",43303 => "01100111",43304 => "00011110",43305 => "01110010",43306 => "10100101",43307 => "01110010",43308 => "01100011",43309 => "00010101",43310 => "10000010",43311 => "10011100",43312 => "01100100",43313 => "01110100",43314 => "01110100",43315 => "01100000",43316 => "00001000",43317 => "00010000",43318 => "10101011",43319 => "10010010",43320 => "01011001",43321 => "00010100",43322 => "00001100",43323 => "01110100",43324 => "00101011",43325 => "01001011",43326 => "10100111",43327 => "11110011",43328 => "10001011",43329 => "11010110",43330 => "11101010",43331 => "10000100",43332 => "00011010",43333 => "00110101",43334 => "00010101",43335 => "11101110",43336 => "10100100",43337 => "00111010",43338 => "01110010",43339 => "01000110",43340 => "11101011",43341 => "00011001",43342 => "10001110",43343 => "10111011",43344 => "00011000",43345 => "11000100",43346 => "01101111",43347 => "01000010",43348 => "10111011",43349 => "10001111",43350 => "01100000",43351 => "00011100",43352 => "01111000",43353 => "11100001",43354 => "11000000",43355 => "00010110",43356 => "01101001",43357 => "00001100",43358 => "00110111",43359 => "00011001",43360 => "11110001",43361 => "00011110",43362 => "10010110",43363 => "00101101",43364 => "10001010",43365 => "11101111",43366 => "10010010",43367 => "01100011",43368 => "01000111",43369 => "10101000",43370 => "01101111",43371 => "10111101",43372 => "01110001",43373 => "00101000",43374 => "11010000",43375 => "10000011",43376 => "10011110",43377 => "11010010",43378 => "00101101",43379 => "00010100",43380 => "11000111",43381 => "11000101",43382 => "01001000",43383 => "01011000",43384 => "00001111",43385 => "00001010",43386 => "00010010",43387 => "10110010",43388 => "10011001",43389 => "01101010",43390 => "11000000",43391 => "11001011",43392 => "01010000",43393 => "01100100",43394 => "11110011",43395 => "00111011",43396 => "01010001",43397 => "00011101",43398 => "11010110",43399 => "11100010",43400 => "01101111",43401 => "00111110",43402 => "01011011",43403 => "00000011",43404 => "10110011",43405 => "11011101",43406 => "10110010",43407 => "11110111",43408 => "10101100",43409 => "10011010",43410 => "00111000",43411 => "00111101",43412 => "01011111",43413 => "11011000",43414 => "00010001",43415 => "01011111",43416 => "01000111",43417 => "01000011",43418 => "11100000",43419 => "10100001",43420 => "10001010",43421 => "01000100",43422 => "01011000",43423 => "01000000",43424 => "00000011",43425 => "00111001",43426 => "00110111",43427 => "01110111",43428 => "11111101",43429 => "10010010",43430 => "10000001",43431 => "00100001",43432 => "10001001",43433 => "00110001",43434 => "01111111",43435 => "01001010",43436 => "11000011",43437 => "01010110",43438 => "00110101",43439 => "10111100",43440 => "10110001",43441 => "01101011",43442 => "10011001",43443 => "00101001",43444 => "11010001",43445 => "01000001",43446 => "11111000",43447 => "10100010",43448 => "11000000",43449 => "11010010",43450 => "01001000",43451 => "00000001",43452 => "10100010",43453 => "01111110",43454 => "01000111",43455 => "10011110",43456 => "11110111",43457 => "10011111",43458 => "11100101",43459 => "00011011",43460 => "10110110",43461 => "01000101",43462 => "10001010",43463 => "01100001",43464 => "01010000",43465 => "10000111",43466 => "11101001",43467 => "11001110",43468 => "10001111",43469 => "00110101",43470 => "01110111",43471 => "00111001",43472 => "01111010",43473 => "00001111",43474 => "01110011",43475 => "00001101",43476 => "01110010",43477 => "10011001",43478 => "01110010",43479 => "01000010",43480 => "01100001",43481 => "01101001",43482 => "01011111",43483 => "01111000",43484 => "00000011",43485 => "00001010",43486 => "00101011",43487 => "00111100",43488 => "11111000",43489 => "00011111",43490 => "00000001",43491 => "00111010",43492 => "10010011",43493 => "00101011",43494 => "00111001",43495 => "00100100",43496 => "00100001",43497 => "11000111",43498 => "00101001",43499 => "11110101",43500 => "11000010",43501 => "00111011",43502 => "01110011",43503 => "10001001",43504 => "11010100",43505 => "00000101",43506 => "10001010",43507 => "01111101",43508 => "11011110",43509 => "01111010",43510 => "10010001",43511 => "00001111",43512 => "10000000",43513 => "00111010",43514 => "10110010",43515 => "01110110",43516 => "10001001",43517 => "10000101",43518 => "00101101",43519 => "00001101",43520 => "11010011",43521 => "11110000",43522 => "00011101",43523 => "11111110",43524 => "00010011",43525 => "11101101",43526 => "11100010",43527 => "00001100",43528 => "11111000",43529 => "01101110",43530 => "00110001",43531 => "01011110",43532 => "00000101",43533 => "11111001",43534 => "10000011",43535 => "00011011",43536 => "11001011",43537 => "01110111",43538 => "00111101",43539 => "11101011",43540 => "00001010",43541 => "11111101",43542 => "10100111",43543 => "11001010",43544 => "11000011",43545 => "01110110",43546 => "01101010",43547 => "10100101",43548 => "01111010",43549 => "10001011",43550 => "01101101",43551 => "11110111",43552 => "11100101",43553 => "01001000",43554 => "10101100",43555 => "00011100",43556 => "10110001",43557 => "11110010",43558 => "00000110",43559 => "11001110",43560 => "01000111",43561 => "00100011",43562 => "10111100",43563 => "01000011",43564 => "00011010",43565 => "01011100",43566 => "11100100",43567 => "00110010",43568 => "00101110",43569 => "11110110",43570 => "11101010",43571 => "01010010",43572 => "01011111",43573 => "11001011",43574 => "01010111",43575 => "01101010",43576 => "00001010",43577 => "00001100",43578 => "01110111",43579 => "01001111",43580 => "10111110",43581 => "11100100",43582 => "10110000",43583 => "10110100",43584 => "11000110",43585 => "10100011",43586 => "10000011",43587 => "00100101",43588 => "11100100",43589 => "10000001",43590 => "11101100",43591 => "00101111",43592 => "10110010",43593 => "10111100",43594 => "01000111",43595 => "01010111",43596 => "00001001",43597 => "01110111",43598 => "01111001",43599 => "01010001",43600 => "01100000",43601 => "11111100",43602 => "01101101",43603 => "11101011",43604 => "10100000",43605 => "10110111",43606 => "01110111",43607 => "11011111",43608 => "01001000",43609 => "10100000",43610 => "11011100",43611 => "10010011",43612 => "00001101",43613 => "00010101",43614 => "00110010",43615 => "10110110",43616 => "00101000",43617 => "11100100",43618 => "00011100",43619 => "01010110",43620 => "11001111",43621 => "01001100",43622 => "01111001",43623 => "10011001",43624 => "00001110",43625 => "11010011",43626 => "00110011",43627 => "01011101",43628 => "10011111",43629 => "11111000",43630 => "00000101",43631 => "00100111",43632 => "10100011",43633 => "01000001",43634 => "11000011",43635 => "00100011",43636 => "00010100",43637 => "01101011",43638 => "01010101",43639 => "01010000",43640 => "01100011",43641 => "00100110",43642 => "11100011",43643 => "10001111",43644 => "10000100",43645 => "01000111",43646 => "01101111",43647 => "11010110",43648 => "10101110",43649 => "10111010",43650 => "10011011",43651 => "11110100",43652 => "00110000",43653 => "00010100",43654 => "00001001",43655 => "00001001",43656 => "00111000",43657 => "00110011",43658 => "00011001",43659 => "01110001",43660 => "10011110",43661 => "01011010",43662 => "10000010",43663 => "11000001",43664 => "00011001",43665 => "10110111",43666 => "00011010",43667 => "11100001",43668 => "01010001",43669 => "01000001",43670 => "10011100",43671 => "11000110",43672 => "01100000",43673 => "00111011",43674 => "01110101",43675 => "11010100",43676 => "01111001",43677 => "01011111",43678 => "00000001",43679 => "11010111",43680 => "01011010",43681 => "00110110",43682 => "10110111",43683 => "00101110",43684 => "11101111",43685 => "10001001",43686 => "10100000",43687 => "10100011",43688 => "01110010",43689 => "10001010",43690 => "11001010",43691 => "00111101",43692 => "11011101",43693 => "11001010",43694 => "01011100",43695 => "10111011",43696 => "10111010",43697 => "00011111",43698 => "01110100",43699 => "11000011",43700 => "00100010",43701 => "01101101",43702 => "10011000",43703 => "01011000",43704 => "10010101",43705 => "10000000",43706 => "11101110",43707 => "10110011",43708 => "00101001",43709 => "10100001",43710 => "10101101",43711 => "10001110",43712 => "00011000",43713 => "10110101",43714 => "00010001",43715 => "10101011",43716 => "10110110",43717 => "10100001",43718 => "11000100",43719 => "00001010",43720 => "00101101",43721 => "11011110",43722 => "01111001",43723 => "00100011",43724 => "11001101",43725 => "00110010",43726 => "10011010",43727 => "11010100",43728 => "11100001",43729 => "01000100",43730 => "10110110",43731 => "11110110",43732 => "10011111",43733 => "11101111",43734 => "01001110",43735 => "01011110",43736 => "01001101",43737 => "01001001",43738 => "10000011",43739 => "01111001",43740 => "01110011",43741 => "00111100",43742 => "00011110",43743 => "01010101",43744 => "01111011",43745 => "01100100",43746 => "00010110",43747 => "10100110",43748 => "00011100",43749 => "01011010",43750 => "11101010",43751 => "11010001",43752 => "01110111",43753 => "11010100",43754 => "11011010",43755 => "11101001",43756 => "01011010",43757 => "11011001",43758 => "11000110",43759 => "01010111",43760 => "11000101",43761 => "10000001",43762 => "11010101",43763 => "00111001",43764 => "01010100",43765 => "01100011",43766 => "11001100",43767 => "10011101",43768 => "11111111",43769 => "10111010",43770 => "01010111",43771 => "00100101",43772 => "11100101",43773 => "10000001",43774 => "00001110",43775 => "01111010",43776 => "10001011",43777 => "11011000",43778 => "01101110",43779 => "10001111",43780 => "01010101",43781 => "00001101",43782 => "11001001",43783 => "11111110",43784 => "01110111",43785 => "10111001",43786 => "10010010",43787 => "10010011",43788 => "00100100",43789 => "11111011",43790 => "10001110",43791 => "10010101",43792 => "00000111",43793 => "01111110",43794 => "10000100",43795 => "10010111",43796 => "01101001",43797 => "00101110",43798 => "00110001",43799 => "01101000",43800 => "01110110",43801 => "00111101",43802 => "01011001",43803 => "00000110",43804 => "11110001",43805 => "10100010",43806 => "01010000",43807 => "10110011",43808 => "01111000",43809 => "10011001",43810 => "11110000",43811 => "00011100",43812 => "01101000",43813 => "11101010",43814 => "10000011",43815 => "01110001",43816 => "01010001",43817 => "01011111",43818 => "00110000",43819 => "01000011",43820 => "01110100",43821 => "00010110",43822 => "01111001",43823 => "10011111",43824 => "11110100",43825 => "10101100",43826 => "01110000",43827 => "10110010",43828 => "01010101",43829 => "00101101",43830 => "11000001",43831 => "01111001",43832 => "11001111",43833 => "01000101",43834 => "10011010",43835 => "10110010",43836 => "11111111",43837 => "10100000",43838 => "10110100",43839 => "01110000",43840 => "00010001",43841 => "10000111",43842 => "10101100",43843 => "00100000",43844 => "10100001",43845 => "11001100",43846 => "11100100",43847 => "00101010",43848 => "10111101",43849 => "10101101",43850 => "11010101",43851 => "00111001",43852 => "01010110",43853 => "01010000",43854 => "11011000",43855 => "01000000",43856 => "10100110",43857 => "10011111",43858 => "10001011",43859 => "10000100",43860 => "10011101",43861 => "10100110",43862 => "10011110",43863 => "10110000",43864 => "01011001",43865 => "11111011",43866 => "01101010",43867 => "11100111",43868 => "01111111",43869 => "01101100",43870 => "00010011",43871 => "11011111",43872 => "11000000",43873 => "10111111",43874 => "10001100",43875 => "11110000",43876 => "00111100",43877 => "01010100",43878 => "11011101",43879 => "11010001",43880 => "10110100",43881 => "11111100",43882 => "00011000",43883 => "11101010",43884 => "01001101",43885 => "01110110",43886 => "10110001",43887 => "01010010",43888 => "10111100",43889 => "10111100",43890 => "01101111",43891 => "10110011",43892 => "11010100",43893 => "11101011",43894 => "01000111",43895 => "01110111",43896 => "10001110",43897 => "10001011",43898 => "10110100",43899 => "01100001",43900 => "10000000",43901 => "10010101",43902 => "11000001",43903 => "01110111",43904 => "10010001",43905 => "11001001",43906 => "10010110",43907 => "11011101",43908 => "11110000",43909 => "00001011",43910 => "00100100",43911 => "11010101",43912 => "11101110",43913 => "10001010",43914 => "01011100",43915 => "00101001",43916 => "01001111",43917 => "00110000",43918 => "10111001",43919 => "01111101",43920 => "10010110",43921 => "01010011",43922 => "11100010",43923 => "11001011",43924 => "11010101",43925 => "10000111",43926 => "01010011",43927 => "01110101",43928 => "11000110",43929 => "11000110",43930 => "01010011",43931 => "10101110",43932 => "00111011",43933 => "10001001",43934 => "11100011",43935 => "11110111",43936 => "10111110",43937 => "01010011",43938 => "10010010",43939 => "00000110",43940 => "11100010",43941 => "10101000",43942 => "11101010",43943 => "11100110",43944 => "01101011",43945 => "00000000",43946 => "11010001",43947 => "11110001",43948 => "10011010",43949 => "10111010",43950 => "10100000",43951 => "01001110",43952 => "11000101",43953 => "11101100",43954 => "10010101",43955 => "10110101",43956 => "11000100",43957 => "01011101",43958 => "00110001",43959 => "11011010",43960 => "11100001",43961 => "10001000",43962 => "10100110",43963 => "00001110",43964 => "01100111",43965 => "11101110",43966 => "11110000",43967 => "11000111",43968 => "01000111",43969 => "01011010",43970 => "01110110",43971 => "11100101",43972 => "00010100",43973 => "00101111",43974 => "01010110",43975 => "11110111",43976 => "00011110",43977 => "10011000",43978 => "10011001",43979 => "11100000",43980 => "10100010",43981 => "01000010",43982 => "11001101",43983 => "11101111",43984 => "10011100",43985 => "01011111",43986 => "00110111",43987 => "11110010",43988 => "10101011",43989 => "11010111",43990 => "11101000",43991 => "01100010",43992 => "10110001",43993 => "00000000",43994 => "10100111",43995 => "10100010",43996 => "01000111",43997 => "10011011",43998 => "00010101",43999 => "11100010",44000 => "10111101",44001 => "01100000",44002 => "01100000",44003 => "11000100",44004 => "10010110",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "10101011" report "FAIL high bits" severity failure;
assert RAM(0) = "11100100" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
