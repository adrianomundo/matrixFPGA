 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "00110000",3 => "00100011",4 => "01111101",5 => "01000000",6 => "10101110",7 => "01101111",8 => "00101000",9 => "01110000",10 => "10101111",11 => "00010100",12 => "01000110",13 => "01110110",14 => "00101100",15 => "10000111",16 => "10111011",17 => "11101011",18 => "10100011",19 => "01011100",20 => "10001010",21 => "00011010",22 => "10011001",23 => "10000111",24 => "00001101",25 => "00011010",26 => "01001000",27 => "11111011",28 => "00100101",29 => "10111000",30 => "01010110",31 => "11111011",32 => "10000100",33 => "10010110",34 => "10100010",35 => "01000000",36 => "10000111",37 => "01011101",38 => "00110110",39 => "01010110",40 => "10000000",41 => "00001010",42 => "01101110",43 => "00010101",44 => "01011110",45 => "01000001",46 => "00001000",47 => "10111110",48 => "11111111",49 => "00101101",50 => "11100111",51 => "10100000",52 => "01111100",53 => "10010000",54 => "00110011",55 => "10100000",56 => "11000011",57 => "10001110",58 => "01010111",59 => "01011001",60 => "11000101",61 => "00100000",62 => "01110011",63 => "00100011",64 => "01111111",65 => "00110001",66 => "01011110",67 => "01110111",68 => "01110000",69 => "01111111",70 => "01110100",71 => "00001111",72 => "10101011",73 => "00110100",74 => "01101011",75 => "10110001",76 => "00110011",77 => "11110101",78 => "10111111",79 => "00010001",80 => "10010000",81 => "10000111",82 => "10001000",83 => "11101011",84 => "10010010",85 => "00011100",86 => "01101110",87 => "01011011",88 => "00110000",89 => "01111000",90 => "10101011",91 => "10100011",92 => "11000101",93 => "00101100",94 => "11011001",95 => "11100011",96 => "11011000",97 => "00000001",98 => "00000110",99 => "01010001",100 => "11111100",101 => "01010110",102 => "00010100",103 => "10111111",104 => "10011110",105 => "00011001",106 => "11000111",107 => "11010101",108 => "00100000",109 => "11000010",110 => "00001000",111 => "00101110",112 => "01111101",113 => "11110100",114 => "00111010",115 => "11100100",116 => "00101110",117 => "11011010",118 => "11110001",119 => "10110110",120 => "10110000",121 => "10000001",122 => "10101111",123 => "01110101",124 => "10110110",125 => "10011101",126 => "10110100",127 => "10000101",128 => "00110101",129 => "01110100",130 => "01001010",131 => "01100001",132 => "11000111",133 => "01011010",134 => "10011101",135 => "00000101",136 => "01110111",137 => "11000100",138 => "00010000",139 => "01001110",140 => "11010011",141 => "00100001",142 => "10000001",143 => "00111011",144 => "00101110",145 => "11011011",146 => "10101111",147 => "01001010",148 => "01110001",149 => "01001000",150 => "01101100",151 => "10100111",152 => "01010011",153 => "10111001",154 => "01101100",155 => "11011000",156 => "11011001",157 => "10101011",158 => "10101000",159 => "10100010",160 => "11101101",161 => "11000011",162 => "01011111",163 => "10100111",164 => "01110000",165 => "00001100",166 => "01011011",167 => "01011011",168 => "01101110",169 => "00111110",170 => "00110011",171 => "01000000",172 => "00110000",173 => "10011010",174 => "00000010",175 => "01100110",176 => "11110011",177 => "11010010",178 => "01001000",179 => "00011101",180 => "10101010",181 => "01101000",182 => "10101101",183 => "01101101",184 => "10001100",185 => "10111101",186 => "11111101",187 => "10110110",188 => "11101111",189 => "10000011",190 => "01101111",191 => "00011011",192 => "00011110",193 => "10100111",194 => "11110011",195 => "10010101",196 => "00000010",197 => "00100000",198 => "01101111",199 => "10100100",200 => "01010001",201 => "10101100",202 => "01001100",203 => "00010100",204 => "00101010",205 => "10011000",206 => "00000110",207 => "10101001",208 => "10100010",209 => "10110001",210 => "00100110",211 => "11111100",212 => "00000110",213 => "10111110",214 => "10000000",215 => "10101011",216 => "11100101",217 => "11110111",218 => "11011111",219 => "01001111",220 => "00011001",221 => "11100100",222 => "11110011",223 => "10001010",224 => "01111101",225 => "11000110",226 => "11110101",227 => "11111111",228 => "01110110",229 => "01111101",230 => "01011000",231 => "10101011",232 => "01100000",233 => "10111110",234 => "00010000",235 => "01000001",236 => "00010010",237 => "10000011",238 => "11011011",239 => "01001011",240 => "01010001",241 => "01101000",242 => "10011110",243 => "11111011",244 => "00011101",245 => "11110110",246 => "11110010",247 => "11011001",248 => "01101110",249 => "01000110",250 => "01000000",251 => "01110100",252 => "10010010",253 => "01010011",254 => "01111110",255 => "10010110",256 => "10011011",257 => "01000011",258 => "10000011",259 => "01100001",260 => "11101011",261 => "01001000",262 => "01100110",263 => "11010111",264 => "00001000",265 => "10010010",266 => "11111010",267 => "00110100",268 => "11101100",269 => "11101111",270 => "00111011",271 => "00110010",272 => "11001100",273 => "01111010",274 => "00101100",275 => "00101100",276 => "10100000",277 => "01011010",278 => "01101100",279 => "10100100",280 => "01010110",281 => "00101011",282 => "00111110",283 => "00000011",284 => "01101010",285 => "11011101",286 => "11010101",287 => "01001111",288 => "00111011",289 => "01010001",290 => "10111110",291 => "01111011",292 => "01010011",293 => "10101110",294 => "10010110",295 => "11110111",296 => "11000101",297 => "01010001",298 => "01000110",299 => "01010011",300 => "11010010",301 => "10010101",302 => "01100100",303 => "01011110",304 => "10110101",305 => "00000001",306 => "11111111",307 => "10001010",308 => "00010111",309 => "00010011",310 => "11000110",311 => "01111110",312 => "01010101",313 => "01111010",314 => "00110010",315 => "11010101",316 => "11100011",317 => "01111101",318 => "11111000",319 => "00011001",320 => "11001110",321 => "11011010",322 => "10010001",323 => "11010010",324 => "00001000",325 => "11110110",326 => "01111111",327 => "11010111",328 => "10000111",329 => "10111010",330 => "11011011",331 => "00000010",332 => "10010100",333 => "00101101",334 => "00001110",335 => "10000100",336 => "00011100",337 => "10000011",338 => "00111101",339 => "01000111",340 => "11001110",341 => "11101010",342 => "10011110",343 => "11100011",344 => "01100010",345 => "01000010",346 => "01010000",347 => "11110011",348 => "11000000",349 => "10011000",350 => "01001001",351 => "10010010",352 => "01110011",353 => "01110011",354 => "01111010",355 => "01010100",356 => "00001111",357 => "01010111",358 => "11000000",359 => "11100011",360 => "01011101",361 => "00011101",362 => "01110011",363 => "10100110",364 => "10001000",365 => "10110001",366 => "10001111",367 => "01010010",368 => "10010100",369 => "11010001",370 => "00000100",371 => "01000111",372 => "10110001",373 => "11011110",374 => "10101001",375 => "11011001",376 => "00001001",377 => "11110100",378 => "00100110",379 => "11100100",380 => "10111000",381 => "01101000",382 => "10000011",383 => "11011011",384 => "11111110",385 => "00000011",386 => "11011001",387 => "10101010",388 => "10101010",389 => "01010000",390 => "11001010",391 => "11011100",392 => "01010100",393 => "00000011",394 => "00110001",395 => "10001001",396 => "10100000",397 => "11010010",398 => "00010011",399 => "00001111",400 => "10101010",401 => "01000111",402 => "00001010",403 => "00011101",404 => "10001010",405 => "01101111",406 => "11011000",407 => "10001100",408 => "11001110",409 => "10000011",410 => "11010010",411 => "11101110",412 => "01101001",413 => "01000110",414 => "10110100",415 => "11111110",416 => "01011110",417 => "01010000",418 => "01011011",419 => "00101001",420 => "10011111",421 => "00110100",422 => "01101111",423 => "11010111",424 => "10010000",425 => "00111010",426 => "10100010",427 => "11100010",428 => "00101000",429 => "01110000",430 => "01110010",431 => "00100001",432 => "11111100",433 => "01000110",434 => "10100001",435 => "11111010",436 => "01010010",437 => "01010001",438 => "01101000",439 => "10110101",440 => "10010000",441 => "11101110",442 => "10111110",443 => "01000100",444 => "10100011",445 => "11011010",446 => "11011111",447 => "10110010",448 => "10100000",449 => "00101101",450 => "01100011",451 => "00001111",452 => "10010001",453 => "11100100",454 => "01101100",455 => "11101101",456 => "00010111",457 => "10010001",458 => "10101110",459 => "00011100",460 => "10101000",461 => "10000100",462 => "11011011",463 => "10000011",464 => "11001011",465 => "00100110",466 => "01101010",467 => "11000110",468 => "10001101",469 => "00110101",470 => "11011110",471 => "11100101",472 => "11001100",473 => "01101011",474 => "00001001",475 => "01111011",476 => "00111001",477 => "11100010",478 => "01100110",479 => "10100101",480 => "10100010",481 => "01011010",482 => "00100001",483 => "00101001",484 => "10111011",485 => "00111100",486 => "10001111",487 => "10000100",488 => "10001110",489 => "00000000",490 => "11111010",491 => "01100101",492 => "00001010",493 => "10010001",494 => "10010010",495 => "00000101",496 => "10111101",497 => "11111011",498 => "01111010",499 => "00010110",500 => "11100101",501 => "01101000",502 => "11001111",503 => "11001100",504 => "11110010",505 => "01111101",506 => "00001011",507 => "01001110",508 => "01000001",509 => "10000010",510 => "10000111",511 => "10101101",512 => "10001001",513 => "10111101",514 => "11111111",515 => "01111111",516 => "01001100",517 => "11000100",518 => "01010101",519 => "10100100",520 => "11000001",521 => "01110110",522 => "11100111",523 => "11111101",524 => "11010100",525 => "11001111",526 => "00001110",527 => "00010010",528 => "10000001",529 => "10101000",530 => "10011110",531 => "01011110",532 => "00111100",533 => "10100110",534 => "01000111",535 => "01001100",536 => "10001111",537 => "10010010",538 => "10111111",539 => "00111100",540 => "11000001",541 => "00010001",542 => "11000111",543 => "01001010",544 => "10000010",545 => "00011111",546 => "11000101",547 => "10011111",548 => "10001110",549 => "00000000",550 => "11000001",551 => "00111010",552 => "01100001",553 => "11111001",554 => "10011101",555 => "11000000",556 => "10010111",557 => "01001101",558 => "10101010",559 => "11001110",560 => "10001000",561 => "01111100",562 => "11000011",563 => "10100010",564 => "10111010",565 => "01010001",566 => "01000000",567 => "01101110",568 => "01000110",569 => "10100010",570 => "10110010",571 => "10101011",572 => "01110001",573 => "11101111",574 => "00010101",575 => "10110000",576 => "10000000",577 => "01110011",578 => "11110100",579 => "01001000",580 => "10010000",581 => "01001011",582 => "11010010",583 => "11011010",584 => "00101010",585 => "00010110",586 => "10010011",587 => "00011111",588 => "00010111",589 => "11011101",590 => "11010100",591 => "10011000",592 => "00010010",593 => "01011000",594 => "10100000",595 => "11010100",596 => "11100111",597 => "00111011",598 => "10011000",599 => "01100110",600 => "01100010",601 => "01000000",602 => "00011000",603 => "00000101",604 => "11110111",605 => "11111110",606 => "11101001",607 => "00011111",608 => "11100001",609 => "10001001",610 => "01010001",611 => "00001000",612 => "00101001",613 => "11101101",614 => "00000110",615 => "11111000",616 => "00011000",617 => "10100010",618 => "00001100",619 => "01010110",620 => "11010100",621 => "10010011",622 => "00001001",623 => "11011111",624 => "10000100",625 => "11010010",626 => "10000010",627 => "01110111",628 => "10010100",629 => "10001001",630 => "01001010",631 => "10111110",632 => "10100100",633 => "01000000",634 => "01100110",635 => "10110001",636 => "01110001",637 => "01101000",638 => "11000011",639 => "00100011",640 => "01001100",641 => "10100111",642 => "00011111",643 => "01100000",644 => "11100011",645 => "11100111",646 => "10111101",647 => "00101010",648 => "01111111",649 => "10110100",650 => "11100001",651 => "01010101",652 => "11010100",653 => "10000011",654 => "01101111",655 => "11111011",656 => "11101100",657 => "11000011",658 => "01111010",659 => "11101111",660 => "11100110",661 => "01101111",662 => "00001111",663 => "01010100",664 => "10011001",665 => "11010001",666 => "10000011",667 => "00100110",668 => "11001001",669 => "10000011",670 => "01101010",671 => "01001000",672 => "00110010",673 => "10011100",674 => "10000000",675 => "11111011",676 => "01000111",677 => "10100010",678 => "01100101",679 => "00110100",680 => "11001001",681 => "00100110",682 => "10100100",683 => "00001011",684 => "11011010",685 => "10000001",686 => "11100100",687 => "11111011",688 => "10111111",689 => "10000000",690 => "11110010",691 => "01101001",692 => "00001110",693 => "00110100",694 => "11010100",695 => "10001100",696 => "10100101",697 => "01000000",698 => "01101110",699 => "00010000",700 => "11011010",701 => "10001101",702 => "00100011",703 => "11001000",704 => "00000000",705 => "10010011",706 => "00100111",707 => "10111101",708 => "01011001",709 => "00001010",710 => "00101111",711 => "10111101",712 => "01010011",713 => "11111111",714 => "10101001",715 => "01000001",716 => "00011010",717 => "10000111",718 => "00010001",719 => "01101010",720 => "00100110",721 => "11111011",722 => "00101010",723 => "10101100",724 => "10011100",725 => "00110000",726 => "11001000",727 => "00001001",728 => "01001110",729 => "10011110",730 => "10010100",731 => "01110010",732 => "01001001",733 => "00110110",734 => "10010100",735 => "01000001",736 => "00011101",737 => "00101010",738 => "10010001",739 => "11010010",740 => "00101111",741 => "11110001",742 => "00110000",743 => "00011100",744 => "11001100",745 => "00101110",746 => "00101011",747 => "00000111",748 => "11100111",749 => "11010111",750 => "10100100",751 => "11110001",752 => "01010001",753 => "11110101",754 => "11010100",755 => "00010011",756 => "00001010",757 => "11000101",758 => "11000101",759 => "11010000",760 => "00011101",761 => "10101001",762 => "00101001",763 => "11000011",764 => "10010011",765 => "01000001",766 => "00000001",767 => "00011010",768 => "11101011",769 => "00110011",770 => "00000111",771 => "10100011",772 => "11101001",773 => "01111010",774 => "10100100",775 => "00001100",776 => "01100001",777 => "00110111",778 => "00111011",779 => "00100101",780 => "11100111",781 => "11110001",782 => "00110100",783 => "11110111",784 => "10011010",785 => "10101010",786 => "01000110",787 => "11111101",788 => "11101000",789 => "01011110",790 => "10101001",791 => "00101010",792 => "11000101",793 => "00110111",794 => "10010111",795 => "01111011",796 => "11100010",797 => "10100101",798 => "01001001",799 => "00110100",800 => "11000111",801 => "10000011",802 => "10010000",803 => "11001101",804 => "01100101",805 => "00010110",806 => "11001000",807 => "01101111",808 => "00001100",809 => "00111100",810 => "00111101",811 => "01110111",812 => "10011011",813 => "00010000",814 => "10111001",815 => "11110000",816 => "11110011",817 => "10111000",818 => "01001001",819 => "01010101",820 => "11100010",821 => "11001010",822 => "01000100",823 => "01100000",824 => "00001011",825 => "01011000",826 => "00001110",827 => "10101010",828 => "01111010",829 => "00110101",830 => "01001100",831 => "10011101",832 => "00101011",833 => "11100011",834 => "00001110",835 => "11011101",836 => "10010101",837 => "10000100",838 => "10010000",839 => "00111010",840 => "11011100",841 => "00001101",842 => "00111010",843 => "00110011",844 => "01101111",845 => "10000011",846 => "00000001",847 => "11010000",848 => "01011000",849 => "00110111",850 => "01101101",851 => "00000000",852 => "01111011",853 => "10001001",854 => "11111001",855 => "10010101",856 => "11000110",857 => "10111011",858 => "10011000",859 => "11111100",860 => "10100111",861 => "11110100",862 => "10101001",863 => "00100010",864 => "01000010",865 => "01001101",866 => "01000001",867 => "00110110",868 => "11111011",869 => "01100011",870 => "01111110",871 => "10000011",872 => "10101110",873 => "01101100",874 => "01101111",875 => "01110101",876 => "10010100",877 => "00001110",878 => "00110011",879 => "11011110",880 => "10110111",881 => "10101111",882 => "00110000",883 => "10111010",884 => "10010011",885 => "11000010",886 => "00011111",887 => "00000111",888 => "11001001",889 => "10100011",890 => "01000010",891 => "10101100",892 => "10001000",893 => "00000111",894 => "11010110",895 => "10001110",896 => "10100100",897 => "01111111",898 => "00011100",899 => "00101110",900 => "11111101",901 => "01101111",902 => "10001010",903 => "11010001",904 => "11011001",905 => "11010010",906 => "01011110",907 => "01010110",908 => "11110001",909 => "01010001",910 => "11011001",911 => "00110100",912 => "10000100",913 => "10001111",914 => "11010011",915 => "10111100",916 => "00011001",917 => "10010011",918 => "01001111",919 => "01100001",920 => "01000001",921 => "01010100",922 => "01000100",923 => "11010100",924 => "00011111",925 => "11001010",926 => "01001010",927 => "11010011",928 => "10010010",929 => "01010110",930 => "11111101",931 => "00111000",932 => "11001011",933 => "00110110",934 => "10001000",935 => "10110000",936 => "01100100",937 => "10011000",938 => "00110011",939 => "01100011",940 => "11101100",941 => "10000001",942 => "11100110",943 => "10010010",944 => "11010010",945 => "10011011",946 => "10100011",947 => "11010100",948 => "11101001",949 => "00011111",950 => "01101110",951 => "00000011",952 => "11111111",953 => "11100011",954 => "11000010",955 => "01011010",956 => "01110000",957 => "01000111",958 => "11010111",959 => "10110010",960 => "11100100",961 => "00110100",962 => "11010100",963 => "01110111",964 => "00100110",965 => "01000111",966 => "00100111",967 => "01100010",968 => "10011110",969 => "01011100",970 => "01111000",971 => "10101001",972 => "00111101",973 => "10001000",974 => "01011001",975 => "01101100",976 => "00100110",977 => "10101010",978 => "11110000",979 => "00100010",980 => "01000111",981 => "00100101",982 => "01101000",983 => "11010011",984 => "10111000",985 => "01110100",986 => "11101001",987 => "10101001",988 => "10010000",989 => "01100011",990 => "11011001",991 => "01010001",992 => "01100110",993 => "11100010",994 => "01001100",995 => "00110111",996 => "11100111",997 => "00010010",998 => "01110111",999 => "01111111",1000 => "01101000",1001 => "00001101",1002 => "10010100",1003 => "01011000",1004 => "01001110",1005 => "10011110",1006 => "11001000",1007 => "01100001",1008 => "10000110",1009 => "00011001",1010 => "11000100",1011 => "10010101",1012 => "01110000",1013 => "11111100",1014 => "11100011",1015 => "10111011",1016 => "01011111",1017 => "01111001",1018 => "10000101",1019 => "10011110",1020 => "01011110",1021 => "10100000",1022 => "11000100",1023 => "00010001",1024 => "00000010",1025 => "01101110",1026 => "10100000",1027 => "11011110",1028 => "11011000",1029 => "10011100",1030 => "10000011",1031 => "01101000",1032 => "10100110",1033 => "10010111",1034 => "11111000",1035 => "00100001",1036 => "11101110",1037 => "01101001",1038 => "01011110",1039 => "00100110",1040 => "10101111",1041 => "11010100",1042 => "00010110",1043 => "00001010",1044 => "11100010",1045 => "11011100",1046 => "10111000",1047 => "01000111",1048 => "00001000",1049 => "00100110",1050 => "00001010",1051 => "00100010",1052 => "01101100",1053 => "00000000",1054 => "11110011",1055 => "11000000",1056 => "11111111",1057 => "10101100",1058 => "10001000",1059 => "01001101",1060 => "10111001",1061 => "10110111",1062 => "11101100",1063 => "11111101",1064 => "00111111",1065 => "00101100",1066 => "10000110",1067 => "01110100",1068 => "00011000",1069 => "10001111",1070 => "00010111",1071 => "00100011",1072 => "01001100",1073 => "11011011",1074 => "00110101",1075 => "01000100",1076 => "10010101",1077 => "01111000",1078 => "00101011",1079 => "00011111",1080 => "01000011",1081 => "01101000",1082 => "11011000",1083 => "10101100",1084 => "11101101",1085 => "00001110",1086 => "11010011",1087 => "10111101",1088 => "01110010",1089 => "01011110",1090 => "11010100",1091 => "00110100",1092 => "00101110",1093 => "01101011",1094 => "01001101",1095 => "00011000",1096 => "01010011",1097 => "00011111",1098 => "01000000",1099 => "10011111",1100 => "10101101",1101 => "01100010",1102 => "11100111",1103 => "11110110",1104 => "00101101",1105 => "01110111",1106 => "11111110",1107 => "01011100",1108 => "00010001",1109 => "00010010",1110 => "00000110",1111 => "01001001",1112 => "10010110",1113 => "00001100",1114 => "01001101",1115 => "01011101",1116 => "01100000",1117 => "10010010",1118 => "11010111",1119 => "00110100",1120 => "01001011",1121 => "01001100",1122 => "11010110",1123 => "11111001",1124 => "11000011",1125 => "11110001",1126 => "10110111",1127 => "10011011",1128 => "01100110",1129 => "00110010",1130 => "00110100",1131 => "01011000",1132 => "00010100",1133 => "01110101",1134 => "00010100",1135 => "01101111",1136 => "10000100",1137 => "01001001",1138 => "00010101",1139 => "00110000",1140 => "10011100",1141 => "00110010",1142 => "01101010",1143 => "00111110",1144 => "00111100",1145 => "10111001",1146 => "11101111",1147 => "10100000",1148 => "10101111",1149 => "10000100",1150 => "11111110",1151 => "01100011",1152 => "00100001",1153 => "10110001",1154 => "11100100",1155 => "10110110",1156 => "10011100",1157 => "10010111",1158 => "00000110",1159 => "11111111",1160 => "00110001",1161 => "01001010",1162 => "10010101",1163 => "01010100",1164 => "10000001",1165 => "10100111",1166 => "10011101",1167 => "11110101",1168 => "01010001",1169 => "01001000",1170 => "10011101",1171 => "11001100",1172 => "00001100",1173 => "01011000",1174 => "11001010",1175 => "10011001",1176 => "11011111",1177 => "00011001",1178 => "11101010",1179 => "11101101",1180 => "00010001",1181 => "01010110",1182 => "10001000",1183 => "10001011",1184 => "10101101",1185 => "00111111",1186 => "10010100",1187 => "11101110",1188 => "01101101",1189 => "10011101",1190 => "11101111",1191 => "10000000",1192 => "11010001",1193 => "11100110",1194 => "01001011",1195 => "11010000",1196 => "11001010",1197 => "10011111",1198 => "01000011",1199 => "00101100",1200 => "11011101",1201 => "11010100",1202 => "10111000",1203 => "01010100",1204 => "00000011",1205 => "10011011",1206 => "00011110",1207 => "00001100",1208 => "11100010",1209 => "10111111",1210 => "01010001",1211 => "01000111",1212 => "11111001",1213 => "00011000",1214 => "01010010",1215 => "10110011",1216 => "00101000",1217 => "01110110",1218 => "01110111",1219 => "10110101",1220 => "10000000",1221 => "11000000",1222 => "01101000",1223 => "10001001",1224 => "11101100",1225 => "11010000",1226 => "01110101",1227 => "01000101",1228 => "01101010",1229 => "00101100",1230 => "01010111",1231 => "11111000",1232 => "00001101",1233 => "00000001",1234 => "10100110",1235 => "01110011",1236 => "11011000",1237 => "01110011",1238 => "01101110",1239 => "01000110",1240 => "10000100",1241 => "11001110",1242 => "11110100",1243 => "11111001",1244 => "11101111",1245 => "10111000",1246 => "01000000",1247 => "01000010",1248 => "11001100",1249 => "11110111",1250 => "11110111",1251 => "00110011",1252 => "00110001",1253 => "01011100",1254 => "11010100",1255 => "10110111",1256 => "11001011",1257 => "11111010",1258 => "10110000",1259 => "11110001",1260 => "01011001",1261 => "10101100",1262 => "01101111",1263 => "01100111",1264 => "11110001",1265 => "11001011",1266 => "10001111",1267 => "00000011",1268 => "11100100",1269 => "01110100",1270 => "10000110",1271 => "10010010",1272 => "11001110",1273 => "11101010",1274 => "10011100",1275 => "11100001",1276 => "01011001",1277 => "11010000",1278 => "01010010",1279 => "10100001",1280 => "01110001",1281 => "01110000",1282 => "00010100",1283 => "01111110",1284 => "01110101",1285 => "11100010",1286 => "10101101",1287 => "10101010",1288 => "11101001",1289 => "11011001",1290 => "11111010",1291 => "00111100",1292 => "01010101",1293 => "00111101",1294 => "00000110",1295 => "00110110",1296 => "10011000",1297 => "11100110",1298 => "00010011",1299 => "00001100",1300 => "01111001",1301 => "11001010",1302 => "11100010",1303 => "01001111",1304 => "11000111",1305 => "10110010",1306 => "10011000",1307 => "11111101",1308 => "11110110",1309 => "11101110",1310 => "01110111",1311 => "00110110",1312 => "00110011",1313 => "00011011",1314 => "00000111",1315 => "00000110",1316 => "10100110",1317 => "01000110",1318 => "11010111",1319 => "11100110",1320 => "10001001",1321 => "01100101",1322 => "10111010",1323 => "10110000",1324 => "11101110",1325 => "10111000",1326 => "00110011",1327 => "10101010",1328 => "01000010",1329 => "11000111",1330 => "11101110",1331 => "01010000",1332 => "10011001",1333 => "00011100",1334 => "01110101",1335 => "00111100",1336 => "01101111",1337 => "11110110",1338 => "01000011",1339 => "10011110",1340 => "10100011",1341 => "10110001",1342 => "10111110",1343 => "01101011",1344 => "11000100",1345 => "10000100",1346 => "11110000",1347 => "01111101",1348 => "01101010",1349 => "00100010",1350 => "00110000",1351 => "01000010",1352 => "11001011",1353 => "10001110",1354 => "11001001",1355 => "00110001",1356 => "11110010",1357 => "11111010",1358 => "11000010",1359 => "11100101",1360 => "11001001",1361 => "10101101",1362 => "10111100",1363 => "00001000",1364 => "01010001",1365 => "10000101",1366 => "00010000",1367 => "01011101",1368 => "00101000",1369 => "11000110",1370 => "00110101",1371 => "10100111",1372 => "01111001",1373 => "10001011",1374 => "10011010",1375 => "10000111",1376 => "01010011",1377 => "01011100",1378 => "10100111",1379 => "10100000",1380 => "00110110",1381 => "01000000",1382 => "01011101",1383 => "10100010",1384 => "00101110",1385 => "10010011",1386 => "01111001",1387 => "01010001",1388 => "01011101",1389 => "10100001",1390 => "10110000",1391 => "01101100",1392 => "00110101",1393 => "01100011",1394 => "10101100",1395 => "00101111",1396 => "00000011",1397 => "11001111",1398 => "01111100",1399 => "10101010",1400 => "11001100",1401 => "11111100",1402 => "11101110",1403 => "11000111",1404 => "01010100",1405 => "10111011",1406 => "11111110",1407 => "00111101",1408 => "01000100",1409 => "11100010",1410 => "10011010",1411 => "00101001",1412 => "01011010",1413 => "01101100",1414 => "11010110",1415 => "11011000",1416 => "11000101",1417 => "01110100",1418 => "10011100",1419 => "01101100",1420 => "01110010",1421 => "01010010",1422 => "01010011",1423 => "00111111",1424 => "01010101",1425 => "11011011",1426 => "01111110",1427 => "10111011",1428 => "11101100",1429 => "00110100",1430 => "10001101",1431 => "10001000",1432 => "10101000",1433 => "00110101",1434 => "11111101",1435 => "00010001",1436 => "10101011",1437 => "01101000",1438 => "11001111",1439 => "11111001",1440 => "01001100",1441 => "11000111",1442 => "00001101",1443 => "11000111",1444 => "10000111",1445 => "10111010",1446 => "01011111",1447 => "00101110",1448 => "00010001",1449 => "11001001",1450 => "10001111",1451 => "00111100",1452 => "00101100",1453 => "11101101",1454 => "00011101",1455 => "00100010",1456 => "01110111",1457 => "10000110",1458 => "10101101",1459 => "10110100",1460 => "00001010",1461 => "01101011",1462 => "10101110",1463 => "01011000",1464 => "01110001",1465 => "00100110",1466 => "10101011",1467 => "10011001",1468 => "00011111",1469 => "10111010",1470 => "00100001",1471 => "00010101",1472 => "01000110",1473 => "01011000",1474 => "11000111",1475 => "00110101",1476 => "10000110",1477 => "01000111",1478 => "01001100",1479 => "01100100",1480 => "11010100",1481 => "10011110",1482 => "11110000",1483 => "01011111",1484 => "01000001",1485 => "10010110",1486 => "00100100",1487 => "11010101",1488 => "01111010",1489 => "00111110",1490 => "11001000",1491 => "00101100",1492 => "01110101",1493 => "01001001",1494 => "11010111",1495 => "11101111",1496 => "00011010",1497 => "00000110",1498 => "00001101",1499 => "01100001",1500 => "10011110",1501 => "10011111",1502 => "11101110",1503 => "11011100",1504 => "11101011",1505 => "11101111",1506 => "10010011",1507 => "11111001",1508 => "01101001",1509 => "01101011",1510 => "00010001",1511 => "10011011",1512 => "10011000",1513 => "10101010",1514 => "11110000",1515 => "00010101",1516 => "00000101",1517 => "00100101",1518 => "00101001",1519 => "11001010",1520 => "10100011",1521 => "00010010",1522 => "10100100",1523 => "01100111",1524 => "10100000",1525 => "10010100",1526 => "11001010",1527 => "01101111",1528 => "11111111",1529 => "00100011",1530 => "00001011",1531 => "10000110",1532 => "00110000",1533 => "01110100",1534 => "11100101",1535 => "10000011",1536 => "11001011",1537 => "10100101",1538 => "00101011",1539 => "10011001",1540 => "01000111",1541 => "01011010",1542 => "00011101",1543 => "01011001",1544 => "00100100",1545 => "00111100",1546 => "10000101",1547 => "01101011",1548 => "00101001",1549 => "11100100",1550 => "00011010",1551 => "11001100",1552 => "11010010",1553 => "01101000",1554 => "10010010",1555 => "00101101",1556 => "00100101",1557 => "10001010",1558 => "01001011",1559 => "10011010",1560 => "10111110",1561 => "00010110",1562 => "10111110",1563 => "01101101",1564 => "11001110",1565 => "01110100",1566 => "01110010",1567 => "11100111",1568 => "10111100",1569 => "01011100",1570 => "11101111",1571 => "10000010",1572 => "11100110",1573 => "11011011",1574 => "11110011",1575 => "01100110",1576 => "00111011",1577 => "01101110",1578 => "01100101",1579 => "11010100",1580 => "11010111",1581 => "01100001",1582 => "01101011",1583 => "01000110",1584 => "10011100",1585 => "10010010",1586 => "01000100",1587 => "00100011",1588 => "11000110",1589 => "11000000",1590 => "10001000",1591 => "11101010",1592 => "01001100",1593 => "01101001",1594 => "01001101",1595 => "00111001",1596 => "00000111",1597 => "11001010",1598 => "00000011",1599 => "10010100",1600 => "00000011",1601 => "10000111",1602 => "11000111",1603 => "11001101",1604 => "10010000",1605 => "11011100",1606 => "01100101",1607 => "10011100",1608 => "01101110",1609 => "11101111",1610 => "11111011",1611 => "10100010",1612 => "11111101",1613 => "10100011",1614 => "10011011",1615 => "00010000",1616 => "10101001",1617 => "10111000",1618 => "01010010",1619 => "11000101",1620 => "00111001",1621 => "11101010",1622 => "00010000",1623 => "01001000",1624 => "11100110",1625 => "01011100",1626 => "01100000",1627 => "00100100",1628 => "01100000",1629 => "01001101",1630 => "11000101",1631 => "10001110",1632 => "11000000",1633 => "00010001",1634 => "01101001",1635 => "10000011",1636 => "11010101",1637 => "11100010",1638 => "11001111",1639 => "10110011",1640 => "10010100",1641 => "11011001",1642 => "00100010",1643 => "10011011",1644 => "10001111",1645 => "01100000",1646 => "10001111",1647 => "01110110",1648 => "11110010",1649 => "01000100",1650 => "00110110",1651 => "01001010",1652 => "10010100",1653 => "01011000",1654 => "11010010",1655 => "01110001",1656 => "00111000",1657 => "11100110",1658 => "00001000",1659 => "00001000",1660 => "01110101",1661 => "10110011",1662 => "00011011",1663 => "11100110",1664 => "01011010",1665 => "10111101",1666 => "10000011",1667 => "00010111",1668 => "00101000",1669 => "10011111",1670 => "10111111",1671 => "11001101",1672 => "10110110",1673 => "01000000",1674 => "11000010",1675 => "10011011",1676 => "01111010",1677 => "11111111",1678 => "10000000",1679 => "11001101",1680 => "01011100",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00000110" report "FAIL high bits" severity failure;
assert RAM(0) = "10010000" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
