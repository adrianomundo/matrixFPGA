 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01010011",3 => "10110100",4 => "10000100",5 => "10011110",6 => "00000001",7 => "10010111",8 => "11110010",9 => "01100101",10 => "10011000",11 => "01100111",12 => "01001100",13 => "10100011",14 => "10010100",15 => "11011101",16 => "10101011",17 => "01000110",18 => "11001001",19 => "01101111",20 => "10100011",21 => "00011110",22 => "00001100",23 => "00010011",24 => "01010110",25 => "00010110",26 => "10111101",27 => "01011111",28 => "00011001",29 => "00100010",30 => "11110111",31 => "10100100",32 => "00110100",33 => "00110111",34 => "01000101",35 => "01101001",36 => "10100111",37 => "10001101",38 => "01110111",39 => "10111011",40 => "11100111",41 => "00100000",42 => "10111100",43 => "10111100",44 => "00110111",45 => "11001101",46 => "11000001",47 => "01011111",48 => "11000000",49 => "00011010",50 => "11011100",51 => "01100011",52 => "11010101",53 => "00100011",54 => "10110001",55 => "00100110",56 => "10011000",57 => "10111110",58 => "00011000",59 => "10000111",60 => "01110100",61 => "00011010",62 => "00101001",63 => "10011100",64 => "00010010",65 => "01110010",66 => "11001011",67 => "10001001",68 => "01100101",69 => "10100011",70 => "00101100",71 => "10100000",72 => "11101000",73 => "11101100",74 => "00001001",75 => "10001010",76 => "01110000",77 => "10011101",78 => "01100110",79 => "00001110",80 => "01001011",81 => "01011101",82 => "10010001",83 => "10110110",84 => "10000101",85 => "01110000",86 => "00110000",87 => "01111001",88 => "10001111",89 => "00000010",90 => "10001100",91 => "00010101",92 => "11100100",93 => "00010010",94 => "11111011",95 => "01110101",96 => "00110011",97 => "01100011",98 => "00011111",99 => "10011011",100 => "01101101",101 => "01010010",102 => "11100001",103 => "10111000",104 => "00101010",105 => "10000001",106 => "01110100",107 => "00101101",108 => "11110111",109 => "10010010",110 => "01101101",111 => "00011011",112 => "11000011",113 => "01001101",114 => "11111110",115 => "11010010",116 => "11110010",117 => "01010001",118 => "00110000",119 => "00000000",120 => "10001011",121 => "10101000",122 => "11100010",123 => "01100101",124 => "11110111",125 => "01010001",126 => "10110110",127 => "10100001",128 => "00111010",129 => "10110100",130 => "10010110",131 => "10001110",132 => "10101000",133 => "00000010",134 => "10111010",135 => "10001011",136 => "11101111",137 => "10000010",138 => "10100000",139 => "01101011",140 => "10111011",141 => "10010000",142 => "01100111",143 => "10000110",144 => "00100011",145 => "00001010",146 => "11100100",147 => "10101100",148 => "01011111",149 => "11001101",150 => "10000100",151 => "11100111",152 => "01101101",153 => "10011110",154 => "11001000",155 => "00011111",156 => "00101000",157 => "11111000",158 => "01110101",159 => "11110010",160 => "11111011",161 => "10010001",162 => "11001000",163 => "10001110",164 => "00101000",165 => "10011111",166 => "01101001",167 => "11001111",168 => "11011100",169 => "01100111",170 => "10111110",171 => "10010001",172 => "00011000",173 => "00100111",174 => "11001011",175 => "10001001",176 => "10001110",177 => "00101011",178 => "11001101",179 => "00011010",180 => "01100001",181 => "11101011",182 => "00011101",183 => "10100010",184 => "11100011",185 => "01100111",186 => "00001101",187 => "00001101",188 => "01000101",189 => "01111111",190 => "11100101",191 => "01000001",192 => "10100110",193 => "00010100",194 => "00011011",195 => "10010111",196 => "01010011",197 => "11000001",198 => "11110001",199 => "01111011",200 => "01111000",201 => "10101110",202 => "11111110",203 => "10001001",204 => "10100110",205 => "01100111",206 => "00000100",207 => "00111101",208 => "10001110",209 => "10100000",210 => "00110110",211 => "00111010",212 => "10001000",213 => "11010101",214 => "11010000",215 => "00100011",216 => "10011111",217 => "11011000",218 => "01100001",219 => "10000111",220 => "00000110",221 => "10010101",222 => "11000110",223 => "11111101",224 => "10001111",225 => "00100100",226 => "01001110",227 => "10101010",228 => "01000100",229 => "11100011",230 => "01111010",231 => "01100111",232 => "01001001",233 => "00101011",234 => "11001110",235 => "01111110",236 => "00101111",237 => "01100001",238 => "01100100",239 => "01101111",240 => "11011011",241 => "10100101",242 => "11111001",243 => "00001000",244 => "10111010",245 => "00101101",246 => "00010100",247 => "11100111",248 => "11110111",249 => "11110010",250 => "01101001",251 => "10001011",252 => "10101011",253 => "00110000",254 => "00011001",255 => "01001100",256 => "11111011",257 => "10000110",258 => "00100110",259 => "00011001",260 => "10010011",261 => "01111011",262 => "01011011",263 => "00100110",264 => "11001110",265 => "01101010",266 => "11011010",267 => "11100010",268 => "01000110",269 => "11001110",270 => "11000000",271 => "10010110",272 => "00110100",273 => "11001100",274 => "10010111",275 => "00111000",276 => "00100000",277 => "11110101",278 => "11000101",279 => "00100011",280 => "00010101",281 => "01110110",282 => "11011000",283 => "00100110",284 => "11001000",285 => "11000101",286 => "11100100",287 => "11101111",288 => "00110001",289 => "11101000",290 => "10000010",291 => "10101001",292 => "00011000",293 => "01111101",294 => "00000000",295 => "00011111",296 => "00001100",297 => "01000110",298 => "10110101",299 => "11100110",300 => "11111100",301 => "01110100",302 => "11011011",303 => "01100100",304 => "10010000",305 => "11010000",306 => "10010110",307 => "10001101",308 => "00011111",309 => "10100100",310 => "10110100",311 => "01000011",312 => "11000000",313 => "11000010",314 => "11100011",315 => "00111011",316 => "00010000",317 => "10100110",318 => "00110100",319 => "00110111",320 => "01100000",321 => "01001100",322 => "00111010",323 => "11011101",324 => "00010010",325 => "01111010",326 => "11110111",327 => "01001011",328 => "00101010",329 => "00010010",330 => "01101111",331 => "11010001",332 => "10011100",333 => "00101000",334 => "10110001",335 => "11110010",336 => "01011001",337 => "11010010",338 => "00101001",339 => "01111000",340 => "10011010",341 => "11100000",342 => "11000101",343 => "00000000",344 => "11110011",345 => "11000100",346 => "01010001",347 => "01100000",348 => "11000011",349 => "01101101",350 => "00010001",351 => "10111011",352 => "11111010",353 => "01000101",354 => "10001110",355 => "10011001",356 => "01000000",357 => "10101000",358 => "01000010",359 => "11000000",360 => "10001001",361 => "11000000",362 => "01000111",363 => "00001001",364 => "00101000",365 => "01101101",366 => "01010100",367 => "00111010",368 => "00110111",369 => "11100100",370 => "00101011",371 => "01110010",372 => "10010010",373 => "00101010",374 => "01101000",375 => "00000111",376 => "11111111",377 => "01011011",378 => "01110001",379 => "00111100",380 => "00110110",381 => "00010001",382 => "10111101",383 => "11111011",384 => "10110111",385 => "01000100",386 => "10101001",387 => "11100000",388 => "00001000",389 => "11111110",390 => "11100110",391 => "00110010",392 => "00000110",393 => "11000100",394 => "01011011",395 => "11000101",396 => "11101010",397 => "00010001",398 => "11101100",399 => "10100110",400 => "10111111",401 => "00111101",402 => "10111011",403 => "00111110",404 => "11000000",405 => "00010110",406 => "11101100",407 => "00101111",408 => "01011011",409 => "01000011",410 => "00100010",411 => "11000110",412 => "10110100",413 => "10010000",414 => "11100100",415 => "11110100",416 => "10101111",417 => "11001000",418 => "11001110",419 => "11111100",420 => "01010011",421 => "10000101",422 => "00001000",423 => "10100111",424 => "00111000",425 => "10110111",426 => "00000101",427 => "11100010",428 => "00010010",429 => "10100010",430 => "00010100",431 => "01001011",432 => "00011101",433 => "00101011",434 => "00011101",435 => "00111100",436 => "11101010",437 => "00001010",438 => "10101100",439 => "01110101",440 => "00010100",441 => "10010111",442 => "11101111",443 => "11101010",444 => "10000011",445 => "11100101",446 => "00010100",447 => "00101011",448 => "10011110",449 => "10101110",450 => "11010110",451 => "01001110",452 => "10011111",453 => "00100001",454 => "11001000",455 => "10000011",456 => "10110010",457 => "11001010",458 => "11001110",459 => "11000011",460 => "00111000",461 => "11111000",462 => "10000011",463 => "01011001",464 => "11101101",465 => "11100110",466 => "10100111",467 => "01100111",468 => "11001000",469 => "11110010",470 => "00110100",471 => "00110101",472 => "00011010",473 => "00100000",474 => "01000010",475 => "00111111",476 => "00010101",477 => "00110111",478 => "00111100",479 => "11101111",480 => "11011111",481 => "11010101",482 => "11010000",483 => "10010101",484 => "01100101",485 => "00100000",486 => "00001000",487 => "10001000",488 => "00011110",489 => "10001010",490 => "11111100",491 => "11011110",492 => "01101010",493 => "00110111",494 => "10110011",495 => "01001101",496 => "00110111",497 => "00001011",498 => "10110111",499 => "01111011",500 => "10010010",501 => "11100100",502 => "01011000",503 => "11001111",504 => "10111011",505 => "10011011",506 => "01101000",507 => "11110011",508 => "00011001",509 => "01000110",510 => "11111001",511 => "00010111",512 => "10000001",513 => "01110101",514 => "01010011",515 => "10110100",516 => "01111001",517 => "10111110",518 => "00000100",519 => "00001100",520 => "11010001",521 => "00001110",522 => "11110011",523 => "11110011",524 => "10000001",525 => "10110101",526 => "11100101",527 => "10110000",528 => "10110011",529 => "00100110",530 => "01001101",531 => "01001000",532 => "01010001",533 => "00010011",534 => "01110011",535 => "11101111",536 => "10100111",537 => "01110110",538 => "10011010",539 => "11100100",540 => "00010010",541 => "11111100",542 => "00111000",543 => "00100100",544 => "10001000",545 => "10100101",546 => "01001001",547 => "11101111",548 => "11010010",549 => "01111010",550 => "11110000",551 => "11000101",552 => "01010111",553 => "01111001",554 => "01011010",555 => "00011100",556 => "00101001",557 => "00101011",558 => "00010110",559 => "00000110",560 => "01111011",561 => "11110111",562 => "10011100",563 => "11010000",564 => "01001000",565 => "00110001",566 => "01000001",567 => "10100101",568 => "11010101",569 => "10000101",570 => "00110111",571 => "10100101",572 => "11001011",573 => "10010000",574 => "10010101",575 => "11100111",576 => "10010101",577 => "01011001",578 => "00111101",579 => "11111101",580 => "11100111",581 => "01100110",582 => "00110101",583 => "00101101",584 => "11110101",585 => "11111100",586 => "01011011",587 => "10010010",588 => "00110110",589 => "11110100",590 => "10011111",591 => "00101011",592 => "10000110",593 => "01001001",594 => "00101010",595 => "11101001",596 => "01001111",597 => "11001011",598 => "01111100",599 => "01101011",600 => "11100100",601 => "01101110",602 => "10110100",603 => "01000000",604 => "00010101",605 => "00110100",606 => "01110000",607 => "00100111",608 => "11000011",609 => "11111101",610 => "11011101",611 => "00010101",612 => "11100000",613 => "11100110",614 => "10101110",615 => "01100111",616 => "01100010",617 => "01100110",618 => "01001010",619 => "01110001",620 => "11100000",621 => "00100001",622 => "00101100",623 => "10000010",624 => "01100110",625 => "00000110",626 => "00110111",627 => "11110101",628 => "10111001",629 => "11010101",630 => "00110010",631 => "00110010",632 => "11110100",633 => "11100000",634 => "11111100",635 => "01010111",636 => "00111101",637 => "10101010",638 => "10100011",639 => "11100110",640 => "01100011",641 => "10010010",642 => "10010000",643 => "01001111",644 => "11101101",645 => "11000100",646 => "01111000",647 => "00101010",648 => "00011110",649 => "00011100",650 => "10110011",651 => "00110101",652 => "11110000",653 => "11000000",654 => "00010010",655 => "11001111",656 => "01111101",657 => "11011000",658 => "10010101",659 => "11100100",660 => "00110101",661 => "10011111",662 => "00111011",663 => "01101001",664 => "11010101",665 => "10000011",666 => "11000001",667 => "11110010",668 => "01101111",669 => "01101011",670 => "00000101",671 => "10010110",672 => "00111101",673 => "10010001",674 => "01000101",675 => "10000110",676 => "11110000",677 => "01101000",678 => "00001110",679 => "11000100",680 => "10100101",681 => "01100100",682 => "01010110",683 => "00010000",684 => "10010001",685 => "00001101",686 => "10100011",687 => "00011101",688 => "01001111",689 => "11000100",690 => "00010100",691 => "10001011",692 => "10010010",693 => "00011101",694 => "01101111",695 => "10001011",696 => "10001000",697 => "11110001",698 => "10111111",699 => "11000001",700 => "10101101",701 => "00000000",702 => "11100101",703 => "10101010",704 => "11011100",705 => "01001010",706 => "10010110",707 => "10011010",708 => "11101111",709 => "00111001",710 => "11100110",711 => "00110100",712 => "00000110",713 => "00001111",714 => "01111101",715 => "11011110",716 => "01110110",717 => "10111011",718 => "00010110",719 => "01101011",720 => "10010000",721 => "00001110",722 => "11100100",723 => "11110110",724 => "00100000",725 => "11000010",726 => "01110010",727 => "11100110",728 => "00000001",729 => "11100011",730 => "00000000",731 => "10111011",732 => "11010110",733 => "10100000",734 => "01111000",735 => "10010011",736 => "11101001",737 => "10000010",738 => "11111111",739 => "11100011",740 => "11001011",741 => "01101010",742 => "00111101",743 => "00101110",744 => "11110000",745 => "01100101",746 => "01100011",747 => "10100111",748 => "01000111",749 => "10101000",750 => "01000110",751 => "11110101",752 => "11111001",753 => "11111000",754 => "10010011",755 => "00000010",756 => "00001011",757 => "10011011",758 => "10010011",759 => "00111000",760 => "01110100",761 => "10111011",762 => "10110001",763 => "01011010",764 => "10110100",765 => "00000101",766 => "01111011",767 => "10110111",768 => "00001000",769 => "01001011",770 => "00100010",771 => "00101100",772 => "00101010",773 => "01011010",774 => "01000111",775 => "11000101",776 => "10000001",777 => "10100010",778 => "11000000",779 => "00100000",780 => "11001101",781 => "00011110",782 => "00000101",783 => "01011001",784 => "00001111",785 => "11010000",786 => "01101100",787 => "01001000",788 => "01001010",789 => "00011100",790 => "01000110",791 => "00011001",792 => "00001001",793 => "00010001",794 => "00000011",795 => "01111001",796 => "10001100",797 => "10110111",798 => "01000100",799 => "10101110",800 => "10001001",801 => "10110011",802 => "11010111",803 => "00111100",804 => "01010011",805 => "10111011",806 => "01110101",807 => "10010110",808 => "11000000",809 => "11010000",810 => "10011001",811 => "11100010",812 => "11110000",813 => "00010010",814 => "11100000",815 => "00100101",816 => "11010100",817 => "10101100",818 => "10100000",819 => "00010011",820 => "00110101",821 => "11101001",822 => "10100000",823 => "10000101",824 => "11111100",825 => "00111010",826 => "00111110",827 => "10000001",828 => "10111110",829 => "01111110",830 => "11101001",831 => "01111000",832 => "10011001",833 => "11000111",834 => "01000101",835 => "10101001",836 => "11110111",837 => "01101100",838 => "10110011",839 => "11011001",840 => "11000111",841 => "10110000",842 => "11010000",843 => "00110110",844 => "00010010",845 => "00101111",846 => "11111001",847 => "00000111",848 => "01000110",849 => "01111110",850 => "10110101",851 => "11000011",852 => "11000111",853 => "11111101",854 => "11000000",855 => "10010001",856 => "01001111",857 => "10011000",858 => "00010011",859 => "11011111",860 => "01110100",861 => "11001000",862 => "10001111",863 => "11011110",864 => "00001000",865 => "11110010",866 => "10100111",867 => "01101110",868 => "00000111",869 => "11100011",870 => "00011011",871 => "01001001",872 => "11100111",873 => "10000100",874 => "11101100",875 => "11101111",876 => "11100110",877 => "11011101",878 => "01110011",879 => "10011100",880 => "11011111",881 => "11001001",882 => "00010001",883 => "10011001",884 => "10101100",885 => "10110111",886 => "00010101",887 => "01010010",888 => "00110001",889 => "10000011",890 => "01001110",891 => "10000011",892 => "01011100",893 => "01011001",894 => "01101010",895 => "10001111",896 => "11000011",897 => "01111000",898 => "01101011",899 => "00110010",900 => "00100001",901 => "10010011",902 => "01111111",903 => "10100011",904 => "10011011",905 => "00100010",906 => "11110101",907 => "01001011",908 => "01000001",909 => "11100011",910 => "11011100",911 => "11011110",912 => "10010101",913 => "01000000",914 => "01011001",915 => "10101111",916 => "11011000",917 => "00101110",918 => "00010000",919 => "11011110",920 => "11000000",921 => "10010111",922 => "01010001",923 => "10100100",924 => "10011000",925 => "11010110",926 => "11100110",927 => "01101011",928 => "11100110",929 => "01110101",930 => "10101010",931 => "11100101",932 => "00000010",933 => "11111010",934 => "11100100",935 => "11000110",936 => "10011101",937 => "10100101",938 => "01110000",939 => "10100100",940 => "10111101",941 => "11011011",942 => "10111000",943 => "11000000",944 => "10011111",945 => "10001110",946 => "01001001",947 => "11001100",948 => "10000100",949 => "11001001",950 => "11011000",951 => "10101101",952 => "00011101",953 => "00011111",954 => "11100101",955 => "10000111",956 => "10110010",957 => "11001111",958 => "01110010",959 => "01001101",960 => "11110100",961 => "10011010",962 => "10100000",963 => "10100110",964 => "10110110",965 => "11010110",966 => "01011000",967 => "11111010",968 => "01111100",969 => "10110010",970 => "10011111",971 => "11011001",972 => "10001000",973 => "11110001",974 => "00011100",975 => "11110110",976 => "11101111",977 => "11100101",978 => "01100101",979 => "01110100",980 => "11100101",981 => "10100001",982 => "01001010",983 => "11111000",984 => "10010101",985 => "01000001",986 => "11111000",987 => "10100001",988 => "11101110",989 => "00010011",990 => "10000000",991 => "00111100",992 => "01100110",993 => "10010001",994 => "11110111",995 => "10101001",996 => "11001010",997 => "00000011",998 => "00101011",999 => "10000011",1000 => "10000010",1001 => "11011000",1002 => "10001000",1003 => "11111110",1004 => "00100000",1005 => "10001001",1006 => "00000110",1007 => "10000000",1008 => "10011111",1009 => "00011000",1010 => "10010011",1011 => "10011100",1012 => "01101110",1013 => "00000000",1014 => "11101011",1015 => "10001101",1016 => "10101110",1017 => "01010111",1018 => "00110011",1019 => "00101001",1020 => "01010101",1021 => "10011001",1022 => "00100000",1023 => "00110011",1024 => "10101011",1025 => "00010001",1026 => "10011000",1027 => "01011110",1028 => "11101001",1029 => "11001000",1030 => "01001100",1031 => "10000100",1032 => "10111010",1033 => "11111011",1034 => "01111010",1035 => "11001111",1036 => "11101110",1037 => "10101011",1038 => "00010111",1039 => "10101010",1040 => "11010001",1041 => "00010100",1042 => "00001000",1043 => "01001110",1044 => "10011111",1045 => "00110100",1046 => "11011010",1047 => "01000001",1048 => "00001000",1049 => "11010010",1050 => "00100110",1051 => "10100101",1052 => "01011001",1053 => "10100101",1054 => "11001111",1055 => "11101110",1056 => "00110000",1057 => "00100000",1058 => "00011001",1059 => "10111111",1060 => "10011010",1061 => "10100001",1062 => "01101010",1063 => "11111100",1064 => "11001101",1065 => "11110011",1066 => "11011001",1067 => "11101100",1068 => "10101110",1069 => "01011011",1070 => "10111011",1071 => "11011010",1072 => "10010110",1073 => "01011100",1074 => "01000101",1075 => "01011011",1076 => "00001110",1077 => "11101010",1078 => "00100111",1079 => "01011110",1080 => "00010010",1081 => "01010010",1082 => "11011001",1083 => "00101111",1084 => "11101101",1085 => "10101011",1086 => "00101111",1087 => "00111001",1088 => "11111100",1089 => "00001101",1090 => "10011001",1091 => "10001000",1092 => "00110101",1093 => "10110000",1094 => "00000111",1095 => "01101111",1096 => "10001111",1097 => "00010100",1098 => "11001001",1099 => "01111000",1100 => "01110110",1101 => "00010000",1102 => "11011110",1103 => "01100000",1104 => "01011001",1105 => "01010010",1106 => "11111000",1107 => "01001000",1108 => "11101100",1109 => "10010011",1110 => "10011100",1111 => "00000001",1112 => "11011000",1113 => "00110100",1114 => "11110100",1115 => "00110101",1116 => "00011100",1117 => "11111001",1118 => "01010101",1119 => "10010101",1120 => "01011011",1121 => "11100011",1122 => "10010001",1123 => "10001100",1124 => "00100010",1125 => "01101000",1126 => "00001010",1127 => "11100001",1128 => "01111000",1129 => "10010011",1130 => "01101010",1131 => "11101011",1132 => "10110101",1133 => "01100011",1134 => "00001010",1135 => "00111110",1136 => "01010001",1137 => "10010110",1138 => "11111000",1139 => "01101011",1140 => "10111100",1141 => "00111010",1142 => "01000010",1143 => "11011100",1144 => "01101010",1145 => "00110001",1146 => "00001111",1147 => "10110011",1148 => "00000011",1149 => "00101100",1150 => "10100000",1151 => "11111010",1152 => "00001100",1153 => "10010010",1154 => "00001001",1155 => "10101111",1156 => "01101010",1157 => "01101101",1158 => "10110101",1159 => "10010010",1160 => "10111110",1161 => "00001101",1162 => "00010100",1163 => "11001100",1164 => "01011110",1165 => "11101100",1166 => "01001110",1167 => "11011000",1168 => "11001101",1169 => "11101100",1170 => "10100111",1171 => "10100000",1172 => "01111101",1173 => "01101110",1174 => "10011001",1175 => "11011101",1176 => "00101101",1177 => "10001001",1178 => "01100001",1179 => "10100110",1180 => "10111100",1181 => "00011100",1182 => "11111001",1183 => "11100101",1184 => "10100011",1185 => "10010011",1186 => "01111111",1187 => "10010111",1188 => "11100111",1189 => "11101000",1190 => "11010100",1191 => "10000110",1192 => "01011101",1193 => "00110100",1194 => "01010110",1195 => "10110010",1196 => "01000011",1197 => "11111111",1198 => "11010100",1199 => "11001011",1200 => "10010001",1201 => "10010111",1202 => "00001001",1203 => "00100110",1204 => "11000100",1205 => "00100010",1206 => "11110011",1207 => "10101001",1208 => "10010010",1209 => "01100111",1210 => "10010010",1211 => "00100100",1212 => "11101011",1213 => "00001000",1214 => "10111111",1215 => "11011000",1216 => "10101001",1217 => "11101111",1218 => "11100100",1219 => "10000101",1220 => "11010100",1221 => "10000010",1222 => "01000101",1223 => "00111011",1224 => "11101010",1225 => "00110000",1226 => "10000010",1227 => "11001110",1228 => "01110111",1229 => "11000111",1230 => "10011001",1231 => "01001110",1232 => "10111111",1233 => "00000111",1234 => "11010010",1235 => "00011000",1236 => "11010111",1237 => "00011100",1238 => "01011000",1239 => "00010001",1240 => "11011000",1241 => "00000111",1242 => "11111001",1243 => "00110100",1244 => "01001110",1245 => "00101001",1246 => "01011000",1247 => "11100100",1248 => "01110110",1249 => "00011111",1250 => "11010101",1251 => "10001101",1252 => "00110100",1253 => "11001000",1254 => "01011011",1255 => "00101111",1256 => "11101111",1257 => "01000100",1258 => "01101001",1259 => "01000011",1260 => "01011001",1261 => "10000001",1262 => "10110100",1263 => "10111101",1264 => "11111010",1265 => "11100100",1266 => "10111111",1267 => "00100010",1268 => "10110111",1269 => "00101011",1270 => "11001110",1271 => "11001100",1272 => "00001101",1273 => "10011101",1274 => "01111000",1275 => "00101000",1276 => "00111100",1277 => "00001101",1278 => "10011101",1279 => "10101100",1280 => "00111101",1281 => "10110111",1282 => "11100110",1283 => "00101101",1284 => "11010111",1285 => "10000101",1286 => "11100000",1287 => "01110001",1288 => "11000111",1289 => "01011011",1290 => "00111100",1291 => "11111000",1292 => "00101010",1293 => "10110100",1294 => "00010001",1295 => "01100000",1296 => "01101000",1297 => "00110011",1298 => "10011010",1299 => "01011101",1300 => "11110101",1301 => "10010100",1302 => "00000000",1303 => "10101001",1304 => "00100100",1305 => "00000100",1306 => "10010110",1307 => "01100100",1308 => "11110011",1309 => "01101111",1310 => "01110010",1311 => "11110101",1312 => "11000110",1313 => "01100100",1314 => "10000101",1315 => "00101000",1316 => "10001100",1317 => "11001100",1318 => "01000010",1319 => "00000101",1320 => "11111010",1321 => "11011001",1322 => "01100110",1323 => "00011001",1324 => "01101110",1325 => "00001111",1326 => "11100111",1327 => "10010101",1328 => "11111101",1329 => "01010100",1330 => "10101010",1331 => "01101011",1332 => "11000001",1333 => "10001111",1334 => "11100001",1335 => "00111011",1336 => "10001000",1337 => "10111011",1338 => "01001110",1339 => "11011111",1340 => "11101100",1341 => "00100100",1342 => "10001111",1343 => "01000000",1344 => "11000110",1345 => "01111001",1346 => "10000111",1347 => "11110101",1348 => "11001101",1349 => "11100100",1350 => "00100101",1351 => "11000100",1352 => "10100111",1353 => "01010101",1354 => "11100111",1355 => "01110110",1356 => "00011001",1357 => "01011001",1358 => "00011111",1359 => "00100101",1360 => "01010101",1361 => "11000101",1362 => "01110101",1363 => "11010111",1364 => "10000100",1365 => "11100111",1366 => "11010000",1367 => "00011111",1368 => "11001010",1369 => "01100010",1370 => "11000100",1371 => "01111111",1372 => "01001101",1373 => "11101111",1374 => "00101111",1375 => "01010110",1376 => "01101100",1377 => "00100100",1378 => "01011110",1379 => "11101010",1380 => "01111000",1381 => "01010110",1382 => "00110101",1383 => "10000100",1384 => "11111001",1385 => "01000000",1386 => "01100000",1387 => "00010000",1388 => "10001101",1389 => "01101111",1390 => "01001001",1391 => "01110001",1392 => "00110001",1393 => "01110001",1394 => "10011110",1395 => "10001111",1396 => "01100011",1397 => "11100101",1398 => "00110010",1399 => "11110010",1400 => "10111000",1401 => "11111011",1402 => "11001100",1403 => "01001111",1404 => "00000111",1405 => "00011011",1406 => "00001101",1407 => "11010110",1408 => "10011011",1409 => "11101000",1410 => "10000011",1411 => "00000110",1412 => "11100110",1413 => "01111111",1414 => "01011111",1415 => "01010111",1416 => "01010111",1417 => "00110111",1418 => "10110000",1419 => "00100010",1420 => "11000111",1421 => "00100101",1422 => "10110100",1423 => "10110111",1424 => "10110101",1425 => "11011111",1426 => "10010000",1427 => "00010011",1428 => "11000111",1429 => "10110001",1430 => "00101101",1431 => "01001100",1432 => "00101011",1433 => "11001001",1434 => "00011010",1435 => "10111101",1436 => "00010010",1437 => "01101001",1438 => "01110110",1439 => "01011111",1440 => "00000101",1441 => "01001100",1442 => "11001111",1443 => "01001110",1444 => "11100011",1445 => "00111001",1446 => "01000010",1447 => "01100011",1448 => "01000011",1449 => "01010110",1450 => "10100111",1451 => "11101011",1452 => "01010010",1453 => "11010001",1454 => "01011010",1455 => "01111100",1456 => "11100001",1457 => "11001010",1458 => "11001111",1459 => "00111100",1460 => "11001011",1461 => "11000110",1462 => "11000000",1463 => "00000100",1464 => "01101000",1465 => "01110000",1466 => "00011010",1467 => "10001011",1468 => "01010100",1469 => "00110110",1470 => "01101100",1471 => "10100001",1472 => "11111010",1473 => "11101010",1474 => "10101001",1475 => "10011011",1476 => "11000111",1477 => "00000110",1478 => "10001000",1479 => "01110101",1480 => "11100001",1481 => "10110111",1482 => "00010010",1483 => "00010110",1484 => "11110000",1485 => "11111010",1486 => "11001110",1487 => "10001010",1488 => "11010001",1489 => "01001101",1490 => "10010010",1491 => "10101010",1492 => "10110110",1493 => "00110101",1494 => "10011101",1495 => "11111000",1496 => "00010010",1497 => "00010000",1498 => "11111001",1499 => "10100111",1500 => "11001101",1501 => "10100110",1502 => "10100000",1503 => "11110111",1504 => "11010000",1505 => "11100001",1506 => "01001100",1507 => "00110111",1508 => "00001100",1509 => "00100000",1510 => "11110111",1511 => "10011001",1512 => "10100111",1513 => "01111010",1514 => "11010111",1515 => "11011000",1516 => "01100100",1517 => "11110100",1518 => "11001101",1519 => "01001000",1520 => "10110111",1521 => "01010001",1522 => "01101011",1523 => "11000111",1524 => "10100010",1525 => "00110000",1526 => "10100000",1527 => "11011111",1528 => "11000011",1529 => "01011101",1530 => "10110001",1531 => "10101000",1532 => "11000110",1533 => "00110000",1534 => "11010001",1535 => "01101001",1536 => "11111111",1537 => "10110110",1538 => "11101101",1539 => "10010100",1540 => "11100111",1541 => "00010001",1542 => "00001001",1543 => "01111101",1544 => "10010100",1545 => "00000011",1546 => "10101111",1547 => "01010000",1548 => "01000100",1549 => "11000000",1550 => "10001000",1551 => "00111000",1552 => "10101011",1553 => "10000011",1554 => "10001100",1555 => "00100110",1556 => "11101100",1557 => "01000101",1558 => "00111110",1559 => "01100101",1560 => "11011110",1561 => "00000001",1562 => "10000010",1563 => "00111110",1564 => "01001101",1565 => "00101111",1566 => "11010011",1567 => "00100101",1568 => "10010001",1569 => "01000101",1570 => "10000000",1571 => "00111010",1572 => "01110110",1573 => "10010110",1574 => "11001000",1575 => "01011111",1576 => "10000011",1577 => "11001001",1578 => "00110110",1579 => "00001001",1580 => "00010011",1581 => "00011110",1582 => "11010110",1583 => "10111100",1584 => "00100101",1585 => "10101010",1586 => "01001011",1587 => "00101001",1588 => "01010100",1589 => "10011101",1590 => "00011110",1591 => "01000000",1592 => "10111000",1593 => "10010011",1594 => "00111110",1595 => "00110110",1596 => "01100010",1597 => "01100110",1598 => "01010001",1599 => "11001110",1600 => "01000000",1601 => "11111010",1602 => "10001110",1603 => "00010110",1604 => "00111111",1605 => "01111110",1606 => "10100001",1607 => "00111111",1608 => "01000111",1609 => "00111111",1610 => "10001001",1611 => "01100011",1612 => "00100111",1613 => "11011011",1614 => "10101100",1615 => "01000111",1616 => "01111001",1617 => "00001111",1618 => "00110001",1619 => "00101100",1620 => "10100000",1621 => "00011000",1622 => "11011101",1623 => "10101110",1624 => "00001110",1625 => "11000010",1626 => "00111010",1627 => "01010111",1628 => "01110011",1629 => "11011100",1630 => "10010101",1631 => "11111101",1632 => "11001111",1633 => "10110010",1634 => "11010101",1635 => "00111100",1636 => "01011111",1637 => "00010001",1638 => "00011011",1639 => "01100011",1640 => "11110100",1641 => "10101000",1642 => "01001010",1643 => "00011111",1644 => "00100110",1645 => "00000001",1646 => "11101010",1647 => "11000100",1648 => "01000011",1649 => "11011100",1650 => "11101110",1651 => "01010100",1652 => "10100110",1653 => "10001010",1654 => "00000111",1655 => "01110101",1656 => "11100000",1657 => "00001111",1658 => "11010100",1659 => "11101000",1660 => "01100000",1661 => "01011110",1662 => "10001101",1663 => "01111000",1664 => "11100101",1665 => "01010010",1666 => "11110000",1667 => "10011011",1668 => "00001101",1669 => "00100000",1670 => "11111111",1671 => "00000001",1672 => "00101001",1673 => "00011110",1674 => "00010100",1675 => "11000110",1676 => "10110011",1677 => "00001011",1678 => "10101001",1679 => "11011001",1680 => "01010101",1681 => "11111010",1682 => "11101110",1683 => "01011011",1684 => "00000001",1685 => "11011010",1686 => "10101101",1687 => "11101110",1688 => "00011110",1689 => "10001010",1690 => "11011000",1691 => "11010000",1692 => "00011111",1693 => "01110001",1694 => "01010110",1695 => "10111101",1696 => "10000001",1697 => "11000100",1698 => "10101111",1699 => "10011111",1700 => "00011111",1701 => "11001010",1702 => "10000111",1703 => "01000101",1704 => "11011111",1705 => "11110010",1706 => "11000101",1707 => "00111111",1708 => "00100001",1709 => "00010100",1710 => "11100101",1711 => "10101100",1712 => "10111100",1713 => "10110010",1714 => "01100111",1715 => "00011110",1716 => "11010011",1717 => "00011000",1718 => "11010100",1719 => "11100011",1720 => "11000001",1721 => "01111110",1722 => "10110001",1723 => "10001100",1724 => "01111101",1725 => "01010000",1726 => "00001011",1727 => "11010011",1728 => "10011101",1729 => "11110000",1730 => "01010111",1731 => "11111100",1732 => "00111001",1733 => "01001010",1734 => "10000011",1735 => "01100010",1736 => "01101011",1737 => "01100100",1738 => "11111111",1739 => "00111001",1740 => "10000001",1741 => "00011100",1742 => "10011110",1743 => "00010101",1744 => "01001000",1745 => "10111100",1746 => "00110101",1747 => "00110011",1748 => "11011010",1749 => "01000000",1750 => "01010001",1751 => "01000010",1752 => "10100011",1753 => "10000101",1754 => "11100011",1755 => "00100111",1756 => "10000101",1757 => "01010100",1758 => "00100100",1759 => "01101101",1760 => "10100011",1761 => "11101111",1762 => "00001000",1763 => "10000000",1764 => "10110010",1765 => "01111011",1766 => "10000100",1767 => "11001111",1768 => "01011111",1769 => "00101010",1770 => "00110110",1771 => "11001001",1772 => "00000001",1773 => "10011000",1774 => "11001000",1775 => "11001110",1776 => "10011011",1777 => "01111011",1778 => "01010110",1779 => "01100111",1780 => "10100000",1781 => "01100100",1782 => "11101011",1783 => "00111110",1784 => "11001101",1785 => "11001110",1786 => "00010001",1787 => "00101100",1788 => "00101000",1789 => "10110010",1790 => "11011010",1791 => "10011111",1792 => "00111111",1793 => "01000101",1794 => "10100010",1795 => "10001100",1796 => "01110111",1797 => "10011110",1798 => "10011011",1799 => "11001111",1800 => "10000101",1801 => "10101101",1802 => "01110111",1803 => "01000110",1804 => "01110001",1805 => "11010100",1806 => "00101111",1807 => "10011001",1808 => "00110101",1809 => "00101011",1810 => "00110101",1811 => "01110101",1812 => "00111001",1813 => "01100110",1814 => "10001010",1815 => "01100110",1816 => "11100010",1817 => "00001010",1818 => "00000101",1819 => "00000001",1820 => "00000111",1821 => "00110100",1822 => "11010001",1823 => "01111110",1824 => "00110111",1825 => "11000001",1826 => "11000011",1827 => "00011001",1828 => "00110010",1829 => "10101111",1830 => "11011000",1831 => "01001110",1832 => "10011011",1833 => "10101111",1834 => "00111110",1835 => "10110000",1836 => "11000110",1837 => "11110011",1838 => "01010110",1839 => "10111000",1840 => "11011001",1841 => "10101100",1842 => "11110101",1843 => "11110110",1844 => "01110001",1845 => "10100100",1846 => "10011001",1847 => "00001100",1848 => "01110001",1849 => "11100110",1850 => "01000010",1851 => "00100100",1852 => "01000110",1853 => "10110111",1854 => "00000111",1855 => "11101100",1856 => "00101111",1857 => "11111100",1858 => "01011000",1859 => "00001001",1860 => "11100111",1861 => "10000000",1862 => "00111111",1863 => "00010111",1864 => "00001101",1865 => "10000110",1866 => "10000110",1867 => "01011110",1868 => "01110110",1869 => "00001111",1870 => "10001111",1871 => "00101101",1872 => "10101100",1873 => "11010111",1874 => "11111000",1875 => "00110011",1876 => "00110111",1877 => "10010010",1878 => "00001001",1879 => "01001100",1880 => "01110100",1881 => "11111010",1882 => "10100100",1883 => "01100110",1884 => "11010011",1885 => "11100001",1886 => "01011010",1887 => "01001101",1888 => "00110111",1889 => "01010010",1890 => "11101000",1891 => "00000011",1892 => "00010000",1893 => "01011111",1894 => "01001001",1895 => "01100101",1896 => "11001101",1897 => "11001011",1898 => "10010000",1899 => "00011011",1900 => "10111111",1901 => "10010011",1902 => "00100001",1903 => "00101101",1904 => "10001011",1905 => "01001111",1906 => "00011001",1907 => "01111110",1908 => "01110110",1909 => "11010111",1910 => "10010100",1911 => "10101001",1912 => "00111010",1913 => "00001100",1914 => "00010110",1915 => "00111101",1916 => "11000011",1917 => "11110101",1918 => "11001100",1919 => "10000110",1920 => "11010100",1921 => "10110010",1922 => "10101001",1923 => "11100001",1924 => "01100001",1925 => "01100010",1926 => "10100111",1927 => "00111010",1928 => "10111101",1929 => "00010011",1930 => "00110101",1931 => "11011101",1932 => "11011111",1933 => "01010010",1934 => "11001111",1935 => "11100100",1936 => "11111110",1937 => "11100000",1938 => "11110101",1939 => "11011100",1940 => "11010110",1941 => "10101111",1942 => "10111101",1943 => "10101111",1944 => "01001101",1945 => "10010110",1946 => "01011001",1947 => "11111001",1948 => "10101100",1949 => "10100011",1950 => "01010110",1951 => "00111000",1952 => "00100001",1953 => "00110110",1954 => "10000011",1955 => "00101100",1956 => "01100111",1957 => "01111000",1958 => "10010000",1959 => "10110100",1960 => "01111110",1961 => "00001011",1962 => "10101010",1963 => "01001111",1964 => "10011010",1965 => "00010000",1966 => "00111000",1967 => "00101010",1968 => "10100010",1969 => "11111110",1970 => "11101111",1971 => "10011100",1972 => "11111011",1973 => "01100101",1974 => "00110110",1975 => "10001011",1976 => "10010000",1977 => "00110100",1978 => "11001101",1979 => "11111000",1980 => "11011010",1981 => "01001000",1982 => "11101000",1983 => "00101000",1984 => "01101110",1985 => "00111111",1986 => "01010010",1987 => "10100010",1988 => "01001101",1989 => "10101110",1990 => "10111010",1991 => "01001010",1992 => "11000100",1993 => "01001000",1994 => "01000001",1995 => "00010000",1996 => "01100001",1997 => "00001010",1998 => "10010001",1999 => "10001110",2000 => "01001110",2001 => "11100101",2002 => "10100001",2003 => "00110000",2004 => "10101100",2005 => "00010011",2006 => "01110000",2007 => "11010101",2008 => "11001111",2009 => "11011100",2010 => "10011101",2011 => "11110100",2012 => "01010111",2013 => "00001100",2014 => "01110101",2015 => "10100010",2016 => "10110111",2017 => "10010011",2018 => "00010100",2019 => "01000010",2020 => "10110010",2021 => "11100110",2022 => "10101011",2023 => "00000011",2024 => "01001111",2025 => "00011010",2026 => "00110011",2027 => "10100111",2028 => "10100001",2029 => "00011111",2030 => "11101101",2031 => "01010000",2032 => "10011101",2033 => "11001000",2034 => "10001011",2035 => "00011100",2036 => "00110100",2037 => "11101010",2038 => "11100100",2039 => "00100100",2040 => "01010101",2041 => "00111000",2042 => "11111110",2043 => "00111001",2044 => "11011100",2045 => "10100111",2046 => "11011010",2047 => "10111111",2048 => "01110110",2049 => "11110101",2050 => "00110110",2051 => "10101001",2052 => "11011001",2053 => "01010100",2054 => "01001001",2055 => "10001110",2056 => "01010100",2057 => "11010010",2058 => "10000010",2059 => "10011100",2060 => "11101000",2061 => "11000011",2062 => "11110010",2063 => "01001010",2064 => "11011000",2065 => "00010000",2066 => "01010010",2067 => "01001000",2068 => "11010000",2069 => "11111011",2070 => "10110001",2071 => "01010000",2072 => "00101001",2073 => "00011000",2074 => "00011011",2075 => "10010100",2076 => "10010001",2077 => "01100011",2078 => "01001010",2079 => "11001100",2080 => "00001011",2081 => "10000101",2082 => "00100111",2083 => "10010111",2084 => "01000101",2085 => "11110001",2086 => "11011000",2087 => "01000111",2088 => "11110110",2089 => "00110100",2090 => "11000011",2091 => "10100000",2092 => "01011101",2093 => "01101101",2094 => "11101010",2095 => "01000011",2096 => "11101101",2097 => "01101010",2098 => "01111000",2099 => "11110100",2100 => "10010110",2101 => "00101111",2102 => "00100000",2103 => "10110011",2104 => "10100001",2105 => "01101000",2106 => "01110000",2107 => "00011000",2108 => "00011001",2109 => "10110101",2110 => "00101011",2111 => "00001110",2112 => "01100110",2113 => "10001000",2114 => "11000101",2115 => "01001001",2116 => "10101111",2117 => "00000111",2118 => "01101111",2119 => "00011010",2120 => "10001100",2121 => "11100100",2122 => "10100010",2123 => "10100110",2124 => "01000111",2125 => "00001000",2126 => "11001111",2127 => "10011011",2128 => "10100100",2129 => "00111010",2130 => "10010110",2131 => "00101100",2132 => "10000110",2133 => "11110011",2134 => "01011010",2135 => "10101011",2136 => "10110111",2137 => "01101110",2138 => "11011010",2139 => "10001000",2140 => "01100110",2141 => "10010000",2142 => "11100000",2143 => "01000111",2144 => "00001001",2145 => "11010101",2146 => "11100110",2147 => "10011001",2148 => "00000010",2149 => "11000100",2150 => "01101111",2151 => "11011101",2152 => "01001100",2153 => "01111001",2154 => "10100110",2155 => "01111111",2156 => "10000011",2157 => "01010111",2158 => "11011110",2159 => "00111101",2160 => "01110101",2161 => "00011100",2162 => "11011011",2163 => "00000001",2164 => "00001101",2165 => "01011011",2166 => "00010011",2167 => "01000101",2168 => "01000010",2169 => "01001110",2170 => "00101101",2171 => "01010111",2172 => "11110100",2173 => "01000100",2174 => "11100000",2175 => "10000010",2176 => "10101001",2177 => "10110110",2178 => "11111000",2179 => "10101011",2180 => "10000100",2181 => "01101110",2182 => "00001000",2183 => "10101101",2184 => "01100000",2185 => "00001111",2186 => "01010001",2187 => "00010001",2188 => "01100111",2189 => "11111011",2190 => "00000110",2191 => "01110001",2192 => "10001111",2193 => "10111000",2194 => "01100011",2195 => "00110000",2196 => "10110110",2197 => "00111000",2198 => "00101110",2199 => "00011011",2200 => "00100100",2201 => "10110101",2202 => "00011001",2203 => "10001100",2204 => "00010100",2205 => "01011011",2206 => "00100010",2207 => "10111111",2208 => "01110000",2209 => "11111010",2210 => "11000110",2211 => "11001010",2212 => "10001000",2213 => "10001100",2214 => "01001101",2215 => "11011011",2216 => "10110110",2217 => "01001011",2218 => "00111011",2219 => "10000111",2220 => "11111010",2221 => "01101001",2222 => "11010101",2223 => "01011010",2224 => "10010001",2225 => "00010101",2226 => "10000001",2227 => "11000010",2228 => "10011110",2229 => "00111101",2230 => "10110000",2231 => "00100011",2232 => "10100110",2233 => "00101101",2234 => "10010010",2235 => "11001101",2236 => "11001110",2237 => "00110010",2238 => "01101010",2239 => "11001011",2240 => "11101110",2241 => "01111101",2242 => "00001011",2243 => "11100100",2244 => "00000000",2245 => "11111100",2246 => "01110110",2247 => "00000010",2248 => "01010000",2249 => "11010111",2250 => "01000110",2251 => "10011000",2252 => "01110001",2253 => "10110000",2254 => "00000000",2255 => "11010110",2256 => "10000111",2257 => "11110001",2258 => "11011101",2259 => "00010011",2260 => "11001000",2261 => "00000010",2262 => "11001010",2263 => "10001111",2264 => "10110100",2265 => "00111010",2266 => "10111001",2267 => "11000011",2268 => "10010000",2269 => "01101000",2270 => "10100010",2271 => "01011001",2272 => "01011110",2273 => "11101100",2274 => "11011010",2275 => "10011111",2276 => "01100110",2277 => "10011110",2278 => "10111100",2279 => "01010010",2280 => "10100111",2281 => "00110001",2282 => "11010110",2283 => "01010000",2284 => "00000100",2285 => "10011001",2286 => "10011000",2287 => "01001001",2288 => "11010101",2289 => "01010111",2290 => "01001001",2291 => "01100100",2292 => "00100011",2293 => "01111000",2294 => "10010110",2295 => "00001001",2296 => "10000110",2297 => "01101111",2298 => "01100101",2299 => "10000011",2300 => "10111000",2301 => "11110111",2302 => "01010000",2303 => "11111111",2304 => "11101011",2305 => "10010101",2306 => "00110011",2307 => "00110001",2308 => "01011000",2309 => "11000110",2310 => "10011001",2311 => "10010011",2312 => "10101010",2313 => "10000101",2314 => "01111001",2315 => "00011011",2316 => "00011000",2317 => "00011011",2318 => "10110101",2319 => "00101110",2320 => "00001001",2321 => "00010110",2322 => "00111110",2323 => "01011111",2324 => "00010000",2325 => "11011011",2326 => "11000010",2327 => "00111110",2328 => "00110111",2329 => "00111101",2330 => "01101010",2331 => "10001100",2332 => "00100010",2333 => "10000001",2334 => "11001010",2335 => "10011110",2336 => "10010010",2337 => "11101001",2338 => "01101100",2339 => "01000001",2340 => "01011100",2341 => "11100110",2342 => "10001001",2343 => "11101000",2344 => "11110101",2345 => "01001101",2346 => "11011111",2347 => "11011010",2348 => "10001011",2349 => "11111100",2350 => "10000110",2351 => "01010000",2352 => "01111011",2353 => "00101011",2354 => "10101101",2355 => "11111011",2356 => "01011001",2357 => "10101010",2358 => "01100000",2359 => "01101001",2360 => "00101000",2361 => "10110011",2362 => "11110011",2363 => "11111010",2364 => "10000111",2365 => "00110111",2366 => "01100000",2367 => "00011010",2368 => "00011100",2369 => "01101101",2370 => "10000101",2371 => "00000111",2372 => "10110110",2373 => "01010101",2374 => "01010000",2375 => "00101111",2376 => "01010101",2377 => "11100000",2378 => "10011100",2379 => "01000111",2380 => "11011100",2381 => "01100010",2382 => "01011110",2383 => "01110100",2384 => "00110111",2385 => "01011010",2386 => "01101011",2387 => "11101001",2388 => "11010011",2389 => "01011011",2390 => "10100101",2391 => "11110110",2392 => "10001001",2393 => "01100110",2394 => "11110011",2395 => "00000110",2396 => "01001110",2397 => "11111110",2398 => "01110100",2399 => "11100110",2400 => "11000110",2401 => "01100100",2402 => "00000000",2403 => "11011111",2404 => "01010010",2405 => "11011000",2406 => "10110010",2407 => "00001101",2408 => "01111110",2409 => "00011001",2410 => "11100001",2411 => "10010110",2412 => "11110100",2413 => "01011001",2414 => "01111110",2415 => "10100011",2416 => "01001010",2417 => "01001000",2418 => "10010101",2419 => "10101100",2420 => "11010111",2421 => "00110001",2422 => "11010011",2423 => "11011101",2424 => "01010110",2425 => "10001000",2426 => "11110111",2427 => "00011100",2428 => "10011110",2429 => "00001101",2430 => "11100101",2431 => "10101001",2432 => "01111001",2433 => "10110001",2434 => "11101100",2435 => "00010000",2436 => "10000111",2437 => "11101101",2438 => "00100011",2439 => "00011010",2440 => "11101111",2441 => "10101000",2442 => "10001101",2443 => "10001101",2444 => "11010000",2445 => "11010000",2446 => "00010010",2447 => "10100111",2448 => "11001100",2449 => "01111101",2450 => "10111101",2451 => "11100001",2452 => "11111100",2453 => "00111100",2454 => "00100100",2455 => "10100101",2456 => "10000101",2457 => "01100000",2458 => "00111100",2459 => "00101100",2460 => "11000111",2461 => "11101011",2462 => "10100111",2463 => "01001000",2464 => "10110100",2465 => "10000001",2466 => "11010010",2467 => "10000110",2468 => "10010110",2469 => "11000001",2470 => "00010001",2471 => "10100101",2472 => "11000110",2473 => "01011110",2474 => "10100010",2475 => "00011010",2476 => "01111111",2477 => "11001111",2478 => "00010110",2479 => "10010100",2480 => "11001011",2481 => "01001000",2482 => "01101001",2483 => "10000001",2484 => "11111111",2485 => "00101001",2486 => "10010010",2487 => "01111011",2488 => "11111110",2489 => "01110101",2490 => "10011011",2491 => "01001110",2492 => "11000010",2493 => "10110010",2494 => "10010011",2495 => "01100100",2496 => "11011000",2497 => "11110110",2498 => "11011111",2499 => "10110000",2500 => "10110110",2501 => "11010000",2502 => "10101111",2503 => "00111111",2504 => "01100110",2505 => "10110111",2506 => "01011101",2507 => "11101110",2508 => "01000110",2509 => "10001101",2510 => "00010000",2511 => "00001110",2512 => "01110100",2513 => "11100010",2514 => "11011011",2515 => "10111110",2516 => "10011111",2517 => "11111101",2518 => "00011101",2519 => "10111000",2520 => "00111110",2521 => "00001011",2522 => "01100010",2523 => "10000011",2524 => "10011000",2525 => "01001100",2526 => "00100000",2527 => "00001111",2528 => "11110000",2529 => "01001011",2530 => "11001001",2531 => "11010010",2532 => "10110000",2533 => "00111110",2534 => "10110110",2535 => "01101001",2536 => "11101110",2537 => "11100001",2538 => "11011010",2539 => "11011101",2540 => "00001010",2541 => "11000011",2542 => "00000101",2543 => "00101101",2544 => "10100001",2545 => "11001101",2546 => "00110100",2547 => "01010101",2548 => "01100100",2549 => "01001111",2550 => "10100110",2551 => "00100110",2552 => "11101011",2553 => "01110111",2554 => "01000000",2555 => "10111110",2556 => "11101000",2557 => "11100000",2558 => "01111100",2559 => "11110011",2560 => "10010011",2561 => "00000010",2562 => "00000011",2563 => "10010110",2564 => "01011100",2565 => "00100111",2566 => "01001111",2567 => "00100111",2568 => "01100000",2569 => "10010001",2570 => "10010110",2571 => "01000000",2572 => "01110010",2573 => "11001100",2574 => "11101100",2575 => "01101001",2576 => "01110010",2577 => "10100100",2578 => "11001011",2579 => "00110000",2580 => "11010001",2581 => "11110010",2582 => "01000000",2583 => "11110110",2584 => "00000111",2585 => "10011000",2586 => "01011110",2587 => "10111101",2588 => "10000001",2589 => "01110111",2590 => "11011010",2591 => "11001001",2592 => "00110111",2593 => "10101100",2594 => "10101110",2595 => "00111101",2596 => "01101010",2597 => "00011011",2598 => "01001000",2599 => "10110110",2600 => "10011001",2601 => "00001011",2602 => "01010001",2603 => "10101100",2604 => "11101001",2605 => "10011010",2606 => "10110111",2607 => "00110010",2608 => "01000010",2609 => "11100000",2610 => "10110000",2611 => "10010101",2612 => "00001111",2613 => "10101100",2614 => "10100001",2615 => "00111100",2616 => "10000000",2617 => "01011010",2618 => "10110011",2619 => "11111010",2620 => "01100101",2621 => "00110001",2622 => "10110110",2623 => "01001101",2624 => "11010111",2625 => "11101110",2626 => "00101101",2627 => "00001010",2628 => "01011001",2629 => "11101000",2630 => "01010101",2631 => "10111100",2632 => "00001101",2633 => "00010011",2634 => "11100100",2635 => "10110110",2636 => "00011011",2637 => "01011100",2638 => "01011010",2639 => "11111000",2640 => "10011010",2641 => "00010111",2642 => "11000111",2643 => "10100100",2644 => "00011000",2645 => "11110001",2646 => "01000110",2647 => "01011110",2648 => "00001101",2649 => "10010110",2650 => "10100000",2651 => "01100100",2652 => "01100100",2653 => "01111110",2654 => "00000101",2655 => "01100101",2656 => "11100001",2657 => "11101100",2658 => "00110101",2659 => "01111101",2660 => "10101001",2661 => "00001000",2662 => "00010101",2663 => "00011101",2664 => "00001010",2665 => "11000010",2666 => "00011110",2667 => "01110001",2668 => "00000001",2669 => "10010100",2670 => "01000001",2671 => "00010110",2672 => "11011011",2673 => "00100100",2674 => "00011000",2675 => "10111011",2676 => "10111110",2677 => "01101010",2678 => "00001010",2679 => "11001010",2680 => "00000000",2681 => "00001001",2682 => "01000001",2683 => "10101001",2684 => "01101000",2685 => "01010100",2686 => "01010100",2687 => "00100001",2688 => "00110011",2689 => "11100101",2690 => "10101010",2691 => "11000110",2692 => "00001010",2693 => "01010001",2694 => "01010000",2695 => "10110101",2696 => "01110010",2697 => "01000001",2698 => "00001101",2699 => "11000010",2700 => "10010001",2701 => "00100111",2702 => "00010101",2703 => "01011000",2704 => "11101001",2705 => "10001010",2706 => "11000001",2707 => "01000111",2708 => "00000110",2709 => "11101001",2710 => "01100000",2711 => "10011011",2712 => "11001101",2713 => "10111110",2714 => "11011111",2715 => "11110010",2716 => "11000100",2717 => "11001111",2718 => "01010100",2719 => "01101100",2720 => "01011100",2721 => "11000100",2722 => "11100101",2723 => "00000111",2724 => "00110101",2725 => "10011111",2726 => "00011100",2727 => "00000010",2728 => "01100100",2729 => "00011111",2730 => "00011110",2731 => "01101000",2732 => "01001100",2733 => "01110111",2734 => "10000011",2735 => "11011100",2736 => "00001101",2737 => "00101010",2738 => "01001110",2739 => "10101101",2740 => "10001101",2741 => "00001101",2742 => "11110000",2743 => "01000011",2744 => "01101000",2745 => "10001000",2746 => "11000001",2747 => "01101011",2748 => "11010011",2749 => "00000001",2750 => "10100010",2751 => "00100110",2752 => "10110111",2753 => "01011101",2754 => "11111110",2755 => "00001011",2756 => "11110100",2757 => "10101011",2758 => "10101011",2759 => "01100110",2760 => "10110111",2761 => "10011001",2762 => "01110011",2763 => "11111110",2764 => "00111111",2765 => "00111000",2766 => "10011110",2767 => "11100010",2768 => "00001001",2769 => "01111010",2770 => "01001110",2771 => "10111110",2772 => "00010000",2773 => "10001100",2774 => "11001011",2775 => "10001110",2776 => "11011000",2777 => "00111001",2778 => "01111000",2779 => "11111101",2780 => "11111000",2781 => "11001100",2782 => "00010101",2783 => "01110101",2784 => "01101011",2785 => "00111000",2786 => "10110001",2787 => "11000110",2788 => "10011010",2789 => "00000011",2790 => "01011100",2791 => "10100110",2792 => "00111101",2793 => "01011101",2794 => "11000100",2795 => "10111101",2796 => "00110000",2797 => "10100100",2798 => "10111101",2799 => "11100111",2800 => "10010000",2801 => "10100110",2802 => "00110111",2803 => "11000001",2804 => "11000111",2805 => "10010000",2806 => "01000000",2807 => "00111000",2808 => "01110110",2809 => "11101110",2810 => "00000100",2811 => "10101100",2812 => "01101000",2813 => "01001011",2814 => "10010111",2815 => "11011010",2816 => "10000010",2817 => "00100001",2818 => "10000010",2819 => "01010001",2820 => "11011101",2821 => "00110001",2822 => "01011111",2823 => "00110111",2824 => "01000011",2825 => "00101100",2826 => "11001010",2827 => "01101110",2828 => "00100100",2829 => "10100011",2830 => "10011111",2831 => "10101101",2832 => "10011011",2833 => "11011110",2834 => "00100010",2835 => "11011011",2836 => "10000101",2837 => "10101000",2838 => "11000100",2839 => "00011011",2840 => "01011011",2841 => "10101000",2842 => "00011010",2843 => "10110010",2844 => "01100011",2845 => "01010110",2846 => "11101011",2847 => "11000111",2848 => "10010111",2849 => "10000000",2850 => "11100011",2851 => "01110101",2852 => "00100001",2853 => "10010011",2854 => "01010001",2855 => "00111011",2856 => "10110000",2857 => "11001111",2858 => "10001101",2859 => "01001111",2860 => "00000001",2861 => "11101001",2862 => "00011101",2863 => "11101000",2864 => "00101001",2865 => "11010111",2866 => "00100111",2867 => "01110110",2868 => "11001001",2869 => "10011010",2870 => "01101100",2871 => "11111001",2872 => "11111100",2873 => "01101000",2874 => "11001001",2875 => "11101001",2876 => "00110100",2877 => "11110111",2878 => "01100111",2879 => "11010100",2880 => "01011010",2881 => "11001010",2882 => "10010001",2883 => "11111000",2884 => "10000111",2885 => "10101001",2886 => "11001001",2887 => "10111101",2888 => "10000110",2889 => "10011101",2890 => "11101000",2891 => "11010101",2892 => "10011111",2893 => "00100101",2894 => "01010011",2895 => "10011011",2896 => "11010100",2897 => "11011101",2898 => "00111101",2899 => "01111011",2900 => "11011000",2901 => "11010011",2902 => "01100000",2903 => "00100001",2904 => "01101100",2905 => "00101001",2906 => "00001111",2907 => "10010110",2908 => "10010010",2909 => "01111000",2910 => "00000110",2911 => "01000101",2912 => "10010101",2913 => "01010010",2914 => "11010111",2915 => "01101100",2916 => "11010100",2917 => "01011011",2918 => "01111110",2919 => "01010011",2920 => "00110101",2921 => "00101110",2922 => "01111100",2923 => "11001000",2924 => "01010000",2925 => "00111100",2926 => "01111100",2927 => "11111001",2928 => "11110001",2929 => "10001001",2930 => "00011000",2931 => "00101010",2932 => "11101111",2933 => "01101011",2934 => "01111011",2935 => "11100111",2936 => "10110011",2937 => "10001111",2938 => "10001010",2939 => "11000000",2940 => "10010010",2941 => "01010010",2942 => "00110110",2943 => "01101111",2944 => "00101011",2945 => "11101011",2946 => "11101011",2947 => "10000000",2948 => "00010010",2949 => "11010010",2950 => "01100110",2951 => "10101010",2952 => "01100111",2953 => "11001011",2954 => "10100100",2955 => "00101011",2956 => "00001110",2957 => "10000000",2958 => "00010001",2959 => "11110111",2960 => "10001010",2961 => "00111111",2962 => "00010110",2963 => "10101011",2964 => "01100111",2965 => "11111101",2966 => "10011001",2967 => "10001111",2968 => "01011100",2969 => "01010100",2970 => "01101101",2971 => "00110111",2972 => "10101010",2973 => "11010100",2974 => "01110110",2975 => "11100010",2976 => "10100100",2977 => "01011101",2978 => "11000111",2979 => "01001111",2980 => "11100010",2981 => "00011100",2982 => "00111111",2983 => "01110011",2984 => "10101011",2985 => "11101001",2986 => "01010100",2987 => "10100010",2988 => "01101010",2989 => "11100011",2990 => "11001000",2991 => "10100101",2992 => "01001010",2993 => "00100001",2994 => "00011100",2995 => "11011101",2996 => "10000111",2997 => "01001010",2998 => "11110101",2999 => "11000011",3000 => "00000100",3001 => "01111111",3002 => "11011110",3003 => "01000100",3004 => "01111000",3005 => "01111111",3006 => "00011010",3007 => "01100110",3008 => "10010011",3009 => "10111010",3010 => "00010111",3011 => "11111011",3012 => "10111011",3013 => "10101000",3014 => "10011000",3015 => "00110010",3016 => "11010111",3017 => "10101011",3018 => "11010110",3019 => "11000000",3020 => "01011100",3021 => "01010000",3022 => "00011111",3023 => "10100011",3024 => "01101101",3025 => "00010000",3026 => "00010000",3027 => "01001011",3028 => "10101111",3029 => "10110110",3030 => "01111010",3031 => "00000000",3032 => "10101101",3033 => "01001001",3034 => "11010110",3035 => "00111001",3036 => "00011100",3037 => "00110110",3038 => "10110010",3039 => "10100101",3040 => "10001110",3041 => "11110000",3042 => "10101100",3043 => "10000111",3044 => "00011011",3045 => "00000011",3046 => "11110011",3047 => "01101100",3048 => "11110011",3049 => "10110100",3050 => "10011001",3051 => "10001111",3052 => "10010000",3053 => "10000011",3054 => "10011110",3055 => "00111010",3056 => "01101110",3057 => "11100100",3058 => "01001100",3059 => "00010110",3060 => "11111110",3061 => "01010111",3062 => "10001110",3063 => "01100100",3064 => "01110000",3065 => "01010011",3066 => "10001101",3067 => "00110100",3068 => "01110110",3069 => "00101011",3070 => "01110000",3071 => "00111111",3072 => "10101010",3073 => "10000010",3074 => "00110100",3075 => "01101000",3076 => "10100100",3077 => "00110010",3078 => "11011010",3079 => "11011010",3080 => "10010110",3081 => "01111001",3082 => "01001101",3083 => "10011101",3084 => "00101110",3085 => "11100011",3086 => "00110110",3087 => "01111010",3088 => "00110110",3089 => "11011100",3090 => "11101100",3091 => "01010001",3092 => "00111110",3093 => "00110010",3094 => "10101010",3095 => "11111011",3096 => "11011000",3097 => "00000011",3098 => "10010011",3099 => "01101111",3100 => "11111011",3101 => "11001000",3102 => "10010000",3103 => "01011011",3104 => "00001000",3105 => "00001111",3106 => "10011110",3107 => "01100101",3108 => "10111100",3109 => "01001100",3110 => "00011100",3111 => "11001011",3112 => "01011110",3113 => "00011111",3114 => "11101101",3115 => "00111111",3116 => "01111101",3117 => "00110101",3118 => "10100100",3119 => "01000111",3120 => "01101101",3121 => "11111100",3122 => "10110101",3123 => "10101010",3124 => "10010011",3125 => "10100010",3126 => "00011010",3127 => "00100101",3128 => "10000100",3129 => "10010011",3130 => "01001010",3131 => "01101001",3132 => "01010011",3133 => "01111101",3134 => "00010110",3135 => "11011001",3136 => "10110110",3137 => "01100000",3138 => "10100011",3139 => "11101101",3140 => "10100001",3141 => "10100101",3142 => "01101011",3143 => "11010111",3144 => "00110001",3145 => "01001011",3146 => "11100000",3147 => "11010110",3148 => "01100100",3149 => "10011000",3150 => "11000111",3151 => "00110101",3152 => "01111111",3153 => "11010101",3154 => "01011011",3155 => "00010110",3156 => "10101101",3157 => "00101110",3158 => "01111011",3159 => "10100111",3160 => "10001110",3161 => "10111100",3162 => "01010111",3163 => "01011001",3164 => "01110010",3165 => "01101101",3166 => "00101000",3167 => "00000111",3168 => "10011000",3169 => "01110100",3170 => "10010001",3171 => "01100100",3172 => "10010101",3173 => "11101000",3174 => "00010111",3175 => "11010000",3176 => "00010100",3177 => "11100100",3178 => "00111011",3179 => "01010101",3180 => "11111001",3181 => "11101000",3182 => "01110010",3183 => "00001111",3184 => "11000110",3185 => "11000010",3186 => "00110011",3187 => "11000100",3188 => "10001111",3189 => "01101111",3190 => "00110011",3191 => "00011111",3192 => "11010111",3193 => "01001100",3194 => "11101110",3195 => "00010001",3196 => "01011001",3197 => "00110110",3198 => "00001101",3199 => "10100110",3200 => "11111101",3201 => "00010011",3202 => "01010110",3203 => "10101110",3204 => "10011010",3205 => "10011101",3206 => "01101011",3207 => "11000011",3208 => "11010110",3209 => "11001001",3210 => "00111001",3211 => "11111000",3212 => "01000010",3213 => "01110111",3214 => "00001101",3215 => "00100010",3216 => "00000011",3217 => "10100100",3218 => "00101000",3219 => "01010101",3220 => "10101001",3221 => "00001000",3222 => "01000001",3223 => "01101000",3224 => "00010010",3225 => "01001010",3226 => "11011011",3227 => "01111000",3228 => "00001011",3229 => "01000100",3230 => "01011111",3231 => "10111010",3232 => "10100110",3233 => "00000110",3234 => "01111001",3235 => "11110110",3236 => "11110110",3237 => "01011101",3238 => "10100100",3239 => "00100110",3240 => "01001000",3241 => "00011010",3242 => "11000101",3243 => "10110111",3244 => "01110000",3245 => "00010001",3246 => "01010100",3247 => "01110010",3248 => "11111110",3249 => "01110001",3250 => "10110011",3251 => "00010010",3252 => "10110011",3253 => "00001001",3254 => "00101110",3255 => "10000100",3256 => "11110010",3257 => "10100001",3258 => "00011001",3259 => "00100000",3260 => "01111111",3261 => "10011010",3262 => "01101110",3263 => "11101101",3264 => "00110110",3265 => "01111111",3266 => "01010100",3267 => "01010110",3268 => "00100100",3269 => "00001111",3270 => "01011011",3271 => "01011010",3272 => "00110011",3273 => "10000100",3274 => "11011011",3275 => "00011011",3276 => "01011110",3277 => "01101000",3278 => "00001001",3279 => "01110110",3280 => "01110110",3281 => "11010100",3282 => "01000110",3283 => "01111000",3284 => "01001010",3285 => "11000001",3286 => "10000011",3287 => "10010010",3288 => "00001110",3289 => "00010111",3290 => "01011110",3291 => "01010101",3292 => "00000100",3293 => "00010011",3294 => "10110100",3295 => "01100110",3296 => "00110110",3297 => "10100010",3298 => "11110100",3299 => "01110111",3300 => "01010001",3301 => "01101101",3302 => "01011101",3303 => "01110001",3304 => "11011000",3305 => "11101100",3306 => "01000100",3307 => "11000001",3308 => "00101111",3309 => "10110111",3310 => "10100001",3311 => "00110000",3312 => "00101010",3313 => "00011000",3314 => "11110001",3315 => "00000001",3316 => "01011000",3317 => "00101100",3318 => "00000111",3319 => "11000110",3320 => "01010001",3321 => "00100010",3322 => "11000000",3323 => "00101101",3324 => "00000001",3325 => "11111011",3326 => "10010011",3327 => "01101110",3328 => "00101011",3329 => "00110111",3330 => "11101001",3331 => "01100001",3332 => "10011101",3333 => "11110100",3334 => "11101011",3335 => "01111001",3336 => "11011111",3337 => "11100100",3338 => "11011011",3339 => "01100001",3340 => "10001110",3341 => "00000011",3342 => "10001111",3343 => "11010011",3344 => "11101100",3345 => "11010011",3346 => "00111001",3347 => "11111001",3348 => "11110100",3349 => "01000101",3350 => "01111100",3351 => "10000110",3352 => "10000111",3353 => "10101000",3354 => "00111111",3355 => "11111100",3356 => "00000111",3357 => "10111101",3358 => "00011001",3359 => "10100111",3360 => "01111100",3361 => "01001111",3362 => "01001111",3363 => "00010001",3364 => "10011011",3365 => "00001011",3366 => "10000001",3367 => "11110011",3368 => "00000011",3369 => "01000011",3370 => "10110011",3371 => "01111111",3372 => "10111001",3373 => "00001101",3374 => "11011111",3375 => "10010000",3376 => "11111011",3377 => "11011101",3378 => "00010101",3379 => "10100001",3380 => "11110010",3381 => "11001000",3382 => "11100101",3383 => "10101101",3384 => "10011000",3385 => "11010101",3386 => "00011011",3387 => "01100011",3388 => "11010101",3389 => "10010000",3390 => "10001011",3391 => "11011111",3392 => "10110011",3393 => "00001110",3394 => "00011101",3395 => "11110111",3396 => "10011010",3397 => "10101010",3398 => "11100010",3399 => "00111101",3400 => "01001011",3401 => "10011100",3402 => "00111101",3403 => "00001110",3404 => "11001011",3405 => "01001010",3406 => "01000110",3407 => "00111010",3408 => "00000001",3409 => "11000001",3410 => "11111011",3411 => "10000011",3412 => "11101111",3413 => "10010111",3414 => "00101000",3415 => "01100011",3416 => "10010101",3417 => "00100011",3418 => "00111111",3419 => "00111111",3420 => "11010000",3421 => "01110001",3422 => "01101011",3423 => "10000011",3424 => "11001101",3425 => "01100001",3426 => "11111000",3427 => "10010101",3428 => "01101100",3429 => "11100010",3430 => "01001100",3431 => "00101000",3432 => "10100011",3433 => "11101001",3434 => "00100110",3435 => "10001111",3436 => "11010001",3437 => "00001110",3438 => "00101010",3439 => "01101000",3440 => "10110011",3441 => "10110100",3442 => "10101011",3443 => "11100001",3444 => "10100011",3445 => "11101101",3446 => "11011100",3447 => "01101000",3448 => "01000000",3449 => "10010010",3450 => "00000101",3451 => "11111011",3452 => "00010011",3453 => "11100100",3454 => "01010101",3455 => "11010000",3456 => "11000100",3457 => "10101010",3458 => "01110111",3459 => "01100010",3460 => "00110010",3461 => "00101111",3462 => "00111001",3463 => "01100010",3464 => "00001101",3465 => "11110011",3466 => "11100010",3467 => "01001001",3468 => "10000001",3469 => "00100100",3470 => "01110010",3471 => "10110101",3472 => "11111001",3473 => "00101011",3474 => "10001101",3475 => "11011100",3476 => "01001100",3477 => "11111011",3478 => "10110100",3479 => "11101101",3480 => "11000111",3481 => "10111011",3482 => "00110101",3483 => "01100010",3484 => "10101100",3485 => "10001010",3486 => "11010111",3487 => "11111011",3488 => "01000101",3489 => "11011000",3490 => "10101110",3491 => "01011011",3492 => "01100111",3493 => "11111000",3494 => "00000010",3495 => "10100110",3496 => "00110000",3497 => "11100001",3498 => "01010110",3499 => "00001111",3500 => "11010111",3501 => "01000110",3502 => "11111110",3503 => "11011011",3504 => "10101001",3505 => "11000001",3506 => "11111101",3507 => "10100101",3508 => "01001011",3509 => "00110010",3510 => "01011011",3511 => "01010000",3512 => "00100110",3513 => "10110011",3514 => "01110000",3515 => "10101101",3516 => "10011011",3517 => "11000010",3518 => "00110100",3519 => "10001111",3520 => "00000110",3521 => "11011110",3522 => "11001011",3523 => "11111011",3524 => "10111110",3525 => "10011101",3526 => "01111000",3527 => "10101000",3528 => "01010001",3529 => "01000010",3530 => "10011111",3531 => "11011111",3532 => "11111010",3533 => "11000010",3534 => "01010010",3535 => "00101101",3536 => "01001000",3537 => "00000100",3538 => "11000010",3539 => "00000100",3540 => "10111111",3541 => "00001011",3542 => "11010101",3543 => "11010101",3544 => "11010111",3545 => "11001011",3546 => "00001011",3547 => "01000110",3548 => "00001001",3549 => "01000111",3550 => "11100101",3551 => "11110011",3552 => "10100000",3553 => "11010100",3554 => "01111110",3555 => "01100010",3556 => "00110101",3557 => "10111111",3558 => "00010010",3559 => "10011111",3560 => "11011010",3561 => "11011111",3562 => "11011001",3563 => "11001011",3564 => "11110001",3565 => "10001000",3566 => "00010001",3567 => "00011110",3568 => "10011100",3569 => "01100110",3570 => "11110111",3571 => "01000001",3572 => "01011100",3573 => "10101001",3574 => "00001011",3575 => "11110000",3576 => "00111001",3577 => "11000111",3578 => "01010100",3579 => "00001101",3580 => "01011101",3581 => "01110011",3582 => "01111001",3583 => "10001011",3584 => "01001010",3585 => "10000000",3586 => "10101011",3587 => "10111111",3588 => "11100101",3589 => "11101000",3590 => "10001010",3591 => "10111011",3592 => "10011110",3593 => "11100111",3594 => "10101011",3595 => "11111001",3596 => "00011001",3597 => "10000111",3598 => "11110001",3599 => "10001001",3600 => "00000001",3601 => "00110000",3602 => "11010000",3603 => "00111110",3604 => "10000100",3605 => "00110101",3606 => "00110011",3607 => "01010100",3608 => "10010101",3609 => "01001001",3610 => "11111111",3611 => "11000110",3612 => "00111101",3613 => "01011001",3614 => "10010010",3615 => "10100101",3616 => "10001100",3617 => "10010100",3618 => "10011111",3619 => "11010000",3620 => "10110001",3621 => "01010101",3622 => "10000100",3623 => "00111111",3624 => "11000011",3625 => "00000000",3626 => "01100100",3627 => "00110000",3628 => "10101100",3629 => "00000101",3630 => "01110111",3631 => "01011000",3632 => "10011100",3633 => "00001111",3634 => "11100001",3635 => "10011110",3636 => "00011010",3637 => "00001101",3638 => "10010100",3639 => "01010101",3640 => "00110100",3641 => "10001111",3642 => "01110001",3643 => "10011010",3644 => "01110010",3645 => "11011011",3646 => "01101101",3647 => "10111100",3648 => "00110011",3649 => "00010010",3650 => "00010010",3651 => "01000001",3652 => "11101101",3653 => "10010000",3654 => "10111011",3655 => "00111011",3656 => "00100010",3657 => "11101001",3658 => "01111011",3659 => "11101100",3660 => "01111001",3661 => "00110111",3662 => "01110100",3663 => "10111100",3664 => "00111110",3665 => "10110000",3666 => "10100011",3667 => "00110001",3668 => "00101011",3669 => "00001010",3670 => "01011101",3671 => "11110111",3672 => "10001110",3673 => "10011001",3674 => "10010110",3675 => "11110011",3676 => "00100111",3677 => "11000001",3678 => "00111101",3679 => "00000011",3680 => "11100101",3681 => "11001001",3682 => "11011111",3683 => "11100010",3684 => "01110100",3685 => "00111001",3686 => "00010000",3687 => "00000111",3688 => "00000100",3689 => "01110010",3690 => "00000111",3691 => "10011000",3692 => "10001001",3693 => "00010000",3694 => "11111110",3695 => "01000110",3696 => "00000010",3697 => "00100110",3698 => "00000111",3699 => "00001001",3700 => "00110010",3701 => "11111001",3702 => "10110111",3703 => "11011111",3704 => "01010101",3705 => "11100010",3706 => "10011010",3707 => "00001011",3708 => "00001001",3709 => "01010111",3710 => "10001101",3711 => "11101100",3712 => "01110111",3713 => "10001011",3714 => "11110101",3715 => "00101010",3716 => "11000101",3717 => "01010110",3718 => "11100010",3719 => "01011010",3720 => "10101000",3721 => "10011001",3722 => "11101001",3723 => "01101011",3724 => "01010010",3725 => "10110110",3726 => "11111110",3727 => "11110101",3728 => "01010100",3729 => "10010001",3730 => "10110110",3731 => "01010100",3732 => "00001000",3733 => "00010100",3734 => "00100000",3735 => "00011000",3736 => "11011010",3737 => "01011011",3738 => "00010001",3739 => "00000001",3740 => "01011111",3741 => "10101110",3742 => "10011100",3743 => "11000001",3744 => "01011001",3745 => "01011010",3746 => "01110111",3747 => "00010000",3748 => "11011101",3749 => "11001010",3750 => "11001000",3751 => "11110001",3752 => "10101010",3753 => "10110101",3754 => "10011101",3755 => "10101011",3756 => "11000010",3757 => "10000001",3758 => "11110010",3759 => "11110100",3760 => "11000001",3761 => "00111111",3762 => "10110111",3763 => "01000110",3764 => "00001101",3765 => "10101011",3766 => "01111010",3767 => "00010111",3768 => "11011011",3769 => "01011011",3770 => "01111000",3771 => "11100110",3772 => "10101010",3773 => "00001001",3774 => "00000111",3775 => "10111001",3776 => "11110000",3777 => "11011111",3778 => "01010100",3779 => "01111111",3780 => "11100010",3781 => "10100011",3782 => "01101000",3783 => "10011110",3784 => "11000011",3785 => "10011001",3786 => "00010111",3787 => "00000010",3788 => "11100011",3789 => "11100101",3790 => "10100100",3791 => "00010111",3792 => "10100110",3793 => "11111000",3794 => "11101001",3795 => "00010011",3796 => "01011010",3797 => "10010100",3798 => "01010000",3799 => "10110001",3800 => "01010010",3801 => "00100101",3802 => "11011101",3803 => "01111111",3804 => "10101011",3805 => "11001010",3806 => "10001100",3807 => "11110000",3808 => "01000100",3809 => "11100101",3810 => "11100010",3811 => "10010001",3812 => "10001010",3813 => "10111111",3814 => "00110100",3815 => "00111001",3816 => "01011000",3817 => "10010101",3818 => "11110001",3819 => "11100111",3820 => "10011010",3821 => "01100001",3822 => "10111000",3823 => "11111111",3824 => "00101110",3825 => "01001101",3826 => "01011111",3827 => "10000000",3828 => "10011010",3829 => "01101111",3830 => "00001011",3831 => "10111100",3832 => "10010110",3833 => "00100010",3834 => "11010010",3835 => "11010010",3836 => "11100001",3837 => "11111110",3838 => "10000000",3839 => "01110110",3840 => "00011100",3841 => "11000111",3842 => "10100001",3843 => "10010010",3844 => "01111001",3845 => "10100111",3846 => "01101101",3847 => "00011111",3848 => "01110100",3849 => "10111110",3850 => "00001101",3851 => "11000111",3852 => "00011111",3853 => "10111111",3854 => "11100101",3855 => "00110010",3856 => "11100001",3857 => "00001011",3858 => "00001101",3859 => "01010010",3860 => "01111100",3861 => "11111000",3862 => "01001111",3863 => "01010000",3864 => "11110011",3865 => "11111000",3866 => "01100101",3867 => "10001100",3868 => "00111011",3869 => "11100110",3870 => "01110010",3871 => "11110011",3872 => "10010110",3873 => "00100111",3874 => "00100111",3875 => "10111101",3876 => "10011101",3877 => "01111100",3878 => "01110110",3879 => "10110011",3880 => "00111001",3881 => "00011111",3882 => "10000001",3883 => "00110110",3884 => "00011101",3885 => "11110100",3886 => "10111101",3887 => "11111101",3888 => "01110111",3889 => "01000011",3890 => "01101100",3891 => "00010100",3892 => "10011010",3893 => "00011110",3894 => "00001010",3895 => "10101011",3896 => "01011000",3897 => "11100111",3898 => "01001000",3899 => "00101000",3900 => "01101111",3901 => "00001001",3902 => "01101000",3903 => "10111001",3904 => "11011101",3905 => "10010100",3906 => "10110010",3907 => "00010000",3908 => "10010100",3909 => "00011001",3910 => "11100001",3911 => "10110101",3912 => "11001110",3913 => "01011101",3914 => "10101111",3915 => "10001111",3916 => "11010001",3917 => "00011100",3918 => "00110010",3919 => "00101110",3920 => "00001011",3921 => "11110001",3922 => "11100111",3923 => "01101011",3924 => "01011010",3925 => "00000101",3926 => "10101001",3927 => "01111000",3928 => "01100000",3929 => "10101001",3930 => "01000111",3931 => "11001010",3932 => "00000000",3933 => "01001010",3934 => "01001001",3935 => "01100000",3936 => "10011011",3937 => "10010011",3938 => "10100110",3939 => "00111111",3940 => "01011000",3941 => "11111001",3942 => "11010111",3943 => "10110111",3944 => "00000010",3945 => "10110100",3946 => "01011100",3947 => "00010110",3948 => "10000101",3949 => "10101100",3950 => "10101001",3951 => "01001101",3952 => "11100110",3953 => "00001110",3954 => "00000110",3955 => "00010111",3956 => "00110001",3957 => "11101111",3958 => "00100011",3959 => "10010100",3960 => "00001111",3961 => "00011101",3962 => "11101101",3963 => "00011101",3964 => "11000101",3965 => "01001100",3966 => "11110100",3967 => "10101011",3968 => "10011011",3969 => "10000000",3970 => "10111111",3971 => "00111101",3972 => "11001010",3973 => "00001001",3974 => "11010101",3975 => "10111110",3976 => "11100001",3977 => "11101100",3978 => "01001110",3979 => "11010101",3980 => "10111111",3981 => "01100011",3982 => "01110110",3983 => "01110001",3984 => "00000010",3985 => "00101111",3986 => "11101001",3987 => "10000101",3988 => "00100101",3989 => "11111100",3990 => "01110100",3991 => "01111111",3992 => "00101000",3993 => "11001010",3994 => "11101010",3995 => "01110110",3996 => "10101001",3997 => "01100011",3998 => "01000110",3999 => "11100000",4000 => "11110110",4001 => "00110001",4002 => "01110110",4003 => "00000001",4004 => "11111011",4005 => "01001001",4006 => "01101100",4007 => "11101010",4008 => "01001101",4009 => "11101001",4010 => "00010010",4011 => "00011101",4012 => "01010000",4013 => "00111110",4014 => "00010011",4015 => "10001110",4016 => "11110100",4017 => "11010110",4018 => "00000101",4019 => "01010010",4020 => "10011010",4021 => "11001001",4022 => "00011011",4023 => "00010110",4024 => "11001110",4025 => "11101000",4026 => "01000001",4027 => "00100000",4028 => "01000110",4029 => "00101111",4030 => "10010101",4031 => "10001010",4032 => "11101010",4033 => "01111111",4034 => "01001011",4035 => "00111111",4036 => "00011010",4037 => "00101101",4038 => "00010100",4039 => "00110001",4040 => "00101111",4041 => "11001000",4042 => "01100010",4043 => "01010001",4044 => "11101111",4045 => "01111110",4046 => "11001100",4047 => "01100111",4048 => "00100101",4049 => "10010110",4050 => "10001101",4051 => "10001111",4052 => "01001001",4053 => "01010101",4054 => "00100001",4055 => "11100100",4056 => "11111010",4057 => "10010011",4058 => "11010100",4059 => "01100111",4060 => "01110010",4061 => "10111001",4062 => "11100001",4063 => "10101000",4064 => "00001000",4065 => "10011011",4066 => "01111101",4067 => "11100100",4068 => "10011111",4069 => "00011011",4070 => "11111111",4071 => "10101100",4072 => "11100010",4073 => "00011011",4074 => "10001101",4075 => "01100101",4076 => "11111010",4077 => "11111001",4078 => "11011100",4079 => "01100010",4080 => "00000011",4081 => "01011100",4082 => "00101101",4083 => "00001100",4084 => "01100011",4085 => "11100101",4086 => "01010110",4087 => "01010110",4088 => "00110010",4089 => "00001101",4090 => "10010001",4091 => "01010001",4092 => "00111110",4093 => "11100101",4094 => "11010011",4095 => "11111011",4096 => "00100000",4097 => "10001000",4098 => "11010000",4099 => "10000101",4100 => "00001000",4101 => "00110010",4102 => "00101110",4103 => "10000111",4104 => "01001010",4105 => "00101011",4106 => "00111100",4107 => "10101101",4108 => "10011000",4109 => "10000000",4110 => "00101010",4111 => "10101011",4112 => "00010001",4113 => "11111001",4114 => "00011100",4115 => "00101000",4116 => "00101001",4117 => "01101101",4118 => "00111111",4119 => "01100111",4120 => "11100111",4121 => "00110110",4122 => "10100010",4123 => "00001101",4124 => "01010111",4125 => "10010001",4126 => "00101000",4127 => "11101110",4128 => "11100110",4129 => "10001011",4130 => "01011101",4131 => "01011001",4132 => "01010101",4133 => "01011100",4134 => "11010001",4135 => "10001011",4136 => "11000111",4137 => "10111111",4138 => "10100101",4139 => "10011010",4140 => "01101000",4141 => "10001001",4142 => "10001010",4143 => "11000100",4144 => "11110111",4145 => "10011111",4146 => "10110100",4147 => "00100001",4148 => "00011111",4149 => "01111100",4150 => "10001011",4151 => "01110010",4152 => "01101110",4153 => "01100111",4154 => "00000011",4155 => "00100010",4156 => "10110100",4157 => "00101010",4158 => "00011000",4159 => "11110100",4160 => "00110011",4161 => "10110011",4162 => "10100000",4163 => "01111000",4164 => "11110101",4165 => "10001010",4166 => "00100011",4167 => "11110111",4168 => "01100000",4169 => "11100101",4170 => "10100001",4171 => "00011001",4172 => "11000111",4173 => "01100100",4174 => "00000111",4175 => "01101101",4176 => "10101011",4177 => "01110111",4178 => "10010001",4179 => "11000100",4180 => "01000010",4181 => "00101101",4182 => "01011101",4183 => "01010011",4184 => "11000010",4185 => "11100010",4186 => "11001001",4187 => "10010010",4188 => "01011100",4189 => "01101101",4190 => "10001111",4191 => "01001000",4192 => "11100000",4193 => "10110011",4194 => "01101100",4195 => "10010110",4196 => "11100101",4197 => "11011001",4198 => "00110001",4199 => "00101110",4200 => "01011010",4201 => "10001110",4202 => "11100110",4203 => "00100101",4204 => "11100111",4205 => "10011110",4206 => "11011001",4207 => "10100000",4208 => "01100101",4209 => "00100001",4210 => "00110000",4211 => "10111000",4212 => "10001110",4213 => "01010000",4214 => "11110001",4215 => "11111010",4216 => "00101111",4217 => "00001100",4218 => "11100000",4219 => "00111100",4220 => "10111110",4221 => "00000010",4222 => "10111001",4223 => "11011011",4224 => "01110110",4225 => "00110100",4226 => "00000011",4227 => "00111001",4228 => "01111000",4229 => "00011000",4230 => "10000011",4231 => "10100101",4232 => "11010110",4233 => "11101001",4234 => "10010110",4235 => "11001110",4236 => "00101001",4237 => "10110000",4238 => "00010100",4239 => "01100000",4240 => "00011110",4241 => "01100001",4242 => "01100101",4243 => "10100011",4244 => "11100101",4245 => "11100001",4246 => "01011000",4247 => "01111011",4248 => "00111110",4249 => "00101100",4250 => "11000111",4251 => "00001100",4252 => "11011011",4253 => "10011000",4254 => "11010000",4255 => "10001101",4256 => "01110110",4257 => "11100010",4258 => "00010000",4259 => "10100111",4260 => "11101100",4261 => "10000001",4262 => "01111001",4263 => "01111000",4264 => "10101000",4265 => "00000011",4266 => "10110001",4267 => "11110000",4268 => "10101001",4269 => "10110000",4270 => "10000110",4271 => "01101100",4272 => "10000111",4273 => "11011110",4274 => "10000101",4275 => "01011000",4276 => "01000100",4277 => "10101101",4278 => "01000011",4279 => "10110101",4280 => "11110100",4281 => "01010011",4282 => "11000011",4283 => "00101100",4284 => "11000000",4285 => "10110000",4286 => "11010011",4287 => "01111101",4288 => "11000011",4289 => "10101011",4290 => "00010010",4291 => "10011100",4292 => "00111011",4293 => "01011010",4294 => "00011001",4295 => "10111111",4296 => "10011011",4297 => "10011101",4298 => "11000011",4299 => "11011001",4300 => "00101111",4301 => "01100000",4302 => "11100100",4303 => "01001010",4304 => "10001111",4305 => "01110110",4306 => "11101100",4307 => "11101001",4308 => "11101001",4309 => "10011101",4310 => "10100100",4311 => "00110011",4312 => "10111000",4313 => "00100100",4314 => "01111010",4315 => "00001001",4316 => "01011101",4317 => "00010111",4318 => "10111100",4319 => "00011111",4320 => "00111010",4321 => "00100010",4322 => "10001000",4323 => "10111001",4324 => "01001001",4325 => "10101100",4326 => "11111000",4327 => "01111100",4328 => "00110000",4329 => "00000100",4330 => "01010111",4331 => "00001001",4332 => "01011110",4333 => "01001010",4334 => "01000000",4335 => "10101111",4336 => "00110000",4337 => "10001111",4338 => "01010010",4339 => "11000100",4340 => "00000011",4341 => "11000011",4342 => "10000010",4343 => "00101100",4344 => "00000110",4345 => "00111001",4346 => "10010111",4347 => "00011011",4348 => "11010000",4349 => "01011111",4350 => "10000110",4351 => "01110111",4352 => "01101110",4353 => "01001111",4354 => "00111000",4355 => "11100110",4356 => "11110000",4357 => "01010100",4358 => "00100000",4359 => "10011100",4360 => "11010011",4361 => "10001000",4362 => "11011010",4363 => "00101001",4364 => "00011101",4365 => "10011110",4366 => "10111010",4367 => "11101011",4368 => "01101011",4369 => "11010010",4370 => "11010000",4371 => "01011111",4372 => "00001000",4373 => "00011100",4374 => "01011000",4375 => "10010111",4376 => "11010010",4377 => "11010111",4378 => "01011110",4379 => "11111111",4380 => "01100001",4381 => "11100000",4382 => "00010001",4383 => "01100101",4384 => "11110100",4385 => "10011000",4386 => "00010110",4387 => "10111000",4388 => "10101011",4389 => "10001011",4390 => "11011110",4391 => "01110110",4392 => "11000011",4393 => "01110111",4394 => "10010110",4395 => "01100111",4396 => "10101000",4397 => "01010110",4398 => "11011010",4399 => "11101111",4400 => "01001110",4401 => "10101110",4402 => "11111010",4403 => "10000011",4404 => "01000101",4405 => "00101100",4406 => "10000100",4407 => "01111101",4408 => "01001010",4409 => "00100111",4410 => "01110110",4411 => "01100110",4412 => "00000010",4413 => "11100101",4414 => "10010010",4415 => "01100000",4416 => "11101000",4417 => "00010111",4418 => "01111000",4419 => "10010101",4420 => "11001100",4421 => "01101000",4422 => "11111100",4423 => "10000011",4424 => "11011011",4425 => "10010110",4426 => "11000101",4427 => "11101110",4428 => "10101100",4429 => "11010100",4430 => "00001101",4431 => "11101110",4432 => "11101100",4433 => "11011010",4434 => "01101011",4435 => "01011101",4436 => "11110101",4437 => "10111010",4438 => "10010011",4439 => "10000101",4440 => "10101101",4441 => "11101111",4442 => "01101001",4443 => "10010111",4444 => "01000100",4445 => "10000011",4446 => "10011101",4447 => "01110111",4448 => "10001110",4449 => "10000110",4450 => "01100010",4451 => "10001000",4452 => "00000101",4453 => "11111010",4454 => "11101000",4455 => "11011001",4456 => "00011101",4457 => "00010011",4458 => "11100111",4459 => "11110111",4460 => "11011100",4461 => "01011101",4462 => "11110101",4463 => "00110011",4464 => "01100111",4465 => "01001000",4466 => "11111010",4467 => "00100110",4468 => "01000100",4469 => "01011110",4470 => "11100100",4471 => "01010101",4472 => "01111000",4473 => "10010101",4474 => "01001111",4475 => "00010010",4476 => "01000110",4477 => "10100111",4478 => "00100100",4479 => "11001100",4480 => "01101111",4481 => "10001101",4482 => "00110110",4483 => "10000111",4484 => "00011010",4485 => "00100001",4486 => "10101110",4487 => "00100000",4488 => "00101101",4489 => "10011101",4490 => "00001110",4491 => "00000001",4492 => "10110101",4493 => "00001101",4494 => "10011100",4495 => "01011101",4496 => "01100111",4497 => "00010010",4498 => "10011001",4499 => "00110101",4500 => "11001010",4501 => "00111100",4502 => "01001001",4503 => "01000111",4504 => "01110100",4505 => "10000010",4506 => "01100110",4507 => "01000111",4508 => "00101110",4509 => "00110010",4510 => "11000100",4511 => "00110011",4512 => "10111101",4513 => "01110100",4514 => "00101111",4515 => "10001100",4516 => "00101001",4517 => "01111100",4518 => "00101101",4519 => "00010000",4520 => "10000110",4521 => "10000001",4522 => "01111111",4523 => "01010000",4524 => "11001110",4525 => "00001100",4526 => "11000110",4527 => "00011111",4528 => "00001100",4529 => "01111101",4530 => "10000110",4531 => "11111101",4532 => "00110101",4533 => "10011101",4534 => "10101000",4535 => "00001111",4536 => "11010101",4537 => "10111011",4538 => "01010110",4539 => "01101101",4540 => "01011100",4541 => "00101101",4542 => "11111111",4543 => "11011011",4544 => "11101001",4545 => "10110011",4546 => "01011101",4547 => "10010001",4548 => "00110011",4549 => "11011000",4550 => "01011001",4551 => "00101111",4552 => "10001110",4553 => "11110011",4554 => "11011110",4555 => "01101011",4556 => "00110010",4557 => "00011110",4558 => "10001001",4559 => "11011011",4560 => "00010000",4561 => "01101111",4562 => "01111011",4563 => "10101101",4564 => "11010100",4565 => "11011110",4566 => "11111110",4567 => "11001111",4568 => "01100111",4569 => "01111100",4570 => "11001101",4571 => "01111101",4572 => "01100000",4573 => "10011111",4574 => "00000000",4575 => "00110111",4576 => "11111010",4577 => "10000001",4578 => "01001001",4579 => "11010000",4580 => "11111000",4581 => "00011111",4582 => "00010010",4583 => "01100001",4584 => "10111011",4585 => "10010010",4586 => "00001111",4587 => "10001001",4588 => "00101000",4589 => "01100111",4590 => "01010001",4591 => "00110011",4592 => "11111000",4593 => "11000001",4594 => "10100011",4595 => "10011001",4596 => "01101101",4597 => "00110000",4598 => "00101111",4599 => "10000111",4600 => "10001111",4601 => "11000100",4602 => "01001010",4603 => "11100100",4604 => "10110111",4605 => "00101110",4606 => "00011011",4607 => "01011110",4608 => "10000101",4609 => "00001010",4610 => "10100001",4611 => "11010101",4612 => "01011001",4613 => "10011000",4614 => "00001111",4615 => "10001011",4616 => "01000100",4617 => "00011101",4618 => "11101101",4619 => "01100101",4620 => "11010111",4621 => "11101101",4622 => "00001110",4623 => "10001010",4624 => "11111110",4625 => "00000111",4626 => "01011100",4627 => "01011110",4628 => "10000110",4629 => "01000010",4630 => "10010110",4631 => "11001101",4632 => "00010111",4633 => "00011100",4634 => "10100100",4635 => "11100110",4636 => "00100110",4637 => "10001010",4638 => "01001011",4639 => "01000001",4640 => "11110001",4641 => "10000110",4642 => "00000000",4643 => "11110111",4644 => "00000100",4645 => "01110010",4646 => "00011110",4647 => "11111101",4648 => "11100011",4649 => "11101100",4650 => "01011010",4651 => "11010111",4652 => "00001100",4653 => "11111100",4654 => "11010100",4655 => "11101111",4656 => "00010000",4657 => "10101011",4658 => "10110110",4659 => "00011100",4660 => "01111011",4661 => "10010111",4662 => "01111111",4663 => "01101001",4664 => "11100110",4665 => "00001100",4666 => "10000110",4667 => "01000000",4668 => "11111011",4669 => "10101110",4670 => "11001001",4671 => "00101100",4672 => "01011110",4673 => "10111110",4674 => "00101111",4675 => "01000001",4676 => "11101010",4677 => "01001011",4678 => "01100100",4679 => "01101011",4680 => "10001000",4681 => "10011011",4682 => "11100010",4683 => "00111110",4684 => "11101111",4685 => "01000100",4686 => "01000010",4687 => "11101100",4688 => "00000010",4689 => "10110001",4690 => "01000111",4691 => "01011110",4692 => "10001111",4693 => "11001110",4694 => "11110011",4695 => "00101010",4696 => "11000011",4697 => "10010111",4698 => "00001001",4699 => "00011011",4700 => "01011000",4701 => "10011011",4702 => "00100111",4703 => "00101001",4704 => "00000101",4705 => "01000000",4706 => "11000001",4707 => "00101010",4708 => "10110111",4709 => "00111010",4710 => "01001111",4711 => "01001010",4712 => "11111000",4713 => "10000000",4714 => "01101111",4715 => "11010010",4716 => "00000110",4717 => "10101011",4718 => "01011110",4719 => "11010011",4720 => "00000110",4721 => "00101101",4722 => "01100010",4723 => "10001110",4724 => "00100111",4725 => "01001001",4726 => "01101100",4727 => "10011011",4728 => "11000111",4729 => "10110010",4730 => "00110000",4731 => "01111010",4732 => "01100110",4733 => "00010101",4734 => "00000110",4735 => "10101010",4736 => "00010010",4737 => "01110110",4738 => "11100001",4739 => "01001101",4740 => "00111011",4741 => "10101101",4742 => "01110011",4743 => "00111111",4744 => "00110110",4745 => "10101010",4746 => "10111110",4747 => "01000101",4748 => "00010110",4749 => "10011101",4750 => "00111001",4751 => "10111011",4752 => "00110001",4753 => "10101010",4754 => "11010000",4755 => "10100111",4756 => "01101111",4757 => "10001110",4758 => "10100000",4759 => "00011101",4760 => "11011100",4761 => "00000111",4762 => "10011011",4763 => "01000000",4764 => "01100001",4765 => "00110011",4766 => "01011100",4767 => "01010100",4768 => "01011000",4769 => "01100110",4770 => "00110110",4771 => "00111001",4772 => "01111001",4773 => "00101000",4774 => "10001011",4775 => "10111000",4776 => "00101111",4777 => "10100000",4778 => "11010001",4779 => "11101110",4780 => "10101010",4781 => "01111100",4782 => "00001111",4783 => "11010000",4784 => "11011010",4785 => "11001111",4786 => "00000111",4787 => "00001000",4788 => "11011101",4789 => "10000011",4790 => "00000011",4791 => "00100000",4792 => "11101010",4793 => "11011011",4794 => "10110100",4795 => "01111011",4796 => "10111010",4797 => "10111001",4798 => "00100011",4799 => "11000001",4800 => "10101000",4801 => "00111100",4802 => "01110000",4803 => "01001001",4804 => "00011001",4805 => "11111001",4806 => "01001001",4807 => "01010100",4808 => "00101101",4809 => "10111100",4810 => "00001101",4811 => "10010100",4812 => "00111101",4813 => "00000100",4814 => "11000100",4815 => "00100111",4816 => "01111001",4817 => "01101100",4818 => "11110100",4819 => "01101011",4820 => "01000110",4821 => "11010001",4822 => "01010101",4823 => "11011100",4824 => "01010110",4825 => "00111000",4826 => "11110010",4827 => "01100101",4828 => "11100101",4829 => "10000011",4830 => "11111000",4831 => "11101100",4832 => "10100110",4833 => "10010100",4834 => "01001101",4835 => "01111011",4836 => "11001010",4837 => "11101110",4838 => "00010110",4839 => "01010110",4840 => "11101010",4841 => "11100100",4842 => "11111011",4843 => "11111100",4844 => "00101000",4845 => "00011000",4846 => "10111110",4847 => "10100110",4848 => "10000010",4849 => "00011011",4850 => "11111110",4851 => "00100000",4852 => "01000000",4853 => "00111000",4854 => "10100101",4855 => "00010010",4856 => "00100110",4857 => "00101100",4858 => "01000101",4859 => "00000010",4860 => "10111001",4861 => "11010101",4862 => "11001000",4863 => "10010101",4864 => "10111110",4865 => "11101001",4866 => "11011100",4867 => "00010110",4868 => "00000101",4869 => "10101000",4870 => "11110101",4871 => "11010011",4872 => "10010101",4873 => "10111000",4874 => "00110010",4875 => "00100011",4876 => "11111011",4877 => "10001110",4878 => "10101111",4879 => "01110101",4880 => "01011111",4881 => "10001011",4882 => "10101101",4883 => "10110111",4884 => "11110000",4885 => "00100111",4886 => "01000001",4887 => "00001000",4888 => "00001110",4889 => "00101111",4890 => "10101000",4891 => "00010011",4892 => "00000001",4893 => "10010001",4894 => "01011101",4895 => "00101000",4896 => "10111110",4897 => "01111100",4898 => "10011100",4899 => "00111110",4900 => "00000011",4901 => "00111101",4902 => "11001100",4903 => "10001001",4904 => "00110010",4905 => "11111010",4906 => "00110001",4907 => "00010010",4908 => "11011101",4909 => "01010000",4910 => "00100100",4911 => "01100100",4912 => "10100011",4913 => "00100000",4914 => "10000001",4915 => "00001010",4916 => "10101100",4917 => "11001001",4918 => "01001010",4919 => "11000001",4920 => "00101100",4921 => "10100010",4922 => "01101001",4923 => "10000111",4924 => "01010111",4925 => "00100100",4926 => "10101111",4927 => "00100000",4928 => "11011111",4929 => "00000100",4930 => "10101111",4931 => "10110000",4932 => "00101111",4933 => "11010100",4934 => "01100101",4935 => "11000001",4936 => "11101001",4937 => "00011101",4938 => "10100101",4939 => "11001111",4940 => "01100111",4941 => "10001011",4942 => "11110111",4943 => "10110101",4944 => "01101001",4945 => "01011101",4946 => "01001011",4947 => "01110111",4948 => "00001011",4949 => "00001011",4950 => "00010111",4951 => "10010100",4952 => "00110011",4953 => "10010010",4954 => "00111111",4955 => "10101001",4956 => "10010110",4957 => "11010101",4958 => "01001101",4959 => "01101111",4960 => "01000000",4961 => "00101001",4962 => "00100110",4963 => "11101111",4964 => "00001111",4965 => "00010000",4966 => "10101100",4967 => "00010111",4968 => "01011110",4969 => "01111010",4970 => "10001000",4971 => "01001000",4972 => "10000000",4973 => "00011011",4974 => "00101110",4975 => "11001011",4976 => "00110000",4977 => "00010010",4978 => "10010111",4979 => "01110101",4980 => "00100001",4981 => "00001110",4982 => "11100100",4983 => "10011010",4984 => "00001001",4985 => "10101011",4986 => "01011001",4987 => "11000100",4988 => "00111100",4989 => "10000100",4990 => "01110001",4991 => "11010001",4992 => "11000001",4993 => "10101100",4994 => "00010111",4995 => "01001000",4996 => "01110000",4997 => "10011110",4998 => "10001111",4999 => "10110010",5000 => "10000000",5001 => "10111001",5002 => "00101011",5003 => "01110000",5004 => "10000100",5005 => "11011110",5006 => "10101000",5007 => "01100011",5008 => "10101101",5009 => "11101111",5010 => "10100001",5011 => "10110101",5012 => "00111000",5013 => "11010100",5014 => "11100011",5015 => "00101010",5016 => "00100100",5017 => "01000101",5018 => "01011101",5019 => "11100011",5020 => "00000001",5021 => "10000000",5022 => "11111000",5023 => "00100110",5024 => "10110100",5025 => "01110010",5026 => "11011110",5027 => "00010011",5028 => "00110100",5029 => "11100111",5030 => "11101110",5031 => "10011110",5032 => "10001110",5033 => "11010001",5034 => "11000011",5035 => "10001110",5036 => "10000110",5037 => "10110010",5038 => "11110011",5039 => "00010011",5040 => "00010101",5041 => "00001110",5042 => "11111001",5043 => "00101000",5044 => "10000011",5045 => "11111101",5046 => "10001011",5047 => "00011101",5048 => "11101100",5049 => "01100111",5050 => "01100001",5051 => "00101100",5052 => "00011010",5053 => "00000011",5054 => "11011001",5055 => "10000001",5056 => "00010101",5057 => "10011110",5058 => "10100101",5059 => "00011101",5060 => "01011000",5061 => "00010110",5062 => "11011101",5063 => "11110101",5064 => "11000101",5065 => "11100101",5066 => "10111111",5067 => "00011110",5068 => "00010001",5069 => "11010010",5070 => "10110010",5071 => "11010101",5072 => "01010001",5073 => "11010010",5074 => "11000000",5075 => "00010001",5076 => "11111101",5077 => "11111011",5078 => "00101011",5079 => "10011001",5080 => "01101111",5081 => "11010100",5082 => "11101000",5083 => "11010110",5084 => "10001000",5085 => "11110100",5086 => "11011111",5087 => "10011110",5088 => "11111111",5089 => "11011111",5090 => "00110111",5091 => "11001011",5092 => "10100000",5093 => "11101101",5094 => "10011010",5095 => "00100111",5096 => "10010000",5097 => "11011101",5098 => "01100110",5099 => "01110100",5100 => "11101111",5101 => "11100001",5102 => "10101011",5103 => "00011111",5104 => "00010110",5105 => "11011010",5106 => "11110110",5107 => "10011010",5108 => "11110001",5109 => "01010010",5110 => "11000010",5111 => "10101111",5112 => "11111011",5113 => "01111110",5114 => "00001111",5115 => "00010111",5116 => "10101110",5117 => "11001100",5118 => "01001100",5119 => "11010011",5120 => "01000001",5121 => "00011000",5122 => "10110111",5123 => "10011010",5124 => "01011000",5125 => "10101110",5126 => "00000110",5127 => "11010001",5128 => "01011011",5129 => "10111100",5130 => "11100011",5131 => "11001100",5132 => "11101010",5133 => "11010011",5134 => "10111111",5135 => "11010000",5136 => "01011100",5137 => "00100101",5138 => "01001010",5139 => "11010010",5140 => "11100101",5141 => "01001110",5142 => "01100100",5143 => "10000101",5144 => "01111100",5145 => "00001110",5146 => "11110110",5147 => "10101100",5148 => "00011110",5149 => "00101011",5150 => "01001011",5151 => "10110011",5152 => "10101001",5153 => "11000100",5154 => "10111111",5155 => "11000100",5156 => "10110100",5157 => "11000010",5158 => "00001101",5159 => "00110010",5160 => "11100101",5161 => "11011111",5162 => "10011000",5163 => "00111000",5164 => "10011100",5165 => "10010000",5166 => "11100000",5167 => "00011110",5168 => "11101010",5169 => "01010111",5170 => "01010101",5171 => "00100110",5172 => "01101001",5173 => "00011110",5174 => "01000111",5175 => "00110010",5176 => "00101101",5177 => "00100111",5178 => "11101000",5179 => "11100110",5180 => "10110011",5181 => "01111101",5182 => "10001010",5183 => "10010010",5184 => "01111010",5185 => "10011000",5186 => "00100011",5187 => "11001000",5188 => "00100001",5189 => "00000110",5190 => "10000100",5191 => "01101001",5192 => "10001011",5193 => "01000110",5194 => "10001000",5195 => "10000011",5196 => "11110111",5197 => "11100110",5198 => "00110101",5199 => "10010101",5200 => "00011011",5201 => "11111111",5202 => "01001100",5203 => "10101110",5204 => "01001110",5205 => "11000010",5206 => "01101011",5207 => "11011110",5208 => "00011010",5209 => "01011011",5210 => "00101011",5211 => "00001100",5212 => "10111101",5213 => "11111000",5214 => "10001011",5215 => "10111101",5216 => "01100101",5217 => "01001010",5218 => "00100100",5219 => "00010100",5220 => "00010101",5221 => "11100001",5222 => "10000010",5223 => "10011111",5224 => "10111010",5225 => "00111000",5226 => "11011111",5227 => "01110000",5228 => "00000111",5229 => "00001011",5230 => "01101101",5231 => "01111000",5232 => "10000111",5233 => "11000011",5234 => "10001110",5235 => "01000011",5236 => "11110011",5237 => "01100010",5238 => "10101110",5239 => "01101100",5240 => "01110010",5241 => "01101101",5242 => "00011101",5243 => "01000001",5244 => "10100001",5245 => "01001000",5246 => "11111111",5247 => "01010101",5248 => "10101001",5249 => "10101100",5250 => "11001001",5251 => "01100100",5252 => "11000101",5253 => "11011110",5254 => "11100011",5255 => "00010010",5256 => "10111110",5257 => "01011111",5258 => "01000001",5259 => "11010101",5260 => "00111011",5261 => "00010010",5262 => "11101100",5263 => "11001100",5264 => "00000101",5265 => "01011100",5266 => "10100100",5267 => "10000011",5268 => "01111010",5269 => "10001111",5270 => "00010010",5271 => "00011101",5272 => "01111001",5273 => "10111010",5274 => "11101101",5275 => "11101111",5276 => "10111100",5277 => "11011001",5278 => "01100100",5279 => "00111100",5280 => "11101000",5281 => "10000011",5282 => "10110101",5283 => "11111101",5284 => "01111100",5285 => "01001000",5286 => "10111010",5287 => "11100000",5288 => "00001000",5289 => "01010010",5290 => "11010111",5291 => "01000000",5292 => "10011111",5293 => "00110010",5294 => "01001101",5295 => "11110010",5296 => "01001010",5297 => "01000000",5298 => "10010111",5299 => "11111010",5300 => "10011011",5301 => "00001100",5302 => "11111111",5303 => "01000010",5304 => "10101100",5305 => "00000101",5306 => "00110110",5307 => "01000000",5308 => "11111100",5309 => "10110100",5310 => "01111010",5311 => "01101110",5312 => "10110111",5313 => "00100011",5314 => "11111101",5315 => "01000111",5316 => "11010101",5317 => "00101110",5318 => "10110101",5319 => "10101001",5320 => "01001111",5321 => "11111101",5322 => "01100000",5323 => "11100010",5324 => "00001001",5325 => "10100100",5326 => "00101010",5327 => "11010011",5328 => "00110101",5329 => "01000110",5330 => "01001010",5331 => "10000100",5332 => "00011110",5333 => "10010110",5334 => "11011001",5335 => "10101000",5336 => "11100111",5337 => "00011111",5338 => "10100011",5339 => "01100010",5340 => "00100100",5341 => "01011000",5342 => "00100011",5343 => "10000000",5344 => "01011110",5345 => "10011101",5346 => "10100000",5347 => "11000000",5348 => "11101111",5349 => "10101110",5350 => "01101101",5351 => "10000111",5352 => "01011000",5353 => "11000110",5354 => "00110100",5355 => "00000101",5356 => "10000010",5357 => "01010111",5358 => "01001111",5359 => "00011110",5360 => "00000100",5361 => "10101010",5362 => "11010101",5363 => "10110001",5364 => "01111101",5365 => "01010111",5366 => "11101111",5367 => "11101010",5368 => "11111111",5369 => "10111010",5370 => "01110111",5371 => "10010011",5372 => "00111000",5373 => "01000100",5374 => "10011011",5375 => "01011100",5376 => "11011110",5377 => "11001010",5378 => "11100111",5379 => "01111000",5380 => "01111010",5381 => "10000110",5382 => "01110111",5383 => "10011011",5384 => "00000001",5385 => "11011011",5386 => "00001001",5387 => "01010001",5388 => "01110011",5389 => "00000010",5390 => "11000011",5391 => "00001110",5392 => "10101011",5393 => "10001110",5394 => "01111110",5395 => "10111101",5396 => "11110111",5397 => "10100010",5398 => "00111111",5399 => "01111010",5400 => "00011100",5401 => "01011100",5402 => "00101000",5403 => "11011110",5404 => "01001110",5405 => "01010101",5406 => "00000000",5407 => "10111000",5408 => "11110000",5409 => "00011001",5410 => "10000000",5411 => "01101101",5412 => "11001111",5413 => "10000011",5414 => "01011011",5415 => "00010111",5416 => "00110110",5417 => "00001011",5418 => "11111100",5419 => "01000110",5420 => "10101010",5421 => "10011001",5422 => "10111101",5423 => "11010010",5424 => "10111111",5425 => "10101001",5426 => "01011010",5427 => "11000001",5428 => "01101011",5429 => "01101111",5430 => "11010001",5431 => "00010010",5432 => "11110011",5433 => "11110110",5434 => "00100001",5435 => "00100010",5436 => "10101101",5437 => "11001011",5438 => "00111110",5439 => "10000010",5440 => "10000101",5441 => "11010000",5442 => "00010101",5443 => "00001000",5444 => "00011000",5445 => "10100110",5446 => "11000010",5447 => "10010001",5448 => "00011001",5449 => "01110000",5450 => "11011000",5451 => "01111001",5452 => "11000001",5453 => "11101111",5454 => "01001001",5455 => "01111000",5456 => "10111001",5457 => "11000101",5458 => "11001001",5459 => "10000110",5460 => "00100101",5461 => "01010111",5462 => "10101010",5463 => "01111100",5464 => "01010000",5465 => "01001100",5466 => "11000100",5467 => "01111110",5468 => "11011101",5469 => "01110101",5470 => "00110011",5471 => "00011000",5472 => "10100000",5473 => "01100011",5474 => "11000001",5475 => "00110000",5476 => "01011111",5477 => "11011100",5478 => "10101110",5479 => "11010011",5480 => "11101101",5481 => "11110110",5482 => "00011001",5483 => "11000010",5484 => "01011110",5485 => "00010101",5486 => "11110100",5487 => "00001100",5488 => "01001111",5489 => "11110000",5490 => "00011100",5491 => "11101011",5492 => "01111001",5493 => "11011101",5494 => "11001111",5495 => "10011010",5496 => "01010001",5497 => "01110101",5498 => "11011010",5499 => "11111111",5500 => "11101110",5501 => "01011001",5502 => "01100011",5503 => "01111100",5504 => "11000001",5505 => "01111011",5506 => "01010011",5507 => "11101100",5508 => "00101100",5509 => "10010010",5510 => "10100110",5511 => "01011010",5512 => "00111100",5513 => "11000000",5514 => "10110000",5515 => "11001011",5516 => "11011110",5517 => "10111011",5518 => "00010000",5519 => "00000001",5520 => "01001010",5521 => "11010001",5522 => "00100000",5523 => "10010101",5524 => "11111010",5525 => "10011011",5526 => "10101000",5527 => "10111100",5528 => "11100010",5529 => "00111011",5530 => "01000110",5531 => "00010101",5532 => "11001010",5533 => "10011100",5534 => "11110010",5535 => "10010010",5536 => "00011101",5537 => "11010000",5538 => "01001000",5539 => "01110110",5540 => "11011101",5541 => "00100001",5542 => "10000010",5543 => "11010111",5544 => "00011000",5545 => "10101001",5546 => "01101101",5547 => "01000100",5548 => "11010101",5549 => "11010001",5550 => "11110001",5551 => "01100111",5552 => "10110010",5553 => "00110000",5554 => "10110110",5555 => "00101000",5556 => "00000101",5557 => "00100110",5558 => "10100111",5559 => "11111100",5560 => "00001010",5561 => "00110001",5562 => "10111110",5563 => "00000111",5564 => "11111100",5565 => "11100011",5566 => "11111111",5567 => "01110100",5568 => "10010011",5569 => "10000110",5570 => "11001000",5571 => "10101010",5572 => "11000111",5573 => "01010000",5574 => "01011111",5575 => "11000100",5576 => "11001111",5577 => "00010101",5578 => "11111111",5579 => "11111010",5580 => "11010101",5581 => "00011011",5582 => "00010000",5583 => "11011010",5584 => "00000000",5585 => "00011110",5586 => "00011010",5587 => "00101001",5588 => "00110001",5589 => "00000000",5590 => "00100111",5591 => "01111010",5592 => "00011111",5593 => "01100111",5594 => "11101110",5595 => "10001110",5596 => "01111100",5597 => "10000110",5598 => "11100000",5599 => "11100000",5600 => "11001111",5601 => "00111000",5602 => "11111100",5603 => "11110110",5604 => "01100100",5605 => "10010111",5606 => "00000000",5607 => "10010110",5608 => "11110111",5609 => "10111010",5610 => "00111100",5611 => "01100110",5612 => "11110101",5613 => "10011010",5614 => "01000101",5615 => "10111010",5616 => "11011111",5617 => "00010000",5618 => "11100011",5619 => "10010110",5620 => "01111011",5621 => "01101100",5622 => "01010011",5623 => "00111100",5624 => "01100100",5625 => "10011110",5626 => "11011011",5627 => "10100000",5628 => "11001000",5629 => "10001010",5630 => "11110001",5631 => "11001001",5632 => "11110011",5633 => "10001101",5634 => "10000011",5635 => "11000110",5636 => "00111001",5637 => "00110010",5638 => "11001011",5639 => "11111101",5640 => "10111001",5641 => "00000000",5642 => "11011101",5643 => "10010100",5644 => "10101110",5645 => "11001001",5646 => "01110100",5647 => "00000010",5648 => "10001001",5649 => "10001101",5650 => "01001001",5651 => "10101111",5652 => "10011011",5653 => "01010001",5654 => "01010111",5655 => "01001101",5656 => "00110101",5657 => "01010001",5658 => "01010111",5659 => "00100010",5660 => "11010110",5661 => "00001111",5662 => "01010001",5663 => "11001010",5664 => "00101100",5665 => "10001010",5666 => "00000110",5667 => "10111110",5668 => "00101001",5669 => "01110100",5670 => "10011001",5671 => "00010010",5672 => "01010100",5673 => "01110111",5674 => "10111111",5675 => "01000111",5676 => "00100110",5677 => "01001001",5678 => "11110000",5679 => "01010100",5680 => "00001100",5681 => "11010000",5682 => "01011011",5683 => "11100100",5684 => "10010000",5685 => "10111110",5686 => "10110101",5687 => "00101101",5688 => "11001001",5689 => "10000100",5690 => "01001110",5691 => "11001001",5692 => "11100111",5693 => "10100011",5694 => "01001110",5695 => "10011110",5696 => "10110001",5697 => "11100001",5698 => "01010100",5699 => "11111100",5700 => "00110011",5701 => "01101111",5702 => "10111110",5703 => "01101000",5704 => "01010001",5705 => "00011000",5706 => "00011010",5707 => "10100000",5708 => "11101111",5709 => "10101011",5710 => "10100010",5711 => "11011111",5712 => "11010111",5713 => "11011100",5714 => "11011010",5715 => "10101101",5716 => "11110000",5717 => "01001011",5718 => "10000101",5719 => "11011110",5720 => "11111110",5721 => "00111000",5722 => "00111111",5723 => "01101011",5724 => "00000001",5725 => "01010000",5726 => "11101011",5727 => "01000011",5728 => "10001101",5729 => "00100011",5730 => "00101010",5731 => "00111001",5732 => "10110110",5733 => "01110110",5734 => "00110111",5735 => "01011111",5736 => "11000000",5737 => "00011000",5738 => "11101101",5739 => "11101101",5740 => "11010100",5741 => "01001111",5742 => "01101011",5743 => "01110111",5744 => "01101110",5745 => "00111100",5746 => "11100010",5747 => "00100100",5748 => "01011100",5749 => "00110101",5750 => "10001010",5751 => "11001101",5752 => "00110010",5753 => "01011000",5754 => "11111110",5755 => "01100000",5756 => "01001111",5757 => "11000001",5758 => "10111101",5759 => "10010011",5760 => "11100111",5761 => "00110111",5762 => "10100101",5763 => "00010111",5764 => "11100111",5765 => "10010111",5766 => "01000111",5767 => "10010101",5768 => "00101000",5769 => "11110000",5770 => "00111001",5771 => "00001111",5772 => "01110001",5773 => "00101111",5774 => "01010111",5775 => "11010011",5776 => "10000011",5777 => "01000110",5778 => "11001110",5779 => "00011110",5780 => "00111100",5781 => "10011100",5782 => "11101101",5783 => "10110010",5784 => "10001100",5785 => "11100100",5786 => "11100100",5787 => "10100010",5788 => "00110000",5789 => "11100111",5790 => "11011110",5791 => "11010111",5792 => "00011001",5793 => "01000110",5794 => "01010110",5795 => "00111111",5796 => "00011010",5797 => "10000101",5798 => "00111011",5799 => "10001000",5800 => "01101110",5801 => "11010110",5802 => "00010101",5803 => "00001000",5804 => "11000111",5805 => "10001100",5806 => "10000111",5807 => "10110100",5808 => "01101110",5809 => "10011000",5810 => "00111000",5811 => "00000110",5812 => "10100011",5813 => "00010001",5814 => "01001000",5815 => "11101101",5816 => "01011001",5817 => "10100011",5818 => "11111110",5819 => "11101111",5820 => "11010101",5821 => "10100011",5822 => "00010110",5823 => "11011111",5824 => "00100001",5825 => "00110110",5826 => "01001010",5827 => "01100001",5828 => "00111011",5829 => "11011010",5830 => "00001000",5831 => "10010111",5832 => "01111001",5833 => "01011001",5834 => "10000011",5835 => "10001111",5836 => "10110011",5837 => "00011000",5838 => "00101001",5839 => "01011100",5840 => "01101101",5841 => "10100100",5842 => "00100010",5843 => "00000111",5844 => "01011100",5845 => "01110000",5846 => "00111001",5847 => "01001010",5848 => "00101011",5849 => "11110010",5850 => "01011000",5851 => "10111010",5852 => "00110010",5853 => "01011010",5854 => "10101010",5855 => "10011010",5856 => "00100001",5857 => "00100111",5858 => "10011001",5859 => "10001110",5860 => "11101111",5861 => "00001010",5862 => "00010101",5863 => "11001111",5864 => "00001111",5865 => "10100101",5866 => "00011011",5867 => "11101000",5868 => "01010110",5869 => "11111110",5870 => "01101000",5871 => "11001010",5872 => "00111111",5873 => "00101011",5874 => "10110101",5875 => "10001111",5876 => "00001110",5877 => "01110011",5878 => "01110110",5879 => "00010100",5880 => "11011010",5881 => "10110100",5882 => "10011000",5883 => "00001100",5884 => "01110001",5885 => "01111000",5886 => "10010010",5887 => "01111110",5888 => "10111010",5889 => "10001000",5890 => "11000100",5891 => "00100001",5892 => "11110001",5893 => "10001000",5894 => "11111010",5895 => "01001001",5896 => "11010110",5897 => "01011110",5898 => "10110000",5899 => "00011011",5900 => "11101000",5901 => "00001000",5902 => "00101010",5903 => "11110111",5904 => "11000011",5905 => "11000101",5906 => "11011011",5907 => "00010011",5908 => "10011111",5909 => "01111010",5910 => "10000001",5911 => "01110011",5912 => "11010001",5913 => "01111111",5914 => "11011010",5915 => "00101111",5916 => "00001001",5917 => "00000101",5918 => "10101000",5919 => "00011000",5920 => "00101100",5921 => "01111000",5922 => "11010110",5923 => "11100100",5924 => "11000000",5925 => "01101101",5926 => "00011010",5927 => "00010000",5928 => "10011110",5929 => "00111101",5930 => "10010101",5931 => "00111001",5932 => "00011110",5933 => "10101111",5934 => "11110001",5935 => "11100101",5936 => "11111110",5937 => "11101110",5938 => "11010101",5939 => "10111001",5940 => "10001110",5941 => "10110001",5942 => "00001011",5943 => "10101100",5944 => "00000011",5945 => "10010000",5946 => "01111010",5947 => "11101001",5948 => "01000011",5949 => "00100100",5950 => "10011011",5951 => "10000010",5952 => "01010110",5953 => "00011111",5954 => "10011111",5955 => "00011011",5956 => "10000001",5957 => "10000001",5958 => "10011110",5959 => "01100010",5960 => "11010011",5961 => "01111001",5962 => "01001100",5963 => "10100110",5964 => "01010011",5965 => "11011000",5966 => "00000110",5967 => "11101011",5968 => "01100110",5969 => "10101101",5970 => "00000111",5971 => "00110000",5972 => "10101010",5973 => "11000101",5974 => "01110110",5975 => "11100111",5976 => "11100001",5977 => "00110100",5978 => "01000111",5979 => "01111101",5980 => "11101111",5981 => "01111001",5982 => "11100100",5983 => "10111000",5984 => "00100101",5985 => "00110110",5986 => "10101111",5987 => "00101011",5988 => "00001000",5989 => "10010110",5990 => "11001111",5991 => "00101001",5992 => "10101011",5993 => "01001000",5994 => "01100101",5995 => "10001100",5996 => "01000101",5997 => "10101111",5998 => "10001110",5999 => "01111000",6000 => "11101110",6001 => "00110010",6002 => "01100110",6003 => "01101101",6004 => "10001110",6005 => "10000101",6006 => "10001000",6007 => "11111100",6008 => "01101100",6009 => "10001100",6010 => "01010100",6011 => "10000000",6012 => "00001001",6013 => "10001100",6014 => "01101111",6015 => "01001111",6016 => "01110100",6017 => "11101110",6018 => "11101000",6019 => "01000110",6020 => "00001000",6021 => "10101101",6022 => "00101111",6023 => "01110101",6024 => "00000000",6025 => "11110000",6026 => "01100010",6027 => "01000101",6028 => "11101101",6029 => "00111000",6030 => "00010111",6031 => "01100111",6032 => "10100000",6033 => "10111011",6034 => "10000010",6035 => "10011000",6036 => "11000011",6037 => "10100110",6038 => "00101111",6039 => "01110101",6040 => "11011101",6041 => "00100001",6042 => "01000111",6043 => "10100100",6044 => "11000110",6045 => "10000001",6046 => "01000001",6047 => "11010100",6048 => "01011000",6049 => "10101011",6050 => "11110011",6051 => "01011110",6052 => "01101010",6053 => "10111110",6054 => "01011011",6055 => "00100000",6056 => "00000111",6057 => "00100001",6058 => "01111001",6059 => "11100110",6060 => "01001000",6061 => "00011100",6062 => "01011100",6063 => "00001001",6064 => "11000000",6065 => "10011000",6066 => "11001110",6067 => "11111110",6068 => "00111010",6069 => "00000010",6070 => "11001010",6071 => "11011011",6072 => "00010000",6073 => "11101111",6074 => "10101110",6075 => "10011101",6076 => "01000111",6077 => "01000101",6078 => "00011100",6079 => "00101011",6080 => "01101110",6081 => "11101001",6082 => "01010000",6083 => "11000111",6084 => "01101011",6085 => "10110011",6086 => "00011100",6087 => "10110111",6088 => "01100000",6089 => "00100100",6090 => "10010001",6091 => "00110011",6092 => "11101111",6093 => "10111110",6094 => "00110000",6095 => "11110010",6096 => "01101001",6097 => "10110110",6098 => "01011100",6099 => "01000100",6100 => "10101001",6101 => "11100011",6102 => "00101011",6103 => "01101101",6104 => "01000101",6105 => "01110000",6106 => "11110000",6107 => "10001101",6108 => "11101101",6109 => "01100111",6110 => "00001001",6111 => "11110110",6112 => "10010010",6113 => "10110101",6114 => "00101011",6115 => "11010011",6116 => "01000000",6117 => "00111110",6118 => "11111000",6119 => "01111011",6120 => "11110110",6121 => "10101010",6122 => "01110111",6123 => "10000011",6124 => "11101100",6125 => "10100100",6126 => "00111000",6127 => "01001001",6128 => "11000000",6129 => "11000000",6130 => "00011101",6131 => "10100101",6132 => "11111011",6133 => "11111110",6134 => "10110111",6135 => "11111011",6136 => "10000110",6137 => "11101011",6138 => "01101011",6139 => "10111010",6140 => "00011101",6141 => "00111011",6142 => "00100110",6143 => "01101111",6144 => "10001001",6145 => "00000000",6146 => "01100101",6147 => "00100010",6148 => "00000001",6149 => "00100001",6150 => "01100110",6151 => "11100110",6152 => "11010001",6153 => "11110010",6154 => "11000001",6155 => "01011111",6156 => "10001110",6157 => "01000110",6158 => "01101001",6159 => "10011110",6160 => "11010000",6161 => "11010101",6162 => "11011001",6163 => "11100000",6164 => "10110110",6165 => "10011001",6166 => "00010000",6167 => "00110100",6168 => "11110111",6169 => "10010101",6170 => "11101001",6171 => "01010110",6172 => "10000110",6173 => "11010111",6174 => "11100010",6175 => "00000110",6176 => "11010001",6177 => "00110001",6178 => "00000011",6179 => "00100001",6180 => "00101010",6181 => "11100111",6182 => "00110110",6183 => "00001101",6184 => "01011011",6185 => "11011011",6186 => "11101111",6187 => "01011100",6188 => "10000001",6189 => "00011001",6190 => "01100100",6191 => "11000001",6192 => "01000101",6193 => "11101111",6194 => "00001011",6195 => "11101110",6196 => "11010101",6197 => "10001011",6198 => "10101100",6199 => "00110101",6200 => "00110010",6201 => "11100011",6202 => "10000010",6203 => "01111111",6204 => "10000101",6205 => "10101111",6206 => "10000011",6207 => "01011011",6208 => "00011011",6209 => "10010011",6210 => "11001100",6211 => "00001110",6212 => "01010001",6213 => "00110011",6214 => "10011100",6215 => "10111101",6216 => "01001010",6217 => "00100011",6218 => "10010011",6219 => "00000010",6220 => "10001011",6221 => "01111001",6222 => "11010011",6223 => "10011101",6224 => "11110110",6225 => "01010011",6226 => "01110010",6227 => "11111100",6228 => "01001001",6229 => "01011101",6230 => "00101010",6231 => "11110100",6232 => "01000011",6233 => "11001100",6234 => "01110111",6235 => "11010100",6236 => "11100100",6237 => "01101111",6238 => "01110011",6239 => "01000001",6240 => "01001101",6241 => "01011110",6242 => "00001111",6243 => "10111011",6244 => "11111100",6245 => "10111100",6246 => "10101000",6247 => "01110001",6248 => "11111101",6249 => "10010001",6250 => "11000101",6251 => "11110010",6252 => "10001000",6253 => "00110010",6254 => "11011100",6255 => "00010111",6256 => "10010011",6257 => "00001010",6258 => "01001100",6259 => "11000000",6260 => "11111001",6261 => "01010000",6262 => "01000001",6263 => "11011111",6264 => "10111111",6265 => "00010000",6266 => "11101110",6267 => "01000101",6268 => "01011000",6269 => "01000010",6270 => "11101101",6271 => "11000101",6272 => "11001011",6273 => "00110101",6274 => "11100100",6275 => "01011000",6276 => "00101011",6277 => "10101111",6278 => "01100101",6279 => "10011010",6280 => "11000001",6281 => "00110011",6282 => "11000011",6283 => "00010110",6284 => "10111001",6285 => "01011011",6286 => "00101110",6287 => "11001001",6288 => "10011101",6289 => "01000011",6290 => "10101011",6291 => "01001100",6292 => "00011011",6293 => "00101100",6294 => "10110011",6295 => "10110110",6296 => "11110110",6297 => "11110111",6298 => "10100000",6299 => "10011011",6300 => "01000011",6301 => "11010100",6302 => "10111100",6303 => "10101100",6304 => "01011110",6305 => "01001111",6306 => "00100011",6307 => "10110111",6308 => "00100011",6309 => "11101011",6310 => "00011110",6311 => "11100000",6312 => "10011011",6313 => "01111011",6314 => "10110011",6315 => "10110100",6316 => "01100010",6317 => "11011110",6318 => "00110101",6319 => "00000100",6320 => "01011110",6321 => "00100000",6322 => "00000101",6323 => "00001001",6324 => "00110001",6325 => "11101100",6326 => "10011101",6327 => "00111001",6328 => "00111100",6329 => "10001001",6330 => "10011110",6331 => "10111110",6332 => "11100011",6333 => "10010100",6334 => "01110110",6335 => "00110111",6336 => "01101010",6337 => "11001101",6338 => "01100100",6339 => "10110101",6340 => "00010111",6341 => "01111001",6342 => "11010101",6343 => "01011111",6344 => "00000001",6345 => "11000111",6346 => "10101101",6347 => "00011000",6348 => "11011101",6349 => "01110111",6350 => "11110011",6351 => "01001111",6352 => "11111001",6353 => "01001010",6354 => "10011111",6355 => "01100100",6356 => "10101100",6357 => "00101101",6358 => "01101101",6359 => "00110000",6360 => "10010100",6361 => "01101010",6362 => "01111011",6363 => "10111010",6364 => "10011011",6365 => "01100011",6366 => "10010000",6367 => "11111110",6368 => "00011110",6369 => "00111101",6370 => "01111110",6371 => "01100100",6372 => "10010001",6373 => "11011100",6374 => "10110110",6375 => "11110011",6376 => "10111000",6377 => "11110101",6378 => "11000100",6379 => "11001011",6380 => "00010011",6381 => "11100100",6382 => "00101001",6383 => "11110100",6384 => "01100000",6385 => "00101011",6386 => "00111010",6387 => "01111101",6388 => "01110101",6389 => "01110000",6390 => "01110110",6391 => "00111010",6392 => "11111110",6393 => "11010011",6394 => "10111011",6395 => "00010110",6396 => "01010001",6397 => "10100100",6398 => "10001011",6399 => "11101100",6400 => "10001111",6401 => "01110001",6402 => "10101101",6403 => "00001100",6404 => "10110000",6405 => "10101110",6406 => "10111011",6407 => "10001000",6408 => "00111010",6409 => "10001101",6410 => "10101100",6411 => "00001010",6412 => "00000100",6413 => "11001000",6414 => "00000110",6415 => "01001111",6416 => "11001000",6417 => "01010010",6418 => "11001011",6419 => "10001001",6420 => "01001100",6421 => "10110111",6422 => "01011101",6423 => "01101101",6424 => "00111001",6425 => "01000000",6426 => "01110110",6427 => "11110101",6428 => "00101111",6429 => "10001110",6430 => "10100111",6431 => "11101001",6432 => "01011110",6433 => "11100110",6434 => "00100111",6435 => "11101001",6436 => "00101111",6437 => "01100000",6438 => "00111111",6439 => "01010011",6440 => "00111110",6441 => "01100111",6442 => "01101100",6443 => "01111011",6444 => "01110011",6445 => "11000101",6446 => "11110100",6447 => "10101011",6448 => "01000001",6449 => "00101110",6450 => "11010111",6451 => "00011011",6452 => "10010101",6453 => "11001010",6454 => "00000100",6455 => "10001101",6456 => "11011110",6457 => "10101111",6458 => "00101000",6459 => "01110010",6460 => "00110101",6461 => "00001001",6462 => "10101100",6463 => "11010001",6464 => "10101011",6465 => "10110110",6466 => "00011101",6467 => "10001011",6468 => "01010101",6469 => "00111100",6470 => "01011010",6471 => "00100100",6472 => "10111001",6473 => "11100111",6474 => "11011000",6475 => "00000111",6476 => "00111011",6477 => "10001100",6478 => "00010001",6479 => "01101111",6480 => "00011100",6481 => "01111111",6482 => "00110000",6483 => "00000011",6484 => "10001011",6485 => "10010111",6486 => "11100010",6487 => "00011010",6488 => "10001100",6489 => "01110010",6490 => "01100000",6491 => "10101001",6492 => "10101111",6493 => "00111111",6494 => "11010000",6495 => "10101111",6496 => "00110000",6497 => "10010010",6498 => "01010001",6499 => "10111011",6500 => "10100111",6501 => "01000110",6502 => "11000001",6503 => "00001010",6504 => "00010110",6505 => "00010000",6506 => "11000001",6507 => "00110000",6508 => "00101011",6509 => "01111101",6510 => "01010101",6511 => "11100100",6512 => "10100111",6513 => "11001111",6514 => "10101100",6515 => "10110001",6516 => "10001100",6517 => "00010100",6518 => "11101000",6519 => "01111100",6520 => "11010000",6521 => "01010000",6522 => "11100011",6523 => "11000010",6524 => "01000111",6525 => "01000110",6526 => "10000011",6527 => "10000100",6528 => "00011110",6529 => "11111011",6530 => "00101011",6531 => "10110010",6532 => "11101110",6533 => "00101100",6534 => "01100010",6535 => "11011111",6536 => "10100000",6537 => "11011100",6538 => "01100100",6539 => "11001110",6540 => "11001101",6541 => "00111101",6542 => "00110011",6543 => "11011000",6544 => "00110010",6545 => "10010010",6546 => "10111101",6547 => "10000110",6548 => "00001000",6549 => "01010100",6550 => "00001110",6551 => "11101000",6552 => "01001111",6553 => "00110000",6554 => "00010101",6555 => "11000100",6556 => "10010001",6557 => "11101110",6558 => "11011001",6559 => "11001011",6560 => "01000001",6561 => "10000100",6562 => "11111001",6563 => "00010000",6564 => "11000011",6565 => "01111000",6566 => "01011001",6567 => "11001100",6568 => "00111100",6569 => "10001100",6570 => "10100110",6571 => "10110111",6572 => "11100001",6573 => "11001111",6574 => "00110101",6575 => "01100101",6576 => "00100000",6577 => "10110101",6578 => "01111100",6579 => "11001111",6580 => "00100100",6581 => "10101101",6582 => "01011110",6583 => "00111111",6584 => "01001100",6585 => "01000101",6586 => "10110000",6587 => "10111100",6588 => "10110111",6589 => "11101001",6590 => "11001000",6591 => "01001101",6592 => "10111010",6593 => "00100001",6594 => "00111000",6595 => "01110011",6596 => "00010111",6597 => "01110001",6598 => "01101000",6599 => "10101001",6600 => "00011000",6601 => "01100111",6602 => "01011010",6603 => "00000010",6604 => "00011110",6605 => "01100111",6606 => "01010111",6607 => "00011010",6608 => "11000100",6609 => "11101001",6610 => "11010111",6611 => "01110101",6612 => "00111111",6613 => "01100010",6614 => "01101011",6615 => "01100001",6616 => "10000111",6617 => "01110001",6618 => "11000111",6619 => "00001010",6620 => "01000101",6621 => "00100110",6622 => "01100110",6623 => "11111000",6624 => "00011011",6625 => "10001110",6626 => "11010000",6627 => "01100101",6628 => "11000001",6629 => "11110011",6630 => "01010001",6631 => "11001101",6632 => "10001100",6633 => "10010001",6634 => "11000000",6635 => "10111101",6636 => "00001111",6637 => "01001001",6638 => "01100110",6639 => "00000010",6640 => "00001001",6641 => "01000100",6642 => "10011100",6643 => "11000010",6644 => "00100000",6645 => "11100100",6646 => "11011001",6647 => "00110110",6648 => "11101001",6649 => "10011100",6650 => "01111000",6651 => "11010111",6652 => "01010000",6653 => "11011001",6654 => "00011111",6655 => "11000000",6656 => "11111101",6657 => "10100001",6658 => "00011011",6659 => "11110010",6660 => "00001111",6661 => "00000000",6662 => "00000000",6663 => "00111100",6664 => "00000101",6665 => "01111011",6666 => "00000111",6667 => "11010100",6668 => "01010110",6669 => "01010100",6670 => "11110111",6671 => "01010110",6672 => "11000011",6673 => "00100100",6674 => "10100011",6675 => "11000010",6676 => "01010011",6677 => "10010111",6678 => "11100000",6679 => "11111011",6680 => "11110000",6681 => "01111010",6682 => "00100010",6683 => "10010011",6684 => "01000011",6685 => "10001101",6686 => "00001010",6687 => "11011100",6688 => "10010101",6689 => "01101000",6690 => "00100001",6691 => "11111010",6692 => "10011001",6693 => "00010011",6694 => "01101111",6695 => "11000101",6696 => "00100101",6697 => "00101000",6698 => "01100011",6699 => "01101100",6700 => "10110001",6701 => "11100011",6702 => "10111100",6703 => "10010101",6704 => "11100010",6705 => "00100010",6706 => "11011000",6707 => "10110001",6708 => "11001000",6709 => "00000111",6710 => "01000111",6711 => "10000000",6712 => "00100000",6713 => "01011101",6714 => "10110001",6715 => "11100000",6716 => "00011000",6717 => "11111101",6718 => "11010101",6719 => "01101100",6720 => "10011000",6721 => "11101100",6722 => "11110011",6723 => "10111001",6724 => "01000100",6725 => "01010011",6726 => "10111010",6727 => "01011100",6728 => "11110000",6729 => "00000000",6730 => "11100011",6731 => "01010010",6732 => "01111110",6733 => "01011011",6734 => "01110001",6735 => "10010110",6736 => "10101100",6737 => "11010111",6738 => "01100011",6739 => "10110010",6740 => "10100010",6741 => "10011001",6742 => "11010101",6743 => "10100110",6744 => "00101000",6745 => "10101110",6746 => "00001010",6747 => "10001111",6748 => "10011100",6749 => "10110001",6750 => "00101000",6751 => "01011111",6752 => "00000001",6753 => "10000010",6754 => "11001001",6755 => "01111111",6756 => "00000010",6757 => "10101000",6758 => "00001010",6759 => "11001111",6760 => "01100100",6761 => "11010110",6762 => "10110010",6763 => "00011001",6764 => "10110111",6765 => "10000010",6766 => "00111111",6767 => "11110001",6768 => "00010101",6769 => "11110011",6770 => "11011101",6771 => "00111011",6772 => "10011010",6773 => "00111010",6774 => "10011001",6775 => "10001101",6776 => "11110111",6777 => "01110111",6778 => "01111110",6779 => "01000010",6780 => "10010011",6781 => "00100000",6782 => "10100100",6783 => "01101011",6784 => "01001011",6785 => "11000111",6786 => "00101110",6787 => "01110110",6788 => "01000101",6789 => "01000000",6790 => "11110100",6791 => "01110101",6792 => "10000101",6793 => "00010000",6794 => "01010111",6795 => "10101111",6796 => "10001110",6797 => "00111111",6798 => "10100011",6799 => "11000111",6800 => "10110110",6801 => "11010001",6802 => "10000110",6803 => "11111100",6804 => "00111000",6805 => "00010000",6806 => "00000100",6807 => "01110011",6808 => "10000001",6809 => "11001001",6810 => "10111010",6811 => "11100101",6812 => "00110010",6813 => "00011100",6814 => "00000111",6815 => "00101001",6816 => "01001100",6817 => "11010101",6818 => "00010100",6819 => "10010110",6820 => "00001110",6821 => "00110011",6822 => "00011001",6823 => "01000100",6824 => "01101100",6825 => "01000101",6826 => "00011111",6827 => "01101100",6828 => "10000111",6829 => "10101100",6830 => "00001101",6831 => "11111111",6832 => "11100001",6833 => "00001000",6834 => "11010110",6835 => "00000011",6836 => "00011000",6837 => "01011101",6838 => "11010011",6839 => "00000001",6840 => "01010110",6841 => "00010111",6842 => "11110111",6843 => "10111101",6844 => "11000000",6845 => "01000011",6846 => "10000010",6847 => "10010100",6848 => "01011001",6849 => "11111110",6850 => "11001110",6851 => "11001110",6852 => "11000101",6853 => "01000000",6854 => "00110101",6855 => "01001000",6856 => "11100011",6857 => "00011100",6858 => "10001010",6859 => "10010000",6860 => "11100010",6861 => "01011010",6862 => "11111011",6863 => "01000111",6864 => "01010110",6865 => "10101111",6866 => "10100101",6867 => "00111011",6868 => "10100110",6869 => "11010000",6870 => "11000111",6871 => "01001111",6872 => "10010001",6873 => "00100011",6874 => "01010110",6875 => "00111000",6876 => "00011111",6877 => "11001110",6878 => "00101001",6879 => "01011110",6880 => "10010001",6881 => "00100101",6882 => "11110010",6883 => "00100011",6884 => "01001111",6885 => "11010011",6886 => "11000100",6887 => "01010110",6888 => "00111110",6889 => "10101000",6890 => "10011001",6891 => "11001110",6892 => "10110100",6893 => "00100111",6894 => "10101011",6895 => "10000101",6896 => "00001010",6897 => "00000110",6898 => "11001000",6899 => "01000110",6900 => "10100111",6901 => "00010100",6902 => "11110000",6903 => "11000111",6904 => "11110111",6905 => "10011000",6906 => "01001111",6907 => "00100010",6908 => "00110011",6909 => "10101010",6910 => "11011101",6911 => "10111110",6912 => "11110101",6913 => "00010010",6914 => "00101111",6915 => "10000100",6916 => "01010000",6917 => "00000010",6918 => "01110010",6919 => "10010000",6920 => "01000110",6921 => "10111110",6922 => "10101001",6923 => "00111010",6924 => "01100101",6925 => "11110010",6926 => "11101011",6927 => "11100001",6928 => "00110010",6929 => "10011101",6930 => "11001110",6931 => "10110101",6932 => "01000111",6933 => "00110101",6934 => "10111110",6935 => "11001010",6936 => "01010010",6937 => "01100010",6938 => "10101100",6939 => "00001010",6940 => "10000100",6941 => "10000010",6942 => "11101100",6943 => "00101011",6944 => "11011001",6945 => "00100001",6946 => "11101101",6947 => "10111000",6948 => "00100111",6949 => "10000001",6950 => "01000111",6951 => "11110000",6952 => "11101001",6953 => "01101110",6954 => "00000010",6955 => "00010100",6956 => "10100101",6957 => "11000010",6958 => "11011001",6959 => "01011011",6960 => "00010001",6961 => "10101001",6962 => "01010101",6963 => "11001111",6964 => "10010101",6965 => "01011111",6966 => "00011100",6967 => "01101101",6968 => "01001001",6969 => "01111011",6970 => "11101101",6971 => "10111010",6972 => "11001001",6973 => "11111110",6974 => "00000110",6975 => "11100000",6976 => "11001011",6977 => "00111100",6978 => "01011011",6979 => "10101100",6980 => "00000101",6981 => "11100101",6982 => "00101001",6983 => "01100001",6984 => "10010011",6985 => "10011000",6986 => "01111000",6987 => "11001011",6988 => "01011000",6989 => "00001010",6990 => "01011010",6991 => "10111010",6992 => "01111110",6993 => "01111110",6994 => "01110011",6995 => "10100000",6996 => "01101010",6997 => "01001110",6998 => "00000011",6999 => "10110000",7000 => "01001100",7001 => "11101100",7002 => "00111001",7003 => "00000100",7004 => "01000101",7005 => "10100110",7006 => "00001100",7007 => "00001000",7008 => "01011110",7009 => "11101000",7010 => "00000010",7011 => "01001011",7012 => "01111100",7013 => "00101010",7014 => "00010000",7015 => "11000000",7016 => "01111111",7017 => "01010111",7018 => "11110001",7019 => "11011000",7020 => "10001011",7021 => "01000001",7022 => "10010010",7023 => "00100000",7024 => "11111011",7025 => "10011001",7026 => "10011000",7027 => "10110010",7028 => "10101011",7029 => "01001110",7030 => "11001000",7031 => "10011101",7032 => "00110011",7033 => "00011000",7034 => "10001000",7035 => "00000010",7036 => "00010000",7037 => "00001000",7038 => "01110110",7039 => "10000110",7040 => "10101000",7041 => "01111111",7042 => "00001111",7043 => "00001001",7044 => "00000000",7045 => "00011001",7046 => "10000010",7047 => "10111110",7048 => "00010101",7049 => "01000011",7050 => "11110100",7051 => "01010000",7052 => "10011010",7053 => "10000010",7054 => "10010100",7055 => "00001000",7056 => "10000111",7057 => "00111100",7058 => "11110010",7059 => "11101101",7060 => "10010110",7061 => "10011111",7062 => "11110010",7063 => "10011001",7064 => "00010111",7065 => "11101000",7066 => "01100111",7067 => "00110110",7068 => "00001111",7069 => "00001101",7070 => "00010110",7071 => "00111111",7072 => "00101101",7073 => "11100100",7074 => "11100110",7075 => "11011110",7076 => "10000111",7077 => "11001111",7078 => "10111001",7079 => "11011011",7080 => "10011100",7081 => "11101000",7082 => "01001110",7083 => "00110111",7084 => "10111000",7085 => "00110110",7086 => "00111000",7087 => "11111100",7088 => "10001101",7089 => "11000001",7090 => "10101001",7091 => "00101110",7092 => "01010111",7093 => "10001010",7094 => "00110001",7095 => "11001001",7096 => "11111001",7097 => "10101010",7098 => "11001010",7099 => "00011011",7100 => "10100000",7101 => "01000000",7102 => "01000101",7103 => "01100011",7104 => "10001001",7105 => "11110101",7106 => "00111010",7107 => "01001101",7108 => "10000101",7109 => "01010111",7110 => "11001001",7111 => "10010000",7112 => "10111111",7113 => "01101000",7114 => "10010110",7115 => "11101000",7116 => "01001110",7117 => "10110010",7118 => "00001101",7119 => "10010010",7120 => "01100110",7121 => "11111000",7122 => "11110111",7123 => "01110100",7124 => "00100110",7125 => "00101000",7126 => "11111100",7127 => "10111101",7128 => "10010010",7129 => "10111011",7130 => "00000101",7131 => "11100110",7132 => "01000101",7133 => "01010111",7134 => "10011101",7135 => "10101010",7136 => "10011111",7137 => "00011011",7138 => "01100111",7139 => "01110100",7140 => "01010101",7141 => "11100010",7142 => "01010001",7143 => "00101001",7144 => "00010101",7145 => "01001110",7146 => "00011111",7147 => "01111101",7148 => "01101000",7149 => "00100110",7150 => "01111110",7151 => "11101110",7152 => "01010001",7153 => "00011011",7154 => "01100001",7155 => "01001011",7156 => "01110001",7157 => "01011100",7158 => "11101001",7159 => "00110000",7160 => "11110100",7161 => "01011011",7162 => "10000010",7163 => "11111100",7164 => "00101110",7165 => "01010001",7166 => "11110010",7167 => "10110000",7168 => "11101110",7169 => "01100001",7170 => "00000010",7171 => "01001001",7172 => "00111111",7173 => "00101000",7174 => "11101110",7175 => "00110101",7176 => "00111101",7177 => "11100111",7178 => "01110100",7179 => "00011110",7180 => "01001001",7181 => "01101101",7182 => "10100111",7183 => "10101100",7184 => "10101010",7185 => "11011011",7186 => "01101111",7187 => "10010010",7188 => "01100011",7189 => "10111001",7190 => "01000100",7191 => "00000011",7192 => "11001001",7193 => "11001110",7194 => "10101011",7195 => "10111110",7196 => "11100111",7197 => "00000101",7198 => "00000111",7199 => "00100000",7200 => "10001101",7201 => "01111101",7202 => "00011101",7203 => "01100001",7204 => "11011110",7205 => "11010000",7206 => "10001001",7207 => "00100111",7208 => "00100011",7209 => "00011110",7210 => "01110111",7211 => "10100111",7212 => "11011001",7213 => "00111001",7214 => "11101110",7215 => "10111111",7216 => "10110100",7217 => "10000110",7218 => "00101100",7219 => "11010001",7220 => "01011100",7221 => "11100110",7222 => "01110000",7223 => "11000000",7224 => "10110011",7225 => "00011111",7226 => "00011000",7227 => "11011110",7228 => "10100001",7229 => "11011100",7230 => "11111101",7231 => "11010011",7232 => "11100111",7233 => "00111011",7234 => "00001000",7235 => "00000101",7236 => "10001011",7237 => "11110000",7238 => "01000110",7239 => "11100111",7240 => "10101000",7241 => "10101001",7242 => "11111001",7243 => "10001101",7244 => "11011111",7245 => "11111010",7246 => "00010100",7247 => "01010111",7248 => "01001000",7249 => "10101001",7250 => "00000000",7251 => "00010011",7252 => "10011001",7253 => "00010001",7254 => "11010001",7255 => "00100101",7256 => "01011101",7257 => "01111011",7258 => "01001100",7259 => "11000000",7260 => "00011101",7261 => "11000111",7262 => "01000000",7263 => "01111001",7264 => "01001110",7265 => "00101101",7266 => "01010000",7267 => "11000110",7268 => "10111011",7269 => "11101100",7270 => "00011100",7271 => "10101100",7272 => "00001000",7273 => "01111111",7274 => "01100001",7275 => "01001111",7276 => "11010000",7277 => "00010101",7278 => "10000001",7279 => "00001000",7280 => "10100110",7281 => "01110001",7282 => "00010011",7283 => "11101010",7284 => "01000011",7285 => "01110101",7286 => "10011101",7287 => "01111100",7288 => "10111110",7289 => "11011001",7290 => "01101001",7291 => "10001110",7292 => "10001111",7293 => "01011101",7294 => "00101100",7295 => "11001110",7296 => "11011110",7297 => "10110110",7298 => "10001100",7299 => "11010010",7300 => "00111100",7301 => "10001010",7302 => "01101111",7303 => "11011001",7304 => "01000011",7305 => "11011011",7306 => "00001101",7307 => "01100111",7308 => "11000001",7309 => "10111111",7310 => "11110100",7311 => "10101010",7312 => "01110111",7313 => "00000011",7314 => "00011101",7315 => "01110110",7316 => "10011001",7317 => "00111011",7318 => "01000001",7319 => "11010001",7320 => "11110110",7321 => "11111001",7322 => "11000101",7323 => "10000000",7324 => "01100101",7325 => "10111101",7326 => "11001011",7327 => "00011011",7328 => "10000100",7329 => "11100101",7330 => "10010000",7331 => "01110100",7332 => "11100011",7333 => "10011000",7334 => "11011001",7335 => "11011011",7336 => "11110001",7337 => "10001010",7338 => "11001011",7339 => "01001110",7340 => "00110111",7341 => "01100110",7342 => "10010101",7343 => "00110011",7344 => "10101100",7345 => "00010100",7346 => "01011001",7347 => "10100111",7348 => "11100011",7349 => "10110001",7350 => "11110110",7351 => "00111110",7352 => "00001111",7353 => "01101110",7354 => "10101110",7355 => "11010101",7356 => "01100001",7357 => "10111011",7358 => "00110111",7359 => "00011001",7360 => "00010001",7361 => "10100110",7362 => "01000100",7363 => "11110010",7364 => "01100101",7365 => "00101100",7366 => "01010111",7367 => "11001001",7368 => "01101110",7369 => "10110100",7370 => "10010000",7371 => "01101100",7372 => "10101000",7373 => "11010010",7374 => "11111000",7375 => "10101011",7376 => "00011101",7377 => "11001010",7378 => "10101101",7379 => "10001100",7380 => "10101101",7381 => "00001010",7382 => "00101010",7383 => "00101010",7384 => "11111010",7385 => "00000101",7386 => "10100101",7387 => "00000011",7388 => "00000000",7389 => "00001100",7390 => "11111110",7391 => "10001111",7392 => "10110110",7393 => "01000101",7394 => "10110101",7395 => "10111000",7396 => "00100010",7397 => "00111100",7398 => "00110111",7399 => "10100101",7400 => "01011011",7401 => "10011011",7402 => "00110111",7403 => "01110010",7404 => "10100111",7405 => "10111000",7406 => "00111100",7407 => "00100011",7408 => "10110110",7409 => "10010011",7410 => "01010110",7411 => "00010000",7412 => "10111110",7413 => "01010101",7414 => "10001000",7415 => "00010010",7416 => "10110101",7417 => "10110001",7418 => "01101101",7419 => "01000000",7420 => "00010000",7421 => "11110100",7422 => "11111100",7423 => "10100011",7424 => "10011110",7425 => "10001011",7426 => "10000000",7427 => "11011111",7428 => "01101001",7429 => "00000010",7430 => "01101010",7431 => "11100011",7432 => "11101110",7433 => "11000001",7434 => "11110111",7435 => "01101110",7436 => "11110011",7437 => "10101111",7438 => "01111111",7439 => "11100000",7440 => "10001010",7441 => "11101111",7442 => "00101000",7443 => "11011011",7444 => "00110100",7445 => "01000101",7446 => "00010001",7447 => "01000001",7448 => "01000111",7449 => "10110101",7450 => "00011111",7451 => "00100000",7452 => "10111010",7453 => "01001001",7454 => "11101011",7455 => "01010000",7456 => "01110101",7457 => "00000101",7458 => "10110100",7459 => "10110100",7460 => "01001111",7461 => "11111011",7462 => "01001111",7463 => "01001110",7464 => "01010011",7465 => "10001011",7466 => "00101110",7467 => "00100110",7468 => "00101010",7469 => "01011111",7470 => "00001011",7471 => "11111011",7472 => "01001011",7473 => "01010110",7474 => "00010011",7475 => "00001001",7476 => "00111111",7477 => "00100001",7478 => "01010111",7479 => "11100001",7480 => "01000100",7481 => "01110001",7482 => "10001010",7483 => "01001011",7484 => "00111011",7485 => "11011010",7486 => "10001111",7487 => "01001001",7488 => "00111101",7489 => "00011110",7490 => "11000011",7491 => "11101000",7492 => "01010101",7493 => "10001110",7494 => "01010010",7495 => "11000110",7496 => "01100110",7497 => "10010011",7498 => "00101010",7499 => "10000000",7500 => "01010100",7501 => "00011111",7502 => "01011001",7503 => "10000100",7504 => "01101001",7505 => "01001011",7506 => "01010011",7507 => "01000001",7508 => "00001101",7509 => "01010110",7510 => "11100010",7511 => "10011111",7512 => "01101111",7513 => "11110011",7514 => "11011110",7515 => "00110011",7516 => "11001100",7517 => "01100001",7518 => "11110010",7519 => "00111010",7520 => "01011000",7521 => "01110110",7522 => "10100101",7523 => "00011011",7524 => "00100010",7525 => "11001011",7526 => "01011100",7527 => "10000010",7528 => "00011111",7529 => "01101001",7530 => "10110100",7531 => "00111011",7532 => "00010001",7533 => "01011100",7534 => "00101111",7535 => "11001101",7536 => "10111010",7537 => "10010111",7538 => "00001101",7539 => "00010110",7540 => "01101100",7541 => "10001110",7542 => "11100101",7543 => "11100101",7544 => "00101110",7545 => "01110111",7546 => "11101001",7547 => "01001010",7548 => "01100001",7549 => "01111101",7550 => "00101011",7551 => "11100111",7552 => "00110001",7553 => "00101111",7554 => "00101000",7555 => "00110100",7556 => "10011100",7557 => "00000110",7558 => "11100100",7559 => "00010101",7560 => "01011011",7561 => "10011000",7562 => "10001001",7563 => "00101111",7564 => "11011100",7565 => "00011110",7566 => "10111110",7567 => "10111111",7568 => "11000010",7569 => "00000010",7570 => "11111001",7571 => "00110111",7572 => "10010010",7573 => "01111100",7574 => "01001001",7575 => "11000111",7576 => "11010100",7577 => "00011110",7578 => "11000000",7579 => "00000000",7580 => "11101110",7581 => "11111001",7582 => "10001111",7583 => "10011111",7584 => "10001011",7585 => "10000000",7586 => "11111010",7587 => "10101110",7588 => "11001101",7589 => "00110100",7590 => "00001011",7591 => "10101010",7592 => "00111001",7593 => "10001111",7594 => "01100011",7595 => "10100001",7596 => "01000011",7597 => "10010001",7598 => "11101000",7599 => "01110110",7600 => "10000100",7601 => "11111000",7602 => "11110111",7603 => "11110100",7604 => "11000010",7605 => "01010011",7606 => "10111110",7607 => "01100101",7608 => "00010101",7609 => "10100000",7610 => "01010001",7611 => "01100011",7612 => "01011001",7613 => "01001010",7614 => "00111011",7615 => "10100010",7616 => "10001001",7617 => "11000100",7618 => "11111110",7619 => "11010010",7620 => "00110111",7621 => "00011010",7622 => "01111000",7623 => "00011011",7624 => "01001111",7625 => "01100000",7626 => "00000011",7627 => "10100101",7628 => "00111010",7629 => "01111001",7630 => "01001001",7631 => "10110010",7632 => "00110110",7633 => "10011000",7634 => "11111011",7635 => "00001110",7636 => "00111110",7637 => "01011101",7638 => "01111011",7639 => "01010001",7640 => "00101001",7641 => "01011110",7642 => "01101110",7643 => "11101111",7644 => "10000000",7645 => "01011011",7646 => "00111110",7647 => "00010100",7648 => "10100101",7649 => "11011000",7650 => "01010010",7651 => "00110000",7652 => "10100010",7653 => "11000011",7654 => "00010000",7655 => "00100110",7656 => "01010111",7657 => "10010110",7658 => "10011001",7659 => "10110111",7660 => "10010000",7661 => "11100110",7662 => "10010101",7663 => "11011100",7664 => "10010010",7665 => "11001100",7666 => "10000111",7667 => "10101001",7668 => "00100011",7669 => "10100010",7670 => "11111101",7671 => "00011001",7672 => "00011011",7673 => "01010101",7674 => "01111100",7675 => "10111101",7676 => "01000100",7677 => "00101101",7678 => "00110100",7679 => "11101001",7680 => "00100101",7681 => "01100111",7682 => "00011110",7683 => "11111101",7684 => "10011011",7685 => "11010110",7686 => "10110001",7687 => "01010111",7688 => "10101011",7689 => "11010011",7690 => "11100000",7691 => "10101100",7692 => "00000101",7693 => "00101001",7694 => "01011000",7695 => "11001110",7696 => "11011011",7697 => "10010010",7698 => "01100001",7699 => "11010101",7700 => "10011100",7701 => "01110110",7702 => "11011000",7703 => "10111000",7704 => "11111011",7705 => "00110000",7706 => "10000100",7707 => "01101001",7708 => "11100111",7709 => "11100001",7710 => "10000001",7711 => "01110111",7712 => "00000000",7713 => "11011100",7714 => "11111100",7715 => "00101001",7716 => "10111011",7717 => "11000000",7718 => "01000100",7719 => "01010100",7720 => "01100001",7721 => "11011000",7722 => "10100100",7723 => "01111001",7724 => "01011111",7725 => "01000000",7726 => "11100010",7727 => "10101000",7728 => "00111011",7729 => "01000100",7730 => "10001010",7731 => "11011101",7732 => "00100011",7733 => "11111101",7734 => "00010010",7735 => "01011001",7736 => "00000001",7737 => "00100000",7738 => "10011010",7739 => "11101000",7740 => "10111101",7741 => "11010110",7742 => "10100000",7743 => "10001111",7744 => "10001011",7745 => "11010110",7746 => "11100110",7747 => "00010001",7748 => "01100111",7749 => "11101010",7750 => "00111111",7751 => "00111000",7752 => "11110001",7753 => "11100111",7754 => "11101010",7755 => "10010111",7756 => "11101110",7757 => "10100010",7758 => "11101100",7759 => "00101100",7760 => "01001100",7761 => "10111111",7762 => "00011111",7763 => "00000001",7764 => "00011101",7765 => "00000011",7766 => "01101101",7767 => "00100010",7768 => "10110010",7769 => "11100010",7770 => "11101110",7771 => "01011001",7772 => "00001011",7773 => "01001011",7774 => "01111001",7775 => "01010010",7776 => "10100101",7777 => "00001101",7778 => "10100010",7779 => "01110010",7780 => "00010100",7781 => "00111010",7782 => "11000100",7783 => "01011010",7784 => "11101010",7785 => "10100001",7786 => "01011110",7787 => "11100000",7788 => "10011110",7789 => "11100101",7790 => "11100000",7791 => "00101011",7792 => "00011101",7793 => "11111110",7794 => "11110110",7795 => "01001011",7796 => "00101100",7797 => "00110101",7798 => "11101000",7799 => "01011010",7800 => "11010100",7801 => "00001101",7802 => "10110111",7803 => "11101001",7804 => "11110000",7805 => "01111010",7806 => "00001011",7807 => "11110100",7808 => "10010111",7809 => "00001110",7810 => "01001100",7811 => "00011010",7812 => "11011110",7813 => "11000101",7814 => "00111100",7815 => "11010001",7816 => "11011110",7817 => "11011111",7818 => "10111001",7819 => "11010000",7820 => "01010011",7821 => "10100101",7822 => "01101001",7823 => "11100101",7824 => "10010101",7825 => "01001011",7826 => "11000111",7827 => "00110010",7828 => "00001110",7829 => "10110111",7830 => "10100110",7831 => "10001110",7832 => "10100110",7833 => "01100101",7834 => "01011101",7835 => "10101101",7836 => "01000100",7837 => "10000100",7838 => "00101001",7839 => "10110101",7840 => "00111001",7841 => "11111011",7842 => "10111011",7843 => "11110000",7844 => "00111111",7845 => "00111111",7846 => "01100111",7847 => "01010001",7848 => "01110010",7849 => "00100000",7850 => "00111110",7851 => "01101000",7852 => "10011101",7853 => "10100011",7854 => "11100010",7855 => "11101110",7856 => "11100010",7857 => "00110110",7858 => "11010011",7859 => "11110101",7860 => "01011000",7861 => "01000110",7862 => "11110100",7863 => "10100111",7864 => "10110110",7865 => "10000010",7866 => "01011010",7867 => "00010101",7868 => "11111001",7869 => "00010011",7870 => "10010101",7871 => "01010000",7872 => "01101010",7873 => "11000101",7874 => "11111101",7875 => "10001111",7876 => "10111100",7877 => "10011000",7878 => "10010010",7879 => "00110111",7880 => "10001101",7881 => "00110111",7882 => "00000111",7883 => "11000111",7884 => "01001001",7885 => "11001001",7886 => "00100100",7887 => "10110011",7888 => "11111001",7889 => "00101011",7890 => "11101111",7891 => "10101001",7892 => "00100110",7893 => "10011010",7894 => "10101100",7895 => "01101110",7896 => "01111100",7897 => "01010011",7898 => "10110101",7899 => "10011101",7900 => "11000110",7901 => "01001100",7902 => "00110001",7903 => "11111101",7904 => "00111001",7905 => "11011100",7906 => "10111010",7907 => "10111100",7908 => "10110011",7909 => "00001000",7910 => "00100110",7911 => "01100010",7912 => "01110100",7913 => "01100110",7914 => "00110000",7915 => "01010010",7916 => "00111101",7917 => "01110110",7918 => "00010000",7919 => "10110010",7920 => "01011001",7921 => "11011010",7922 => "10110001",7923 => "01100011",7924 => "01010011",7925 => "01100100",7926 => "11010010",7927 => "01010110",7928 => "11000011",7929 => "00010110",7930 => "10111110",7931 => "01111101",7932 => "01001001",7933 => "01100101",7934 => "11010001",7935 => "01010110",7936 => "00110101",7937 => "11010010",7938 => "01100011",7939 => "10011100",7940 => "11001011",7941 => "00010000",7942 => "00011010",7943 => "11000010",7944 => "00101010",7945 => "11010011",7946 => "00011100",7947 => "01000001",7948 => "00000000",7949 => "11100101",7950 => "01000010",7951 => "01001101",7952 => "01100100",7953 => "00001100",7954 => "00000010",7955 => "10011101",7956 => "11101101",7957 => "11000100",7958 => "00010000",7959 => "00111010",7960 => "00000011",7961 => "11101000",7962 => "01100010",7963 => "00100100",7964 => "10100101",7965 => "10011010",7966 => "10001001",7967 => "11100011",7968 => "11101111",7969 => "01010101",7970 => "00101010",7971 => "01011100",7972 => "10101111",7973 => "00110010",7974 => "00110010",7975 => "00011100",7976 => "11011111",7977 => "00101010",7978 => "10000010",7979 => "11101110",7980 => "01001101",7981 => "00010111",7982 => "00111101",7983 => "00010001",7984 => "00110111",7985 => "10000011",7986 => "01010101",7987 => "10000100",7988 => "00011101",7989 => "11101111",7990 => "01100011",7991 => "00001111",7992 => "11101010",7993 => "11100101",7994 => "01011010",7995 => "00001001",7996 => "01101100",7997 => "10001000",7998 => "11100011",7999 => "01010111",8000 => "10001001",8001 => "01110010",8002 => "01111111",8003 => "10000011",8004 => "10101111",8005 => "01010101",8006 => "10010001",8007 => "11011000",8008 => "10110001",8009 => "00001101",8010 => "00101110",8011 => "00001011",8012 => "11101101",8013 => "11001110",8014 => "10010000",8015 => "11111001",8016 => "11000101",8017 => "10100101",8018 => "10010100",8019 => "11101000",8020 => "01110101",8021 => "11111000",8022 => "01100000",8023 => "11110101",8024 => "01100111",8025 => "00111110",8026 => "10000001",8027 => "01101000",8028 => "11110011",8029 => "11010110",8030 => "01111011",8031 => "01111011",8032 => "00001100",8033 => "01111101",8034 => "01101001",8035 => "11001001",8036 => "10110100",8037 => "10000100",8038 => "11100011",8039 => "01001110",8040 => "01110100",8041 => "00011010",8042 => "11100001",8043 => "10011110",8044 => "00001100",8045 => "01000000",8046 => "10101100",8047 => "00111011",8048 => "11010100",8049 => "10000001",8050 => "11001111",8051 => "10000101",8052 => "10001100",8053 => "00111011",8054 => "11111100",8055 => "11111101",8056 => "10001100",8057 => "10100101",8058 => "11010100",8059 => "00111011",8060 => "11000000",8061 => "01011100",8062 => "01001110",8063 => "01101000",8064 => "00100001",8065 => "11010101",8066 => "01000101",8067 => "01001110",8068 => "01101101",8069 => "10001110",8070 => "01101011",8071 => "11011000",8072 => "10101010",8073 => "10010001",8074 => "00101001",8075 => "01011100",8076 => "01110011",8077 => "10010101",8078 => "00101111",8079 => "01110011",8080 => "10011001",8081 => "01000100",8082 => "10101000",8083 => "01100111",8084 => "00001000",8085 => "10111111",8086 => "10101111",8087 => "11101111",8088 => "11000010",8089 => "01101111",8090 => "00011111",8091 => "01110101",8092 => "11101001",8093 => "10001100",8094 => "10110010",8095 => "00111110",8096 => "10101001",8097 => "01000110",8098 => "10111010",8099 => "01011111",8100 => "11101010",8101 => "01000000",8102 => "01110010",8103 => "11010110",8104 => "10010100",8105 => "10000001",8106 => "11110010",8107 => "00110111",8108 => "01100111",8109 => "01011100",8110 => "01111100",8111 => "00101100",8112 => "00010001",8113 => "11011110",8114 => "10010011",8115 => "01101101",8116 => "10101101",8117 => "11000011",8118 => "10011101",8119 => "01000110",8120 => "11101011",8121 => "00001001",8122 => "10111101",8123 => "11010010",8124 => "00000001",8125 => "11001010",8126 => "00001000",8127 => "11000010",8128 => "01010111",8129 => "10111111",8130 => "10011111",8131 => "01111100",8132 => "00100011",8133 => "10010100",8134 => "11001000",8135 => "00011101",8136 => "01110000",8137 => "10001101",8138 => "10011011",8139 => "00111011",8140 => "00001010",8141 => "10010001",8142 => "00110100",8143 => "01101101",8144 => "10010110",8145 => "01010010",8146 => "00111011",8147 => "01011010",8148 => "01000110",8149 => "10011011",8150 => "01010011",8151 => "00011001",8152 => "11111100",8153 => "01001101",8154 => "00001110",8155 => "01100000",8156 => "00111011",8157 => "00001010",8158 => "11000101",8159 => "11111111",8160 => "01001001",8161 => "11010101",8162 => "10001011",8163 => "10001011",8164 => "11011101",8165 => "00111111",8166 => "01000011",8167 => "00110110",8168 => "10101011",8169 => "11110000",8170 => "00111111",8171 => "11101011",8172 => "01100101",8173 => "11110010",8174 => "01110011",8175 => "00111100",8176 => "01000000",8177 => "01011100",8178 => "10101010",8179 => "10011010",8180 => "10001111",8181 => "01000100",8182 => "01111110",8183 => "11011010",8184 => "00000110",8185 => "11001000",8186 => "01111010",8187 => "01111111",8188 => "01011001",8189 => "00001101",8190 => "10101111",8191 => "01000101",8192 => "10111010",8193 => "00110100",8194 => "10110001",8195 => "01011001",8196 => "01101110",8197 => "00111111",8198 => "10101101",8199 => "00000101",8200 => "01011101",8201 => "11100001",8202 => "00001100",8203 => "11010100",8204 => "10000001",8205 => "11101011",8206 => "00011101",8207 => "00101011",8208 => "10010001",8209 => "01101001",8210 => "11111000",8211 => "11001010",8212 => "10100111",8213 => "10101011",8214 => "01000111",8215 => "11101100",8216 => "01110111",8217 => "10010111",8218 => "00000111",8219 => "00010101",8220 => "10001110",8221 => "00111000",8222 => "01111100",8223 => "00010010",8224 => "00111011",8225 => "01001011",8226 => "11011101",8227 => "00100111",8228 => "10000011",8229 => "01111100",8230 => "11000101",8231 => "10010101",8232 => "01111001",8233 => "11111000",8234 => "11011010",8235 => "01001100",8236 => "01111100",8237 => "01101101",8238 => "01111001",8239 => "01100010",8240 => "01100100",8241 => "00100100",8242 => "01111001",8243 => "11000010",8244 => "00010011",8245 => "11100100",8246 => "10101101",8247 => "10010000",8248 => "01001000",8249 => "10010111",8250 => "10001110",8251 => "10100011",8252 => "11110011",8253 => "10000000",8254 => "10111001",8255 => "00110011",8256 => "11011011",8257 => "01011111",8258 => "01011011",8259 => "00011001",8260 => "01011010",8261 => "00001100",8262 => "01010110",8263 => "00000011",8264 => "00110110",8265 => "11111001",8266 => "00110111",8267 => "11001000",8268 => "01011100",8269 => "11111101",8270 => "00010101",8271 => "01111001",8272 => "11101001",8273 => "01001001",8274 => "11011101",8275 => "10011100",8276 => "10101110",8277 => "11001000",8278 => "10001011",8279 => "10001111",8280 => "00010000",8281 => "00011010",8282 => "01101100",8283 => "11011011",8284 => "01111100",8285 => "11101010",8286 => "01110110",8287 => "11011100",8288 => "00011011",8289 => "11001010",8290 => "10000011",8291 => "10001100",8292 => "11100010",8293 => "01100100",8294 => "01001000",8295 => "10111111",8296 => "11011011",8297 => "11111111",8298 => "11011101",8299 => "11001110",8300 => "11110000",8301 => "00110111",8302 => "10010000",8303 => "01001100",8304 => "00011100",8305 => "01111000",8306 => "11111010",8307 => "10101111",8308 => "00100111",8309 => "00011001",8310 => "01001110",8311 => "01100111",8312 => "10001001",8313 => "01110000",8314 => "01011001",8315 => "11100100",8316 => "10111100",8317 => "00100010",8318 => "11100011",8319 => "00011001",8320 => "01011010",8321 => "01111011",8322 => "11010000",8323 => "11000010",8324 => "01110010",8325 => "01100010",8326 => "10001010",8327 => "11001010",8328 => "00100110",8329 => "00101000",8330 => "00101111",8331 => "11001011",8332 => "10000111",8333 => "00111101",8334 => "00101101",8335 => "00010000",8336 => "00100111",8337 => "00100100",8338 => "01110001",8339 => "10011111",8340 => "10010110",8341 => "01100010",8342 => "01010011",8343 => "01111011",8344 => "01101111",8345 => "00100101",8346 => "10000011",8347 => "11001101",8348 => "00000000",8349 => "01111101",8350 => "00100100",8351 => "10101101",8352 => "10011011",8353 => "01011000",8354 => "00000100",8355 => "01001101",8356 => "00000001",8357 => "11001110",8358 => "10111001",8359 => "11101011",8360 => "01110110",8361 => "00001111",8362 => "00110100",8363 => "00100110",8364 => "10001011",8365 => "10100110",8366 => "10011011",8367 => "10001111",8368 => "10011101",8369 => "01110011",8370 => "00100111",8371 => "00100101",8372 => "01001011",8373 => "10001001",8374 => "00111010",8375 => "01011100",8376 => "10100110",8377 => "01110000",8378 => "11000100",8379 => "00110101",8380 => "11101010",8381 => "11111001",8382 => "11010111",8383 => "11101100",8384 => "10110011",8385 => "10100011",8386 => "10100010",8387 => "01010111",8388 => "11100101",8389 => "10101100",8390 => "01100000",8391 => "10010000",8392 => "00011101",8393 => "11010000",8394 => "11000101",8395 => "00100000",8396 => "00110001",8397 => "00100010",8398 => "00111100",8399 => "10111010",8400 => "01010001",8401 => "01011001",8402 => "10000101",8403 => "10100111",8404 => "10110111",8405 => "01100111",8406 => "00101010",8407 => "01001110",8408 => "01010001",8409 => "00001111",8410 => "01001111",8411 => "10100001",8412 => "00110010",8413 => "11100101",8414 => "10100000",8415 => "00100010",8416 => "11010101",8417 => "01011110",8418 => "11100110",8419 => "00111001",8420 => "00110100",8421 => "00011000",8422 => "10010101",8423 => "10100110",8424 => "00001010",8425 => "00100010",8426 => "00101000",8427 => "10011100",8428 => "10010011",8429 => "01011110",8430 => "00001000",8431 => "01011101",8432 => "00111001",8433 => "11110100",8434 => "11001110",8435 => "11111101",8436 => "01101000",8437 => "11111010",8438 => "10110110",8439 => "01111110",8440 => "00000000",8441 => "11100001",8442 => "10001011",8443 => "00100110",8444 => "01000101",8445 => "10001110",8446 => "01011000",8447 => "11011001",8448 => "11100001",8449 => "00111010",8450 => "01100101",8451 => "10000101",8452 => "00010000",8453 => "11010011",8454 => "10001011",8455 => "01011111",8456 => "10110001",8457 => "11111100",8458 => "00000111",8459 => "01010101",8460 => "10010111",8461 => "11100110",8462 => "11101000",8463 => "10000101",8464 => "11010000",8465 => "11101001",8466 => "11101011",8467 => "00010011",8468 => "11100011",8469 => "00111001",8470 => "00100101",8471 => "10100111",8472 => "01011111",8473 => "11110011",8474 => "10100001",8475 => "01011111",8476 => "11010001",8477 => "10110100",8478 => "10000101",8479 => "11101101",8480 => "01000001",8481 => "11010000",8482 => "01101010",8483 => "00010110",8484 => "10101111",8485 => "01101010",8486 => "11011010",8487 => "00111101",8488 => "01111001",8489 => "10010111",8490 => "10010001",8491 => "00001010",8492 => "11101111",8493 => "10100000",8494 => "00011000",8495 => "10100101",8496 => "01001011",8497 => "00100010",8498 => "00011110",8499 => "10111100",8500 => "10100000",8501 => "00101000",8502 => "11001101",8503 => "10000010",8504 => "00010110",8505 => "00110100",8506 => "01001000",8507 => "11001101",8508 => "01101101",8509 => "11100101",8510 => "10100110",8511 => "10101110",8512 => "01100010",8513 => "10111100",8514 => "01000110",8515 => "00000100",8516 => "00111100",8517 => "10000110",8518 => "01101001",8519 => "10001100",8520 => "10001101",8521 => "00001000",8522 => "01101010",8523 => "11110111",8524 => "10010100",8525 => "00101110",8526 => "01100101",8527 => "01100101",8528 => "11100000",8529 => "11111101",8530 => "10000110",8531 => "00101110",8532 => "10100011",8533 => "00010100",8534 => "10101110",8535 => "10011101",8536 => "00100100",8537 => "01011000",8538 => "00010100",8539 => "00011001",8540 => "11000101",8541 => "00111111",8542 => "11101111",8543 => "01110010",8544 => "01001011",8545 => "10011111",8546 => "10100111",8547 => "10010100",8548 => "11111101",8549 => "01001011",8550 => "10011010",8551 => "01010011",8552 => "10010111",8553 => "00001000",8554 => "01010011",8555 => "11110101",8556 => "11001011",8557 => "10101110",8558 => "10110011",8559 => "01010100",8560 => "00111110",8561 => "11011001",8562 => "11110011",8563 => "01100110",8564 => "01110000",8565 => "10111101",8566 => "11011000",8567 => "00111010",8568 => "10011001",8569 => "11100000",8570 => "10111100",8571 => "10011111",8572 => "01101110",8573 => "10111100",8574 => "11100100",8575 => "01101110",8576 => "11001001",8577 => "00101001",8578 => "01101110",8579 => "11010110",8580 => "10100101",8581 => "01111010",8582 => "11001000",8583 => "00001110",8584 => "01010101",8585 => "00110100",8586 => "11011000",8587 => "10110011",8588 => "11011001",8589 => "01110100",8590 => "11010101",8591 => "10000001",8592 => "10010110",8593 => "01111010",8594 => "10100001",8595 => "11101101",8596 => "00101010",8597 => "01010101",8598 => "00001111",8599 => "01011000",8600 => "10100010",8601 => "00001010",8602 => "10101001",8603 => "01101101",8604 => "00110011",8605 => "10000001",8606 => "01001101",8607 => "01100011",8608 => "11111010",8609 => "01111011",8610 => "01101101",8611 => "00100000",8612 => "10010111",8613 => "00011001",8614 => "01011011",8615 => "11010001",8616 => "00100000",8617 => "00011011",8618 => "11101101",8619 => "01101001",8620 => "00001001",8621 => "11000011",8622 => "11100000",8623 => "10001101",8624 => "10010111",8625 => "10101000",8626 => "10110100",8627 => "10100000",8628 => "10001111",8629 => "00100101",8630 => "10000111",8631 => "11011011",8632 => "01101100",8633 => "10011000",8634 => "10001000",8635 => "11010101",8636 => "11100111",8637 => "11001010",8638 => "11011110",8639 => "11101101",8640 => "00011110",8641 => "01111011",8642 => "01000101",8643 => "00110001",8644 => "11010100",8645 => "01010011",8646 => "11110010",8647 => "10101010",8648 => "11100110",8649 => "01011101",8650 => "00101011",8651 => "11010000",8652 => "00010101",8653 => "01000000",8654 => "01100000",8655 => "10010100",8656 => "00010000",8657 => "11011110",8658 => "00001001",8659 => "01100001",8660 => "10010011",8661 => "00000111",8662 => "01110100",8663 => "11101111",8664 => "10101000",8665 => "00100000",8666 => "11101010",8667 => "01100001",8668 => "01110011",8669 => "00101001",8670 => "11100010",8671 => "01110100",8672 => "01111101",8673 => "01000011",8674 => "01101011",8675 => "00000011",8676 => "10011101",8677 => "01110011",8678 => "11010011",8679 => "01100100",8680 => "00001011",8681 => "01011111",8682 => "10000000",8683 => "11000010",8684 => "01000100",8685 => "01000100",8686 => "01110001",8687 => "11001010",8688 => "00110111",8689 => "00011100",8690 => "11111111",8691 => "01101000",8692 => "11111110",8693 => "11110110",8694 => "01100000",8695 => "01010111",8696 => "01010000",8697 => "10101010",8698 => "11010101",8699 => "00010001",8700 => "10010111",8701 => "10000010",8702 => "01110110",8703 => "00000100",8704 => "11000100",8705 => "00001010",8706 => "01000001",8707 => "00101100",8708 => "01110111",8709 => "00001001",8710 => "10011101",8711 => "10110001",8712 => "11100011",8713 => "01010110",8714 => "11010111",8715 => "11011110",8716 => "11110101",8717 => "10100010",8718 => "10011000",8719 => "10001111",8720 => "00110000",8721 => "11001011",8722 => "10100011",8723 => "10011101",8724 => "11110000",8725 => "01001100",8726 => "01110111",8727 => "10110101",8728 => "01110110",8729 => "11011110",8730 => "11100001",8731 => "00010110",8732 => "11001011",8733 => "00110000",8734 => "10100010",8735 => "00101011",8736 => "00100000",8737 => "10000000",8738 => "11011101",8739 => "01100001",8740 => "00111000",8741 => "11110100",8742 => "00111011",8743 => "11011010",8744 => "01111011",8745 => "10111011",8746 => "00010001",8747 => "11100110",8748 => "00010000",8749 => "01011001",8750 => "00110111",8751 => "01000001",8752 => "10011110",8753 => "10011010",8754 => "01111011",8755 => "10001110",8756 => "01000000",8757 => "01111101",8758 => "01100011",8759 => "01010001",8760 => "01011110",8761 => "10010110",8762 => "00100011",8763 => "10100000",8764 => "11110000",8765 => "11100010",8766 => "11111010",8767 => "01011101",8768 => "00100001",8769 => "01110000",8770 => "00000011",8771 => "01100111",8772 => "10011000",8773 => "00000101",8774 => "01111110",8775 => "00011010",8776 => "11000011",8777 => "10011001",8778 => "11100101",8779 => "10011100",8780 => "00111000",8781 => "10010011",8782 => "11110011",8783 => "01010010",8784 => "01010111",8785 => "01011111",8786 => "11000011",8787 => "00000011",8788 => "11000001",8789 => "11010110",8790 => "01101000",8791 => "01011001",8792 => "01110011",8793 => "01010101",8794 => "00101111",8795 => "10110101",8796 => "10101001",8797 => "01001100",8798 => "01011010",8799 => "01011011",8800 => "01010110",8801 => "10110101",8802 => "10111101",8803 => "10110111",8804 => "11010001",8805 => "00101000",8806 => "00001100",8807 => "00100100",8808 => "00011111",8809 => "01011100",8810 => "00011100",8811 => "10101010",8812 => "00011110",8813 => "10100110",8814 => "10101000",8815 => "11011011",8816 => "00111011",8817 => "00111101",8818 => "01010110",8819 => "11110110",8820 => "01110001",8821 => "10101010",8822 => "11011001",8823 => "11001101",8824 => "00011010",8825 => "10110000",8826 => "10101000",8827 => "01101011",8828 => "11000011",8829 => "10100010",8830 => "00110111",8831 => "01101110",8832 => "00011011",8833 => "00100111",8834 => "11001110",8835 => "11010111",8836 => "01010010",8837 => "11000010",8838 => "10010000",8839 => "11111110",8840 => "00111010",8841 => "00101111",8842 => "11011000",8843 => "00101000",8844 => "01001011",8845 => "01111111",8846 => "01001110",8847 => "00100010",8848 => "00111001",8849 => "11101111",8850 => "01101010",8851 => "11011000",8852 => "11101100",8853 => "01010000",8854 => "01110011",8855 => "10110101",8856 => "00101111",8857 => "01101010",8858 => "11000010",8859 => "01101111",8860 => "00000010",8861 => "11010011",8862 => "10110111",8863 => "00111100",8864 => "11100101",8865 => "00100110",8866 => "10000010",8867 => "01111101",8868 => "00111100",8869 => "11110110",8870 => "11001010",8871 => "01111000",8872 => "11101000",8873 => "11001011",8874 => "11001110",8875 => "01010110",8876 => "01011010",8877 => "10101011",8878 => "01111110",8879 => "01111111",8880 => "00011000",8881 => "11001010",8882 => "01111001",8883 => "11000001",8884 => "11010111",8885 => "10110100",8886 => "11111000",8887 => "10010110",8888 => "10111100",8889 => "10001100",8890 => "01010000",8891 => "01011101",8892 => "01000011",8893 => "10111100",8894 => "00000101",8895 => "11101111",8896 => "10110100",8897 => "10101110",8898 => "01110100",8899 => "01001011",8900 => "10100111",8901 => "00001011",8902 => "11111000",8903 => "01010110",8904 => "00100011",8905 => "00011100",8906 => "01110000",8907 => "01101100",8908 => "00101111",8909 => "11110010",8910 => "00110111",8911 => "10100111",8912 => "11001011",8913 => "11110011",8914 => "01010111",8915 => "00001111",8916 => "00110100",8917 => "00000110",8918 => "10011111",8919 => "00100100",8920 => "10010010",8921 => "11100110",8922 => "01010110",8923 => "11010110",8924 => "11000000",8925 => "11100000",8926 => "11000101",8927 => "00001101",8928 => "10110101",8929 => "00001101",8930 => "11100110",8931 => "01110100",8932 => "01101100",8933 => "00110000",8934 => "00100111",8935 => "10111001",8936 => "00011010",8937 => "11011001",8938 => "10101111",8939 => "11001010",8940 => "01010110",8941 => "01111101",8942 => "10011111",8943 => "01110101",8944 => "00111000",8945 => "01011110",8946 => "00011001",8947 => "01001111",8948 => "10100111",8949 => "01010100",8950 => "01101100",8951 => "00111110",8952 => "01101000",8953 => "00110101",8954 => "10110000",8955 => "10011111",8956 => "11110111",8957 => "01101101",8958 => "01101101",8959 => "01011001",8960 => "11100100",8961 => "11010111",8962 => "00110001",8963 => "10110011",8964 => "01010111",8965 => "01100111",8966 => "01100101",8967 => "10100010",8968 => "11100000",8969 => "11011101",8970 => "01000001",8971 => "11010001",8972 => "11001001",8973 => "10110111",8974 => "10000111",8975 => "11000111",8976 => "11110000",8977 => "00111100",8978 => "01111001",8979 => "11001010",8980 => "10001100",8981 => "11001110",8982 => "01000010",8983 => "11011101",8984 => "00100100",8985 => "01011101",8986 => "00010011",8987 => "00110111",8988 => "10110111",8989 => "11001111",8990 => "01111000",8991 => "11001000",8992 => "10100110",8993 => "01100000",8994 => "11010001",8995 => "11101110",8996 => "11011111",8997 => "00011010",8998 => "01101100",8999 => "10111001",9000 => "11011001",9001 => "10101111",9002 => "00011111",9003 => "11010011",9004 => "10000010",9005 => "10001101",9006 => "11010101",9007 => "11010000",9008 => "00000101",9009 => "10101111",9010 => "00000011",9011 => "11000010",9012 => "01011111",9013 => "11010100",9014 => "11000001",9015 => "10100101",9016 => "01111001",9017 => "01000110",9018 => "10100100",9019 => "11000011",9020 => "10111011",9021 => "11111110",9022 => "11001000",9023 => "01011101",9024 => "01111010",9025 => "01000011",9026 => "11110101",9027 => "01001010",9028 => "00101101",9029 => "01101000",9030 => "01100010",9031 => "11101000",9032 => "11100110",9033 => "00000100",9034 => "11100100",9035 => "10101101",9036 => "01101101",9037 => "10011010",9038 => "01101001",9039 => "00111010",9040 => "00001101",9041 => "00010100",9042 => "10010110",9043 => "10001100",9044 => "11101000",9045 => "01111011",9046 => "10001101",9047 => "01110110",9048 => "10000100",9049 => "00011101",9050 => "00011111",9051 => "01101001",9052 => "01100101",9053 => "00010101",9054 => "01110011",9055 => "01001001",9056 => "01100111",9057 => "11010101",9058 => "00000000",9059 => "11110101",9060 => "11101100",9061 => "00100110",9062 => "00100101",9063 => "00010110",9064 => "11011000",9065 => "11111101",9066 => "10111101",9067 => "01001111",9068 => "11011111",9069 => "00000011",9070 => "01111001",9071 => "11101001",9072 => "01110001",9073 => "01001001",9074 => "11011100",9075 => "01011100",9076 => "01000111",9077 => "11100110",9078 => "10110110",9079 => "11111100",9080 => "11011110",9081 => "00100000",9082 => "01101011",9083 => "00101111",9084 => "10011010",9085 => "11111010",9086 => "11110010",9087 => "01110001",9088 => "11000100",9089 => "01111000",9090 => "10101000",9091 => "11000011",9092 => "00111011",9093 => "01111100",9094 => "11011110",9095 => "11110001",9096 => "10110011",9097 => "11111010",9098 => "10011001",9099 => "11111001",9100 => "01111010",9101 => "10001010",9102 => "10001100",9103 => "00110001",9104 => "11101011",9105 => "00011011",9106 => "11011001",9107 => "01100001",9108 => "00101000",9109 => "00010111",9110 => "10000001",9111 => "11101011",9112 => "00110110",9113 => "01111101",9114 => "01011101",9115 => "01110101",9116 => "11000111",9117 => "00100011",9118 => "00000001",9119 => "10111010",9120 => "10000101",9121 => "11110001",9122 => "00101110",9123 => "00000000",9124 => "01011001",9125 => "11011011",9126 => "10101110",9127 => "01000011",9128 => "10101100",9129 => "10101101",9130 => "11101000",9131 => "11101101",9132 => "00101001",9133 => "10110111",9134 => "00101100",9135 => "01001000",9136 => "00010110",9137 => "10111001",9138 => "10101111",9139 => "01110100",9140 => "00011010",9141 => "00110001",9142 => "00100111",9143 => "10001111",9144 => "01010000",9145 => "01000100",9146 => "01000111",9147 => "01100010",9148 => "11001010",9149 => "01111100",9150 => "11001101",9151 => "01111110",9152 => "11110011",9153 => "01000101",9154 => "10001101",9155 => "11101011",9156 => "00000010",9157 => "10100000",9158 => "00111110",9159 => "01011100",9160 => "10100100",9161 => "10100101",9162 => "11110110",9163 => "01110111",9164 => "11001001",9165 => "11100111",9166 => "10111011",9167 => "01010100",9168 => "10111001",9169 => "11100100",9170 => "11101101",9171 => "10011010",9172 => "00110001",9173 => "10011111",9174 => "01111010",9175 => "00000100",9176 => "10100110",9177 => "00011101",9178 => "10011100",9179 => "00011111",9180 => "01010001",9181 => "10001110",9182 => "11101001",9183 => "11100101",9184 => "01101101",9185 => "10010000",9186 => "01011110",9187 => "01011111",9188 => "00100001",9189 => "00000100",9190 => "11110111",9191 => "01101001",9192 => "00100110",9193 => "01111010",9194 => "00101011",9195 => "10111010",9196 => "10111100",9197 => "01000011",9198 => "00111011",9199 => "01000011",9200 => "10101000",9201 => "10010111",9202 => "00010111",9203 => "01111010",9204 => "01011011",9205 => "01010010",9206 => "11000100",9207 => "11010000",9208 => "01001000",9209 => "11101110",9210 => "11101100",9211 => "00000000",9212 => "11001000",9213 => "11000000",9214 => "00001101",9215 => "11101010",9216 => "10101010",9217 => "11000000",9218 => "10000001",9219 => "11001100",9220 => "00010000",9221 => "11111001",9222 => "11011001",9223 => "11111110",9224 => "10101101",9225 => "00111010",9226 => "10000110",9227 => "10101111",9228 => "01001101",9229 => "01100101",9230 => "00001011",9231 => "11101111",9232 => "11000100",9233 => "01010011",9234 => "01101000",9235 => "10010110",9236 => "01010011",9237 => "01111000",9238 => "11110111",9239 => "10100110",9240 => "00111010",9241 => "00010111",9242 => "01001011",9243 => "11011011",9244 => "11100011",9245 => "00110100",9246 => "00100110",9247 => "11011010",9248 => "01011010",9249 => "00011010",9250 => "10001000",9251 => "10100000",9252 => "00010001",9253 => "00010111",9254 => "01100010",9255 => "11110001",9256 => "00101110",9257 => "11000101",9258 => "00101110",9259 => "00110110",9260 => "11000101",9261 => "01011000",9262 => "11110110",9263 => "10011000",9264 => "00111111",9265 => "01001101",9266 => "01110000",9267 => "10010100",9268 => "10100000",9269 => "11010110",9270 => "10011000",9271 => "00101101",9272 => "10100011",9273 => "10001111",9274 => "11110111",9275 => "10110010",9276 => "00000000",9277 => "00100100",9278 => "10110001",9279 => "11011010",9280 => "00011110",9281 => "10011101",9282 => "11011101",9283 => "00101011",9284 => "01001011",9285 => "11000001",9286 => "10000111",9287 => "00001000",9288 => "01100111",9289 => "00110110",9290 => "01001011",9291 => "00010001",9292 => "00111001",9293 => "01101010",9294 => "00010010",9295 => "01110000",9296 => "10101000",9297 => "01001010",9298 => "10110101",9299 => "10010100",9300 => "11100110",9301 => "01011110",9302 => "01111000",9303 => "10011000",9304 => "10000001",9305 => "01000000",9306 => "01000101",9307 => "00110010",9308 => "11100101",9309 => "00111011",9310 => "10110110",9311 => "01110111",9312 => "10011100",9313 => "10000001",9314 => "00001010",9315 => "10110001",9316 => "01111101",9317 => "10001101",9318 => "00000010",9319 => "00101000",9320 => "10001101",9321 => "00000011",9322 => "00010110",9323 => "00111110",9324 => "10011011",9325 => "10110001",9326 => "10000100",9327 => "11001010",9328 => "10001101",9329 => "11000000",9330 => "10001011",9331 => "11110010",9332 => "01111010",9333 => "10110100",9334 => "01110111",9335 => "11101011",9336 => "11000001",9337 => "10101001",9338 => "11101110",9339 => "11001010",9340 => "00011101",9341 => "01101001",9342 => "00010101",9343 => "11001000",9344 => "00100011",9345 => "10110011",9346 => "01111001",9347 => "01000101",9348 => "11101100",9349 => "11110111",9350 => "01010001",9351 => "01010111",9352 => "10111111",9353 => "11101100",9354 => "00101100",9355 => "10011001",9356 => "11001101",9357 => "11100000",9358 => "01011111",9359 => "11011110",9360 => "10001111",9361 => "11100011",9362 => "11010101",9363 => "10110001",9364 => "01111011",9365 => "00001100",9366 => "10101001",9367 => "10100110",9368 => "00100011",9369 => "11001100",9370 => "11011100",9371 => "01110110",9372 => "00010000",9373 => "00110110",9374 => "11000111",9375 => "10011111",9376 => "00111011",9377 => "11101110",9378 => "00011001",9379 => "00110111",9380 => "10110000",9381 => "10110001",9382 => "00111010",9383 => "10000100",9384 => "00110000",9385 => "01001111",9386 => "01001100",9387 => "00010011",9388 => "11100011",9389 => "11001100",9390 => "01000000",9391 => "01101101",9392 => "00100001",9393 => "01100010",9394 => "10111000",9395 => "11000100",9396 => "11010000",9397 => "11011111",9398 => "10101011",9399 => "00101000",9400 => "00111011",9401 => "00011110",9402 => "10101110",9403 => "11011110",9404 => "11100110",9405 => "10110101",9406 => "11010111",9407 => "00110011",9408 => "10111011",9409 => "11000000",9410 => "01110011",9411 => "10010100",9412 => "10101100",9413 => "00001000",9414 => "11011010",9415 => "00011100",9416 => "10101001",9417 => "01100110",9418 => "11101101",9419 => "01000001",9420 => "01101010",9421 => "01101000",9422 => "00110010",9423 => "11111101",9424 => "01000011",9425 => "00010011",9426 => "01101010",9427 => "11100110",9428 => "11000100",9429 => "10010101",9430 => "00001011",9431 => "11001101",9432 => "01101011",9433 => "11111011",9434 => "00000100",9435 => "01011100",9436 => "00101010",9437 => "00111000",9438 => "00011000",9439 => "00001101",9440 => "11010100",9441 => "01110101",9442 => "00100010",9443 => "00110111",9444 => "01101101",9445 => "00010011",9446 => "01011000",9447 => "10101110",9448 => "10001111",9449 => "11010010",9450 => "00011100",9451 => "01101000",9452 => "10100100",9453 => "00101100",9454 => "00001011",9455 => "01100110",9456 => "11101001",9457 => "11010010",9458 => "10110010",9459 => "01101001",9460 => "10001011",9461 => "11111110",9462 => "01010110",9463 => "01101110",9464 => "00000001",9465 => "01100100",9466 => "01001000",9467 => "01110011",9468 => "01001111",9469 => "10011101",9470 => "11111010",9471 => "10101001",9472 => "01011011",9473 => "11000000",9474 => "01001100",9475 => "00011001",9476 => "10111111",9477 => "00000010",9478 => "11101010",9479 => "10111110",9480 => "01110110",9481 => "11010000",9482 => "00011100",9483 => "01101100",9484 => "11111010",9485 => "10000001",9486 => "00001101",9487 => "00011111",9488 => "00110111",9489 => "00001000",9490 => "00101101",9491 => "00101101",9492 => "00010110",9493 => "10101001",9494 => "11101010",9495 => "11111011",9496 => "10001101",9497 => "00111110",9498 => "01000101",9499 => "01011011",9500 => "00010100",9501 => "11110110",9502 => "11110010",9503 => "00111011",9504 => "11001101",9505 => "11110011",9506 => "01000010",9507 => "01111001",9508 => "01100001",9509 => "01000001",9510 => "01111000",9511 => "11000000",9512 => "01110111",9513 => "11000001",9514 => "11011100",9515 => "01000010",9516 => "00110100",9517 => "10001001",9518 => "01110111",9519 => "10100000",9520 => "01101011",9521 => "10101111",9522 => "10100110",9523 => "00001011",9524 => "10011100",9525 => "01101111",9526 => "11100001",9527 => "11101111",9528 => "10101111",9529 => "10011100",9530 => "10011011",9531 => "10000001",9532 => "10010110",9533 => "00110000",9534 => "11010000",9535 => "00101000",9536 => "01000110",9537 => "01110100",9538 => "10010011",9539 => "10010011",9540 => "10111110",9541 => "01011111",9542 => "01000011",9543 => "11001101",9544 => "10011000",9545 => "10101110",9546 => "01101101",9547 => "01001111",9548 => "11100010",9549 => "00100011",9550 => "00111011",9551 => "11100101",9552 => "01011111",9553 => "11110111",9554 => "00011110",9555 => "01110100",9556 => "10001010",9557 => "11011001",9558 => "11001001",9559 => "10000011",9560 => "11100101",9561 => "10010001",9562 => "10111010",9563 => "11100010",9564 => "01111111",9565 => "01010001",9566 => "11011110",9567 => "00110110",9568 => "00111110",9569 => "00000101",9570 => "11010110",9571 => "11110110",9572 => "00111111",9573 => "11001000",9574 => "11011000",9575 => "10111100",9576 => "01100101",9577 => "01010011",9578 => "01000011",9579 => "11110001",9580 => "00101101",9581 => "00011100",9582 => "11010011",9583 => "01110100",9584 => "01010101",9585 => "11011110",9586 => "01100110",9587 => "11110101",9588 => "10010111",9589 => "01011001",9590 => "00000111",9591 => "11101000",9592 => "01010000",9593 => "01110011",9594 => "10010010",9595 => "00110010",9596 => "01011110",9597 => "11100100",9598 => "01001011",9599 => "00000011",9600 => "10100001",9601 => "01001111",9602 => "11111111",9603 => "10011000",9604 => "00011000",9605 => "11010000",9606 => "10100001",9607 => "11110010",9608 => "11000001",9609 => "10011111",9610 => "11011100",9611 => "11010011",9612 => "01000011",9613 => "00011101",9614 => "00100110",9615 => "11100010",9616 => "11001010",9617 => "11010010",9618 => "01100010",9619 => "01111111",9620 => "10101001",9621 => "00111101",9622 => "01001100",9623 => "10111001",9624 => "10010100",9625 => "10110001",9626 => "10010000",9627 => "00101001",9628 => "00110000",9629 => "10111011",9630 => "00001111",9631 => "10010000",9632 => "01010011",9633 => "01010110",9634 => "10001101",9635 => "11000100",9636 => "10110001",9637 => "01010001",9638 => "11000110",9639 => "10101001",9640 => "10100101",9641 => "00101100",9642 => "11100000",9643 => "11010001",9644 => "11111000",9645 => "11101010",9646 => "10100000",9647 => "01001110",9648 => "00011001",9649 => "10010010",9650 => "10101111",9651 => "00010111",9652 => "10101011",9653 => "11010011",9654 => "01101110",9655 => "00100110",9656 => "11010000",9657 => "10010101",9658 => "10101011",9659 => "01100110",9660 => "00011011",9661 => "11001111",9662 => "01110101",9663 => "10101010",9664 => "01100010",9665 => "01100001",9666 => "10111110",9667 => "00101001",9668 => "00101101",9669 => "10100000",9670 => "00110011",9671 => "10000001",9672 => "01011010",9673 => "10111101",9674 => "11100011",9675 => "00010110",9676 => "01000001",9677 => "11010000",9678 => "00110010",9679 => "10110001",9680 => "10010011",9681 => "01000101",9682 => "11101001",9683 => "10001101",9684 => "10011010",9685 => "01100111",9686 => "00010010",9687 => "01010000",9688 => "10110001",9689 => "11111101",9690 => "10101011",9691 => "00110100",9692 => "11010001",9693 => "01111100",9694 => "11000011",9695 => "01100011",9696 => "10010001",9697 => "11010101",9698 => "10110010",9699 => "01010110",9700 => "11100011",9701 => "10010011",9702 => "00110010",9703 => "11101100",9704 => "11010001",9705 => "01001010",9706 => "11011010",9707 => "01010010",9708 => "00110110",9709 => "00110111",9710 => "11101001",9711 => "10010110",9712 => "01010010",9713 => "01000001",9714 => "11110010",9715 => "11011011",9716 => "00010001",9717 => "11000111",9718 => "11111000",9719 => "01011011",9720 => "01111110",9721 => "11101111",9722 => "10110011",9723 => "01100101",9724 => "11010011",9725 => "01011011",9726 => "01111100",9727 => "00111111",9728 => "11011110",9729 => "11001111",9730 => "00100010",9731 => "00100111",9732 => "11110101",9733 => "00000001",9734 => "10000111",9735 => "10111100",9736 => "10111101",9737 => "10110011",9738 => "01001101",9739 => "10011110",9740 => "01110101",9741 => "01101001",9742 => "10010000",9743 => "00110001",9744 => "10101111",9745 => "10101010",9746 => "11000100",9747 => "11101000",9748 => "01100110",9749 => "10101100",9750 => "01010101",9751 => "10101110",9752 => "01011101",9753 => "01011100",9754 => "00110000",9755 => "01111111",9756 => "11100110",9757 => "00011111",9758 => "01101101",9759 => "01011010",9760 => "01000011",9761 => "00101010",9762 => "10001101",9763 => "10110000",9764 => "10011000",9765 => "01000111",9766 => "11001101",9767 => "01111000",9768 => "01100111",9769 => "01100100",9770 => "00010110",9771 => "01100110",9772 => "10000010",9773 => "01000010",9774 => "00000010",9775 => "10001000",9776 => "10110001",9777 => "01000100",9778 => "11000010",9779 => "00010011",9780 => "01101000",9781 => "10111111",9782 => "11001010",9783 => "10100100",9784 => "10110001",9785 => "10011000",9786 => "01011101",9787 => "00101111",9788 => "11101110",9789 => "10111001",9790 => "11010100",9791 => "10111011",9792 => "11110111",9793 => "10110000",9794 => "11110001",9795 => "11100100",9796 => "00111000",9797 => "00111001",9798 => "10100110",9799 => "01000011",9800 => "11011100",9801 => "11111100",9802 => "10001010",9803 => "00001100",9804 => "10011101",9805 => "00001001",9806 => "10111100",9807 => "11001001",9808 => "10010110",9809 => "10110101",9810 => "11100110",9811 => "11111011",9812 => "11100111",9813 => "10000000",9814 => "10000111",9815 => "11110001",9816 => "10010110",9817 => "11011011",9818 => "10111010",9819 => "00101101",9820 => "11111101",9821 => "10000001",9822 => "00001100",9823 => "01010110",9824 => "00001111",9825 => "00110000",9826 => "00001011",9827 => "10011111",9828 => "00101010",9829 => "00011001",9830 => "10001110",9831 => "00101010",9832 => "11101010",9833 => "11011001",9834 => "00011100",9835 => "01100111",9836 => "11110010",9837 => "00010010",9838 => "10010111",9839 => "10110111",9840 => "11011010",9841 => "11000011",9842 => "10101101",9843 => "11011011",9844 => "00011001",9845 => "00010101",9846 => "01001000",9847 => "01101111",9848 => "01111010",9849 => "10010110",9850 => "01011011",9851 => "01101111",9852 => "10100111",9853 => "11101101",9854 => "00100000",9855 => "01010111",9856 => "10110001",9857 => "00111111",9858 => "11100000",9859 => "10111000",9860 => "10100001",9861 => "11000110",9862 => "11110001",9863 => "11011000",9864 => "00001110",9865 => "10100010",9866 => "01100110",9867 => "11010101",9868 => "10100100",9869 => "01111011",9870 => "10010001",9871 => "10111100",9872 => "01100011",9873 => "11010111",9874 => "01100101",9875 => "11001011",9876 => "11100010",9877 => "10101000",9878 => "11001000",9879 => "11000100",9880 => "10001100",9881 => "10111001",9882 => "10011101",9883 => "10101001",9884 => "10111111",9885 => "10010110",9886 => "01001010",9887 => "00001010",9888 => "10101101",9889 => "11110111",9890 => "00011110",9891 => "01110111",9892 => "11100111",9893 => "01000011",9894 => "11001101",9895 => "01011001",9896 => "10010010",9897 => "10001110",9898 => "00010101",9899 => "10101000",9900 => "01011101",9901 => "10000001",9902 => "11010111",9903 => "10100000",9904 => "11111000",9905 => "10011110",9906 => "11101101",9907 => "01110011",9908 => "11110111",9909 => "01110000",9910 => "01110000",9911 => "00100100",9912 => "00000111",9913 => "10100000",9914 => "11011111",9915 => "01011111",9916 => "00011010",9917 => "11111111",9918 => "11100010",9919 => "00100000",9920 => "10111110",9921 => "00100010",9922 => "00101000",9923 => "00111000",9924 => "00110110",9925 => "11011100",9926 => "11001001",9927 => "10111101",9928 => "11011101",9929 => "10000101",9930 => "10110100",9931 => "00110000",9932 => "10101011",9933 => "10001101",9934 => "11010011",9935 => "11000101",9936 => "10011001",9937 => "00111110",9938 => "00110111",9939 => "10100000",9940 => "11011101",9941 => "00111110",9942 => "11000000",9943 => "00001001",9944 => "11100110",9945 => "10101000",9946 => "10101000",9947 => "00010111",9948 => "00001111",9949 => "10110110",9950 => "00111101",9951 => "00111000",9952 => "00100110",9953 => "10110000",9954 => "10110110",9955 => "10110111",9956 => "00011000",9957 => "00011110",9958 => "10001010",9959 => "00001111",9960 => "10010110",9961 => "11000111",9962 => "10111000",9963 => "10001010",9964 => "01111000",9965 => "00110000",9966 => "00110111",9967 => "11010111",9968 => "00100101",9969 => "10000001",9970 => "10111111",9971 => "10010001",9972 => "00011101",9973 => "10000011",9974 => "10111110",9975 => "01010100",9976 => "11111000",9977 => "00001110",9978 => "00011000",9979 => "10011000",9980 => "11010010",9981 => "01101100",9982 => "10011111",9983 => "10000111",9984 => "10100111",9985 => "01011101",9986 => "01100100",9987 => "10100001",9988 => "11111100",9989 => "10010001",9990 => "10100000",9991 => "10101100",9992 => "11111100",9993 => "00111011",9994 => "01010110",9995 => "01010100",9996 => "11001010",9997 => "01010111",9998 => "01000110",9999 => "01111111",10000 => "11100101",10001 => "01010011",10002 => "11111010",10003 => "10101100",10004 => "01010000",10005 => "10010011",10006 => "11111110",10007 => "10110011",10008 => "01111001",10009 => "10110111",10010 => "00010100",10011 => "11010110",10012 => "00100010",10013 => "00111100",10014 => "01110001",10015 => "10010111",10016 => "01101110",10017 => "10000101",10018 => "01001101",10019 => "01000111",10020 => "01010011",10021 => "11000000",10022 => "01011110",10023 => "10010101",10024 => "01001000",10025 => "10100110",10026 => "11001001",10027 => "10100100",10028 => "11110100",10029 => "10001100",10030 => "11100111",10031 => "01011100",10032 => "10101100",10033 => "01101000",10034 => "00010001",10035 => "10100101",10036 => "11001010",10037 => "00001010",10038 => "11011001",10039 => "00110010",10040 => "10110101",10041 => "11010011",10042 => "11110110",10043 => "01110100",10044 => "10000001",10045 => "10000000",10046 => "01010001",10047 => "00001101",10048 => "10010010",10049 => "00111100",10050 => "11111110",10051 => "11000010",10052 => "01011110",10053 => "11111111",10054 => "10011010",10055 => "01100110",10056 => "11001101",10057 => "10111111",10058 => "01110111",10059 => "00101011",10060 => "11111001",10061 => "10011100",10062 => "11110010",10063 => "01010011",10064 => "00000000",10065 => "01001000",10066 => "00101000",10067 => "10111001",10068 => "01010011",10069 => "11001001",10070 => "01101101",10071 => "01100001",10072 => "01010110",10073 => "11111011",10074 => "01111100",10075 => "11010100",10076 => "00110111",10077 => "01101001",10078 => "01111100",10079 => "01000100",10080 => "00011000",10081 => "00111001",10082 => "11110010",10083 => "10000111",10084 => "10000101",10085 => "11010000",10086 => "10011001",10087 => "11010011",10088 => "01100010",10089 => "00001101",10090 => "11000100",10091 => "00011100",10092 => "11110100",10093 => "01001011",10094 => "01101011",10095 => "01111000",10096 => "00111100",10097 => "10000101",10098 => "01010001",10099 => "11111010",10100 => "10101101",10101 => "00000010",10102 => "11001111",10103 => "10010100",10104 => "01111010",10105 => "00000110",10106 => "10110000",10107 => "10111110",10108 => "10110011",10109 => "00110011",10110 => "10011101",10111 => "10101011",10112 => "11111110",10113 => "01010011",10114 => "00001011",10115 => "11111101",10116 => "00110100",10117 => "00100111",10118 => "10000001",10119 => "10011011",10120 => "11011000",10121 => "00000111",10122 => "00101111",10123 => "01110100",10124 => "10001100",10125 => "00101010",10126 => "01001000",10127 => "11101010",10128 => "11101001",10129 => "11001101",10130 => "11101001",10131 => "10101000",10132 => "01100010",10133 => "10101010",10134 => "11100011",10135 => "10111001",10136 => "10001111",10137 => "00010110",10138 => "11101111",10139 => "01110111",10140 => "01001101",10141 => "11001000",10142 => "01100100",10143 => "00001000",10144 => "01100010",10145 => "11110010",10146 => "10011011",10147 => "10100010",10148 => "10011001",10149 => "00000011",10150 => "10110010",10151 => "11011010",10152 => "11011001",10153 => "01111100",10154 => "11110110",10155 => "11001100",10156 => "00111010",10157 => "01010010",10158 => "00011110",10159 => "01000101",10160 => "10011110",10161 => "11000010",10162 => "11001110",10163 => "11000111",10164 => "00110111",10165 => "00011100",10166 => "10100011",10167 => "10011010",10168 => "01100101",10169 => "00011100",10170 => "00001110",10171 => "01000110",10172 => "01001011",10173 => "11011010",10174 => "10110110",10175 => "11100101",10176 => "00110010",10177 => "01110010",10178 => "10000101",10179 => "00001011",10180 => "01011111",10181 => "01011000",10182 => "01011100",10183 => "00011000",10184 => "11001010",10185 => "00011100",10186 => "10000010",10187 => "00001010",10188 => "01110001",10189 => "01011100",10190 => "01111101",10191 => "00101001",10192 => "10000100",10193 => "00101111",10194 => "01101000",10195 => "10011001",10196 => "11111101",10197 => "11010011",10198 => "01100000",10199 => "01110111",10200 => "00010011",10201 => "10000011",10202 => "11010100",10203 => "00100010",10204 => "01001110",10205 => "10111100",10206 => "11111000",10207 => "01011111",10208 => "01010010",10209 => "10100110",10210 => "10101010",10211 => "00100110",10212 => "11110111",10213 => "00111001",10214 => "01000110",10215 => "01101100",10216 => "10000110",10217 => "10100001",10218 => "01000000",10219 => "00110101",10220 => "00000011",10221 => "00001100",10222 => "10101110",10223 => "00011011",10224 => "10110100",10225 => "10000100",10226 => "10010110",10227 => "01111100",10228 => "10001101",10229 => "00110000",10230 => "00100000",10231 => "11001111",10232 => "01101001",10233 => "00011100",10234 => "10111100",10235 => "01000100",10236 => "10010110",10237 => "00001001",10238 => "10011000",10239 => "00100110",10240 => "00101101",10241 => "01010011",10242 => "00001100",10243 => "01101101",10244 => "00111101",10245 => "10010010",10246 => "01100010",10247 => "11101111",10248 => "01010110",10249 => "01111101",10250 => "11111110",10251 => "00010100",10252 => "00111110",10253 => "01001000",10254 => "10111110",10255 => "00000010",10256 => "01100001",10257 => "00111111",10258 => "10011111",10259 => "10011011",10260 => "01011100",10261 => "00100010",10262 => "10001100",10263 => "10010110",10264 => "11111011",10265 => "11000111",10266 => "11010010",10267 => "10101110",10268 => "11001001",10269 => "01010100",10270 => "10110111",10271 => "00100100",10272 => "00111101",10273 => "01001101",10274 => "10011000",10275 => "10011100",10276 => "00111101",10277 => "11101110",10278 => "11011110",10279 => "01000110",10280 => "11101011",10281 => "01010100",10282 => "00010111",10283 => "11011101",10284 => "10110101",10285 => "10100001",10286 => "01011110",10287 => "01100100",10288 => "01010101",10289 => "00101011",10290 => "10010100",10291 => "10101001",10292 => "01100001",10293 => "10111111",10294 => "11011001",10295 => "10010000",10296 => "10011001",10297 => "00110100",10298 => "11100111",10299 => "10010000",10300 => "01011011",10301 => "01000111",10302 => "10000101",10303 => "00011100",10304 => "11111001",10305 => "11011111",10306 => "11101111",10307 => "00111110",10308 => "01100011",10309 => "10100001",10310 => "11100111",10311 => "01100000",10312 => "10111110",10313 => "11101110",10314 => "10110100",10315 => "10000010",10316 => "01010000",10317 => "10000110",10318 => "11110001",10319 => "01110110",10320 => "11100000",10321 => "10010110",10322 => "11000110",10323 => "00011001",10324 => "11010110",10325 => "00001001",10326 => "01010101",10327 => "10110101",10328 => "10111001",10329 => "11011011",10330 => "01101010",10331 => "01111001",10332 => "00000100",10333 => "00001100",10334 => "01000101",10335 => "10001001",10336 => "11110000",10337 => "00010101",10338 => "01000010",10339 => "10011101",10340 => "10000111",10341 => "01101100",10342 => "10010010",10343 => "10110010",10344 => "11111101",10345 => "10110111",10346 => "11000111",10347 => "01100110",10348 => "10100110",10349 => "11000100",10350 => "01111001",10351 => "10011111",10352 => "00010011",10353 => "00011000",10354 => "00001010",10355 => "00101110",10356 => "01001110",10357 => "10001100",10358 => "00011001",10359 => "00010101",10360 => "01110001",10361 => "01000101",10362 => "10011100",10363 => "10000000",10364 => "00100010",10365 => "11011101",10366 => "00000110",10367 => "01011111",10368 => "11101100",10369 => "10110101",10370 => "10000111",10371 => "00111001",10372 => "01011100",10373 => "11001111",10374 => "01110100",10375 => "00000011",10376 => "11110111",10377 => "11100111",10378 => "10100111",10379 => "11001100",10380 => "01001101",10381 => "10110010",10382 => "01001110",10383 => "11110000",10384 => "11101010",10385 => "11110000",10386 => "10010100",10387 => "10111111",10388 => "11111110",10389 => "10010010",10390 => "01000110",10391 => "10001100",10392 => "10111100",10393 => "10011110",10394 => "10111100",10395 => "01111101",10396 => "10000100",10397 => "10001000",10398 => "11001001",10399 => "01110011",10400 => "01110111",10401 => "10001111",10402 => "00101010",10403 => "00101111",10404 => "01000000",10405 => "10111100",10406 => "10110100",10407 => "10110100",10408 => "00111110",10409 => "11000000",10410 => "11001101",10411 => "01111001",10412 => "10110000",10413 => "01011101",10414 => "11000110",10415 => "10011101",10416 => "10100111",10417 => "00010110",10418 => "11001100",10419 => "11100101",10420 => "10000100",10421 => "10011001",10422 => "00000010",10423 => "01111001",10424 => "11101110",10425 => "01110000",10426 => "10010101",10427 => "11001100",10428 => "01110111",10429 => "10111111",10430 => "00100111",10431 => "10010101",10432 => "00010111",10433 => "10010111",10434 => "00101010",10435 => "11010111",10436 => "11100101",10437 => "10010101",10438 => "11110101",10439 => "01100101",10440 => "01100001",10441 => "00001001",10442 => "01000000",10443 => "01111011",10444 => "00001100",10445 => "00011001",10446 => "00101011",10447 => "01010111",10448 => "11111100",10449 => "11011000",10450 => "11001111",10451 => "01101000",10452 => "00011011",10453 => "01110100",10454 => "10110011",10455 => "10111000",10456 => "01100111",10457 => "01101011",10458 => "11010100",10459 => "10101011",10460 => "11101100",10461 => "01110110",10462 => "11110100",10463 => "10110100",10464 => "10110101",10465 => "10001111",10466 => "00010110",10467 => "00010011",10468 => "11100011",10469 => "01110011",10470 => "10000100",10471 => "11010101",10472 => "01011000",10473 => "10110111",10474 => "10000101",10475 => "10001111",10476 => "00111110",10477 => "00001011",10478 => "01100100",10479 => "11101010",10480 => "11011010",10481 => "11100011",10482 => "00100111",10483 => "01011111",10484 => "00000110",10485 => "10010000",10486 => "10110000",10487 => "10000001",10488 => "11111111",10489 => "01100001",10490 => "01000111",10491 => "01110110",10492 => "11001100",10493 => "00100011",10494 => "11111111",10495 => "11111101",10496 => "10000000",10497 => "00010000",10498 => "11101010",10499 => "10000110",10500 => "00101110",10501 => "11100100",10502 => "00101011",10503 => "00110001",10504 => "00010001",10505 => "10111101",10506 => "00011110",10507 => "01000011",10508 => "10100110",10509 => "11001111",10510 => "10100001",10511 => "01101111",10512 => "10010000",10513 => "01001101",10514 => "01001010",10515 => "11110100",10516 => "00011011",10517 => "01010000",10518 => "10101011",10519 => "11000011",10520 => "10101010",10521 => "10001111",10522 => "10011110",10523 => "10011010",10524 => "00011111",10525 => "01011101",10526 => "10111110",10527 => "10100111",10528 => "10111110",10529 => "10011000",10530 => "00011000",10531 => "00101100",10532 => "01111101",10533 => "01011010",10534 => "01010111",10535 => "10011111",10536 => "01111010",10537 => "01101110",10538 => "00000010",10539 => "00011000",10540 => "00100111",10541 => "10010010",10542 => "11101111",10543 => "10000111",10544 => "00001000",10545 => "00001101",10546 => "10111101",10547 => "01111101",10548 => "00011001",10549 => "00110100",10550 => "10010100",10551 => "00001000",10552 => "11110110",10553 => "10111100",10554 => "11000110",10555 => "10000110",10556 => "11111101",10557 => "01001101",10558 => "00010100",10559 => "00011111",10560 => "00001100",10561 => "01100001",10562 => "01011011",10563 => "01001001",10564 => "10110011",10565 => "00101100",10566 => "01101000",10567 => "01111011",10568 => "00111100",10569 => "01111000",10570 => "10010011",10571 => "11000111",10572 => "00111111",10573 => "01001100",10574 => "01101100",10575 => "10101100",10576 => "11100100",10577 => "10001011",10578 => "01101111",10579 => "10100010",10580 => "11110101",10581 => "11010010",10582 => "10000100",10583 => "10100111",10584 => "11001001",10585 => "10000110",10586 => "00111110",10587 => "11000001",10588 => "01101010",10589 => "01011111",10590 => "00000011",10591 => "10101001",10592 => "10100011",10593 => "01110110",10594 => "01010110",10595 => "10011001",10596 => "10110110",10597 => "01010001",10598 => "00000010",10599 => "00001010",10600 => "11100101",10601 => "11000001",10602 => "11101001",10603 => "00000010",10604 => "01101011",10605 => "01111011",10606 => "01011111",10607 => "11101110",10608 => "01101000",10609 => "10111101",10610 => "01000100",10611 => "10000111",10612 => "00110000",10613 => "01001111",10614 => "00011001",10615 => "10010111",10616 => "10010100",10617 => "01110010",10618 => "11111000",10619 => "01110000",10620 => "10110000",10621 => "00010111",10622 => "10111111",10623 => "10001000",10624 => "11100010",10625 => "00001011",10626 => "01110010",10627 => "11101010",10628 => "10111010",10629 => "01000101",10630 => "11000010",10631 => "11001111",10632 => "11110010",10633 => "00101010",10634 => "01101000",10635 => "00101100",10636 => "10001111",10637 => "00010101",10638 => "01110100",10639 => "01011111",10640 => "00100010",10641 => "10000001",10642 => "10100011",10643 => "11110111",10644 => "00110101",10645 => "10101001",10646 => "01011001",10647 => "01010110",10648 => "01011101",10649 => "00101101",10650 => "00101011",10651 => "00110010",10652 => "00001100",10653 => "00101110",10654 => "01010000",10655 => "11101001",10656 => "10100111",10657 => "00000100",10658 => "11101100",10659 => "11100010",10660 => "11101011",10661 => "10101101",10662 => "10111011",10663 => "11011101",10664 => "01110111",10665 => "10011110",10666 => "00101000",10667 => "10110001",10668 => "00100110",10669 => "00001110",10670 => "00000100",10671 => "00001001",10672 => "01101000",10673 => "00000011",10674 => "10000010",10675 => "10110011",10676 => "01101001",10677 => "10110010",10678 => "11000101",10679 => "00010101",10680 => "01011111",10681 => "00111000",10682 => "00101010",10683 => "00010001",10684 => "01110000",10685 => "10100010",10686 => "10101111",10687 => "00111100",10688 => "10111100",10689 => "10111001",10690 => "11100000",10691 => "01100011",10692 => "11110010",10693 => "01010010",10694 => "01100110",10695 => "01100001",10696 => "00011100",10697 => "00100111",10698 => "10101110",10699 => "11101000",10700 => "10010110",10701 => "11011111",10702 => "00010101",10703 => "11001001",10704 => "01010001",10705 => "11101011",10706 => "00011000",10707 => "10010010",10708 => "11011101",10709 => "00010111",10710 => "10111010",10711 => "11110010",10712 => "01100100",10713 => "00000100",10714 => "01001001",10715 => "10011110",10716 => "10011011",10717 => "00110011",10718 => "11011001",10719 => "10100010",10720 => "00110111",10721 => "11110011",10722 => "01010011",10723 => "01000000",10724 => "00110010",10725 => "01111111",10726 => "10110001",10727 => "00001001",10728 => "11001011",10729 => "00110111",10730 => "01000001",10731 => "00111010",10732 => "00111011",10733 => "00001011",10734 => "00110111",10735 => "10100101",10736 => "11110010",10737 => "11001111",10738 => "00110011",10739 => "00001110",10740 => "11100111",10741 => "10100111",10742 => "10111010",10743 => "00110011",10744 => "00110110",10745 => "10101101",10746 => "11111111",10747 => "10010100",10748 => "00111011",10749 => "00010000",10750 => "10000000",10751 => "00011000",10752 => "01010001",10753 => "00100010",10754 => "10011011",10755 => "00100110",10756 => "01101111",10757 => "01000100",10758 => "01101100",10759 => "00101101",10760 => "00101100",10761 => "10111001",10762 => "01001111",10763 => "11111010",10764 => "00110010",10765 => "11110000",10766 => "11111110",10767 => "00001101",10768 => "00001100",10769 => "01000001",10770 => "01000101",10771 => "00000110",10772 => "00100111",10773 => "00010110",10774 => "10000101",10775 => "00111101",10776 => "01101011",10777 => "01101001",10778 => "00110110",10779 => "00001110",10780 => "10110111",10781 => "00101101",10782 => "01010000",10783 => "10011111",10784 => "01101011",10785 => "11011011",10786 => "11010110",10787 => "10000101",10788 => "11010001",10789 => "00001010",10790 => "11100111",10791 => "11011100",10792 => "11001001",10793 => "00110110",10794 => "00011001",10795 => "10011011",10796 => "10100111",10797 => "11100011",10798 => "10011010",10799 => "01101111",10800 => "00110010",10801 => "00101111",10802 => "01000011",10803 => "11101001",10804 => "11110110",10805 => "11101000",10806 => "11101010",10807 => "10001110",10808 => "01000010",10809 => "00000110",10810 => "11110001",10811 => "10100000",10812 => "10000101",10813 => "11100001",10814 => "01001111",10815 => "00001111",10816 => "10001110",10817 => "01010000",10818 => "10110010",10819 => "00010110",10820 => "01010010",10821 => "00101010",10822 => "11000001",10823 => "10101111",10824 => "10011101",10825 => "00100011",10826 => "10110011",10827 => "01000001",10828 => "11010111",10829 => "01111000",10830 => "00100110",10831 => "10110010",10832 => "10111001",10833 => "10110100",10834 => "01101111",10835 => "01011111",10836 => "10111010",10837 => "01000100",10838 => "11001110",10839 => "10111111",10840 => "00011101",10841 => "11010011",10842 => "10100011",10843 => "10111011",10844 => "11010111",10845 => "11010011",10846 => "01111111",10847 => "00010101",10848 => "00110000",10849 => "01100010",10850 => "11100010",10851 => "01101101",10852 => "01001100",10853 => "10001000",10854 => "01101101",10855 => "11111101",10856 => "01110111",10857 => "10000011",10858 => "00011111",10859 => "01000011",10860 => "10111010",10861 => "00010010",10862 => "01011000",10863 => "11010011",10864 => "00001100",10865 => "00110101",10866 => "01100000",10867 => "00111001",10868 => "00000001",10869 => "00111111",10870 => "11001111",10871 => "00101000",10872 => "10010101",10873 => "01000100",10874 => "11000111",10875 => "10010001",10876 => "01111001",10877 => "10000010",10878 => "01100111",10879 => "00010111",10880 => "01111111",10881 => "11101001",10882 => "10001001",10883 => "11000110",10884 => "01000010",10885 => "00111000",10886 => "00110101",10887 => "10000000",10888 => "11011010",10889 => "11001011",10890 => "11111110",10891 => "00010000",10892 => "00000100",10893 => "01011001",10894 => "01100101",10895 => "10000001",10896 => "10001001",10897 => "10110100",10898 => "01000001",10899 => "10101110",10900 => "00111101",10901 => "11110010",10902 => "11111000",10903 => "00111101",10904 => "11010101",10905 => "00111101",10906 => "10101110",10907 => "11100011",10908 => "00000011",10909 => "11101111",10910 => "00011001",10911 => "10001110",10912 => "00101101",10913 => "00111011",10914 => "00100100",10915 => "10011100",10916 => "01001110",10917 => "11000101",10918 => "10101100",10919 => "10001011",10920 => "00111001",10921 => "01011101",10922 => "11111000",10923 => "11010000",10924 => "01000001",10925 => "01111001",10926 => "00101111",10927 => "00111111",10928 => "10011011",10929 => "10001011",10930 => "00110100",10931 => "00100001",10932 => "10100001",10933 => "11001110",10934 => "10101010",10935 => "01010011",10936 => "10010101",10937 => "10110111",10938 => "00001011",10939 => "11011001",10940 => "01001101",10941 => "11011100",10942 => "00101100",10943 => "00111101",10944 => "00011010",10945 => "00001110",10946 => "11001101",10947 => "10001001",10948 => "00110010",10949 => "00000101",10950 => "10010101",10951 => "00011010",10952 => "00011111",10953 => "11111111",10954 => "01000010",10955 => "10000110",10956 => "11100101",10957 => "01000110",10958 => "10011000",10959 => "01011101",10960 => "00111100",10961 => "10010100",10962 => "10011100",10963 => "00101101",10964 => "00010000",10965 => "01100111",10966 => "01101111",10967 => "01111110",10968 => "11000010",10969 => "00000111",10970 => "01111000",10971 => "10000010",10972 => "00100101",10973 => "11001011",10974 => "01101011",10975 => "01110110",10976 => "01001000",10977 => "10011111",10978 => "01011100",10979 => "01110101",10980 => "10110000",10981 => "00100100",10982 => "00100001",10983 => "00101110",10984 => "01001111",10985 => "01011100",10986 => "00111111",10987 => "01010101",10988 => "10100010",10989 => "01010010",10990 => "11111110",10991 => "11101010",10992 => "10100110",10993 => "00011010",10994 => "10011001",10995 => "01101001",10996 => "01110101",10997 => "00010101",10998 => "01100110",10999 => "00001010",11000 => "00101111",11001 => "10011110",11002 => "01110000",11003 => "00111111",11004 => "11000110",11005 => "10100000",11006 => "00111000",11007 => "00001111",11008 => "00010011",11009 => "11101000",11010 => "00100111",11011 => "11111001",11012 => "11111101",11013 => "00000110",11014 => "10110110",11015 => "00100011",11016 => "00111001",11017 => "01010101",11018 => "10111001",11019 => "00000111",11020 => "00111010",11021 => "01011000",11022 => "11010110",11023 => "01000010",11024 => "10010010",11025 => "01110010",11026 => "11101011",11027 => "01001101",11028 => "10011111",11029 => "01001000",11030 => "00000000",11031 => "10010110",11032 => "11100101",11033 => "00001010",11034 => "00010101",11035 => "10101111",11036 => "10001000",11037 => "00110111",11038 => "10000010",11039 => "10111010",11040 => "11101010",11041 => "11101101",11042 => "11000000",11043 => "01111101",11044 => "01101100",11045 => "00000110",11046 => "01000000",11047 => "10010101",11048 => "00001001",11049 => "10100101",11050 => "10011101",11051 => "10101101",11052 => "00000010",11053 => "11101111",11054 => "10011111",11055 => "00111000",11056 => "01100100",11057 => "00011110",11058 => "00001010",11059 => "10110110",11060 => "11100011",11061 => "10101101",11062 => "11010010",11063 => "10011100",11064 => "00001111",11065 => "00000011",11066 => "10011111",11067 => "01111100",11068 => "01100111",11069 => "10010101",11070 => "00110011",11071 => "00010011",11072 => "10101100",11073 => "00000001",11074 => "10011101",11075 => "01011001",11076 => "01101100",11077 => "11110010",11078 => "01110101",11079 => "10011100",11080 => "11000100",11081 => "11011010",11082 => "10101111",11083 => "01100011",11084 => "01111000",11085 => "00111011",11086 => "10111010",11087 => "11001001",11088 => "00111100",11089 => "10101101",11090 => "10100100",11091 => "00010011",11092 => "11110110",11093 => "11111101",11094 => "01001011",11095 => "10111101",11096 => "10101101",11097 => "00110001",11098 => "11011101",11099 => "10111110",11100 => "00001110",11101 => "01110001",11102 => "10111100",11103 => "11111010",11104 => "01110010",11105 => "00101110",11106 => "10100000",11107 => "01110101",11108 => "10111010",11109 => "11110001",11110 => "10110010",11111 => "10110110",11112 => "00010100",11113 => "01011000",11114 => "01001101",11115 => "11000011",11116 => "11010110",11117 => "00111011",11118 => "11110100",11119 => "10101000",11120 => "01010010",11121 => "10111010",11122 => "10100001",11123 => "01001101",11124 => "10010011",11125 => "01011101",11126 => "01110111",11127 => "10010010",11128 => "11001010",11129 => "00010111",11130 => "11111101",11131 => "11010110",11132 => "00110010",11133 => "11110101",11134 => "11001011",11135 => "00011100",11136 => "00000001",11137 => "11001001",11138 => "00110011",11139 => "01101001",11140 => "01101111",11141 => "01100111",11142 => "01110110",11143 => "01101000",11144 => "10111011",11145 => "11010010",11146 => "01000001",11147 => "10111101",11148 => "00111110",11149 => "01100010",11150 => "10101011",11151 => "11101100",11152 => "00000001",11153 => "10010101",11154 => "10101010",11155 => "00101000",11156 => "01111001",11157 => "01001000",11158 => "11011001",11159 => "11010010",11160 => "10010000",11161 => "10000000",11162 => "01001010",11163 => "00111001",11164 => "00110001",11165 => "01010110",11166 => "00101011",11167 => "11101000",11168 => "01101110",11169 => "11100101",11170 => "00000110",11171 => "11000101",11172 => "01111110",11173 => "11101101",11174 => "11100011",11175 => "10001010",11176 => "01111000",11177 => "10010010",11178 => "01000000",11179 => "10111001",11180 => "01101011",11181 => "00101110",11182 => "11111000",11183 => "10010111",11184 => "10110001",11185 => "10010111",11186 => "11000001",11187 => "00011010",11188 => "11110000",11189 => "01011111",11190 => "11111110",11191 => "10100110",11192 => "01111101",11193 => "11100111",11194 => "01001011",11195 => "11110111",11196 => "01111110",11197 => "01000100",11198 => "01011011",11199 => "10011010",11200 => "10110000",11201 => "10000011",11202 => "01111001",11203 => "11010100",11204 => "00000001",11205 => "01011011",11206 => "10001111",11207 => "00000001",11208 => "10111101",11209 => "00110100",11210 => "01000110",11211 => "10101010",11212 => "10111110",11213 => "00101010",11214 => "01010000",11215 => "00100101",11216 => "10101001",11217 => "00110110",11218 => "10011111",11219 => "10011001",11220 => "01010000",11221 => "01000111",11222 => "00111000",11223 => "10110010",11224 => "11110000",11225 => "11100101",11226 => "00111101",11227 => "11111111",11228 => "01011010",11229 => "11110111",11230 => "10101101",11231 => "11000010",11232 => "10010001",11233 => "01100000",11234 => "11011010",11235 => "11110101",11236 => "01000000",11237 => "00000110",11238 => "10111011",11239 => "10111001",11240 => "10010100",11241 => "01111010",11242 => "00011000",11243 => "01000000",11244 => "11010001",11245 => "01011010",11246 => "01111101",11247 => "11001000",11248 => "10100101",11249 => "01111101",11250 => "01011110",11251 => "01010111",11252 => "10000000",11253 => "11011101",11254 => "01010100",11255 => "10101111",11256 => "00101100",11257 => "11110000",11258 => "00001100",11259 => "11000110",11260 => "10010100",11261 => "10011010",11262 => "11100101",11263 => "01011100",11264 => "01011101",11265 => "00001100",11266 => "11110010",11267 => "01001010",11268 => "00101111",11269 => "01100000",11270 => "00000111",11271 => "11101010",11272 => "00100010",11273 => "11110111",11274 => "01000111",11275 => "10000111",11276 => "11001001",11277 => "10001011",11278 => "00001001",11279 => "00011110",11280 => "01001010",11281 => "00000001",11282 => "01001000",11283 => "00001101",11284 => "11010111",11285 => "10000001",11286 => "10000111",11287 => "01011000",11288 => "10010111",11289 => "00010100",11290 => "10011101",11291 => "11100100",11292 => "11001111",11293 => "01110100",11294 => "00110100",11295 => "00000110",11296 => "11110001",11297 => "11100010",11298 => "10111110",11299 => "01100011",11300 => "01000110",11301 => "11110110",11302 => "11101100",11303 => "10010011",11304 => "00100101",11305 => "11000000",11306 => "11100010",11307 => "01111111",11308 => "00100110",11309 => "01101111",11310 => "10100110",11311 => "11011110",11312 => "11100100",11313 => "10110111",11314 => "11011001",11315 => "10101001",11316 => "01110010",11317 => "11001011",11318 => "00101000",11319 => "11100011",11320 => "00011001",11321 => "00011001",11322 => "10010111",11323 => "11100000",11324 => "01111010",11325 => "10100011",11326 => "10110100",11327 => "00011100",11328 => "11110011",11329 => "10110100",11330 => "00000001",11331 => "11110010",11332 => "01010010",11333 => "01001101",11334 => "01101110",11335 => "10111100",11336 => "01101110",11337 => "01010110",11338 => "11110010",11339 => "01101111",11340 => "00000011",11341 => "00101011",11342 => "00010000",11343 => "01101111",11344 => "00010110",11345 => "11101100",11346 => "11111100",11347 => "11101110",11348 => "11001001",11349 => "00111111",11350 => "00111011",11351 => "00101001",11352 => "00100110",11353 => "11010100",11354 => "11110110",11355 => "10011010",11356 => "10110011",11357 => "11000010",11358 => "11110000",11359 => "00000111",11360 => "11111010",11361 => "00100000",11362 => "11011011",11363 => "01110100",11364 => "01101010",11365 => "10101110",11366 => "00000111",11367 => "11000001",11368 => "00110001",11369 => "10101001",11370 => "11010000",11371 => "01011111",11372 => "10010000",11373 => "10000101",11374 => "01011101",11375 => "11111101",11376 => "11111001",11377 => "11000000",11378 => "01100100",11379 => "01000010",11380 => "11111110",11381 => "01100001",11382 => "01100111",11383 => "10111011",11384 => "11111100",11385 => "01111100",11386 => "00001101",11387 => "00100100",11388 => "11001100",11389 => "00110011",11390 => "00001110",11391 => "10100110",11392 => "11011111",11393 => "01111101",11394 => "00111111",11395 => "00101011",11396 => "10000111",11397 => "11011111",11398 => "10111101",11399 => "10100100",11400 => "10101001",11401 => "11111001",11402 => "01011010",11403 => "11000110",11404 => "00111110",11405 => "00111100",11406 => "11011010",11407 => "01000111",11408 => "10100001",11409 => "00110001",11410 => "11011111",11411 => "10101001",11412 => "10000011",11413 => "00001000",11414 => "10111111",11415 => "10010001",11416 => "11011001",11417 => "01000001",11418 => "11101111",11419 => "11100111",11420 => "11000011",11421 => "11011010",11422 => "10100010",11423 => "11001001",11424 => "01100000",11425 => "01100011",11426 => "01001100",11427 => "11011100",11428 => "00011111",11429 => "10100101",11430 => "11000000",11431 => "01111000",11432 => "10110110",11433 => "01101001",11434 => "00111000",11435 => "01000011",11436 => "00101100",11437 => "11010111",11438 => "00100001",11439 => "11001001",11440 => "10001001",11441 => "11110101",11442 => "11100100",11443 => "11110001",11444 => "11111011",11445 => "01100110",11446 => "01011111",11447 => "01011000",11448 => "00001101",11449 => "11010000",11450 => "00010001",11451 => "10101000",11452 => "01100000",11453 => "01000110",11454 => "11011111",11455 => "00011110",11456 => "01010111",11457 => "11001001",11458 => "11001010",11459 => "11010111",11460 => "11011011",11461 => "11110010",11462 => "11101011",11463 => "10001001",11464 => "11100001",11465 => "01110000",11466 => "10100100",11467 => "01110111",11468 => "11111111",11469 => "11101011",11470 => "01110001",11471 => "01011010",11472 => "10111010",11473 => "11000010",11474 => "11010001",11475 => "00100110",11476 => "11111111",11477 => "01000000",11478 => "00000100",11479 => "10101011",11480 => "10001000",11481 => "00010011",11482 => "11111100",11483 => "00001110",11484 => "10101010",11485 => "01111001",11486 => "11100011",11487 => "11100010",11488 => "01000011",11489 => "10011101",11490 => "11101100",11491 => "01001000",11492 => "10101111",11493 => "11100101",11494 => "01111011",11495 => "01100000",11496 => "00000111",11497 => "11011010",11498 => "10010010",11499 => "11010110",11500 => "01010000",11501 => "00100001",11502 => "00111011",11503 => "10111111",11504 => "00101111",11505 => "00111100",11506 => "01110110",11507 => "00011011",11508 => "01100100",11509 => "00101001",11510 => "01111111",11511 => "01100111",11512 => "01101011",11513 => "11000001",11514 => "01110011",11515 => "01010010",11516 => "00111000",11517 => "00011001",11518 => "10011011",11519 => "01001100",11520 => "10100011",11521 => "01010100",11522 => "00101101",11523 => "10011000",11524 => "10101010",11525 => "01101000",11526 => "11111111",11527 => "01000101",11528 => "11011100",11529 => "01010101",11530 => "11000000",11531 => "10101011",11532 => "11111110",11533 => "10011111",11534 => "11010010",11535 => "10011100",11536 => "01101010",11537 => "01111110",11538 => "00110111",11539 => "01101110",11540 => "01000010",11541 => "00001010",11542 => "01010001",11543 => "00010101",11544 => "11000010",11545 => "01111110",11546 => "01111001",11547 => "10100000",11548 => "10111101",11549 => "11100011",11550 => "01011101",11551 => "10101000",11552 => "00100000",11553 => "01111101",11554 => "11000011",11555 => "01010011",11556 => "11110001",11557 => "11001101",11558 => "00110110",11559 => "11111001",11560 => "01010010",11561 => "10011110",11562 => "10110011",11563 => "00001010",11564 => "11101010",11565 => "11101101",11566 => "10111000",11567 => "10001000",11568 => "11101111",11569 => "11010010",11570 => "10100010",11571 => "01010111",11572 => "00010111",11573 => "00001100",11574 => "10010111",11575 => "01001101",11576 => "10001011",11577 => "01101011",11578 => "00001001",11579 => "00110010",11580 => "10101111",11581 => "10010010",11582 => "01111110",11583 => "01100110",11584 => "01110111",11585 => "00111000",11586 => "00011101",11587 => "01000001",11588 => "01111111",11589 => "10011010",11590 => "00111110",11591 => "11101011",11592 => "10010000",11593 => "10101010",11594 => "01100110",11595 => "01101111",11596 => "01010011",11597 => "01000010",11598 => "10111101",11599 => "01110001",11600 => "11100010",11601 => "10101111",11602 => "10010111",11603 => "00110000",11604 => "11000110",11605 => "01101111",11606 => "11000011",11607 => "11111110",11608 => "00011010",11609 => "00001100",11610 => "00001010",11611 => "01001000",11612 => "11111010",11613 => "10111011",11614 => "01000111",11615 => "10001111",11616 => "00011010",11617 => "11110011",11618 => "00010000",11619 => "00101101",11620 => "11110100",11621 => "11101001",11622 => "00110010",11623 => "01101111",11624 => "01010110",11625 => "11001101",11626 => "01011100",11627 => "00001111",11628 => "01110110",11629 => "11110010",11630 => "11001000",11631 => "11010100",11632 => "10001111",11633 => "11011100",11634 => "11100010",11635 => "01011110",11636 => "11000111",11637 => "01101010",11638 => "00111011",11639 => "10111110",11640 => "00110101",11641 => "10111001",11642 => "11011101",11643 => "11000101",11644 => "00110110",11645 => "11101010",11646 => "10000000",11647 => "11100111",11648 => "10011100",11649 => "10011101",11650 => "11101100",11651 => "11101111",11652 => "01111010",11653 => "11000000",11654 => "10111010",11655 => "10010110",11656 => "11101010",11657 => "10100010",11658 => "01101011",11659 => "10000101",11660 => "11001011",11661 => "01101111",11662 => "10000110",11663 => "10111100",11664 => "01011111",11665 => "10010111",11666 => "01100010",11667 => "00000110",11668 => "01110101",11669 => "11010010",11670 => "01000010",11671 => "11000001",11672 => "10100011",11673 => "10011111",11674 => "00111010",11675 => "10111101",11676 => "01001011",11677 => "11110000",11678 => "01110110",11679 => "01111001",11680 => "10101110",11681 => "00110110",11682 => "11000011",11683 => "01011100",11684 => "11111111",11685 => "00110100",11686 => "00010100",11687 => "01011110",11688 => "11000011",11689 => "00100110",11690 => "10110011",11691 => "00000111",11692 => "00011101",11693 => "11010011",11694 => "10010001",11695 => "10100001",11696 => "00100101",11697 => "11110111",11698 => "10111000",11699 => "00100010",11700 => "10011001",11701 => "11100100",11702 => "10110010",11703 => "10101100",11704 => "01000101",11705 => "11010011",11706 => "10100001",11707 => "01010111",11708 => "10101111",11709 => "00000101",11710 => "10100110",11711 => "10010011",11712 => "11100100",11713 => "11001011",11714 => "01011010",11715 => "10010100",11716 => "10101011",11717 => "11111010",11718 => "10001111",11719 => "00100010",11720 => "10110100",11721 => "01011111",11722 => "01100010",11723 => "00000010",11724 => "01001010",11725 => "11101011",11726 => "01111010",11727 => "01111110",11728 => "00011100",11729 => "01010111",11730 => "01110110",11731 => "11011101",11732 => "01100101",11733 => "10111110",11734 => "11100001",11735 => "00110101",11736 => "11110001",11737 => "00100000",11738 => "01111101",11739 => "00010111",11740 => "10101101",11741 => "11000011",11742 => "01101000",11743 => "01010001",11744 => "00100001",11745 => "10100011",11746 => "10110011",11747 => "01110110",11748 => "11000011",11749 => "11110001",11750 => "10111010",11751 => "00010010",11752 => "11100101",11753 => "11100011",11754 => "01101110",11755 => "01100011",11756 => "01110110",11757 => "11100000",11758 => "00001100",11759 => "00110010",11760 => "10011001",11761 => "01111100",11762 => "11111101",11763 => "11110111",11764 => "10000011",11765 => "11001110",11766 => "01100110",11767 => "01000110",11768 => "10011110",11769 => "01101101",11770 => "11011000",11771 => "00011011",11772 => "01000110",11773 => "00100110",11774 => "11000001",11775 => "10001100",11776 => "10000111",11777 => "10110101",11778 => "00000100",11779 => "01110100",11780 => "00000001",11781 => "11011100",11782 => "01000110",11783 => "10000100",11784 => "00110111",11785 => "00000011",11786 => "10001101",11787 => "10111110",11788 => "11100101",11789 => "01100101",11790 => "10010010",11791 => "00001100",11792 => "01010011",11793 => "00000111",11794 => "11100100",11795 => "10101111",11796 => "10100111",11797 => "10101000",11798 => "00000001",11799 => "11111011",11800 => "01000010",11801 => "01011110",11802 => "11100010",11803 => "01111000",11804 => "11110111",11805 => "01111011",11806 => "10001110",11807 => "00010111",11808 => "01011100",11809 => "01100011",11810 => "01110011",11811 => "11100101",11812 => "10110101",11813 => "00110111",11814 => "01011101",11815 => "11100111",11816 => "10111100",11817 => "00100101",11818 => "00001101",11819 => "00101110",11820 => "01111000",11821 => "11101000",11822 => "11001110",11823 => "00100010",11824 => "10100111",11825 => "00101111",11826 => "11010001",11827 => "01001100",11828 => "00010111",11829 => "01101110",11830 => "01001000",11831 => "10100101",11832 => "10100111",11833 => "01100111",11834 => "00010000",11835 => "01111001",11836 => "11110110",11837 => "00011111",11838 => "11000010",11839 => "00111001",11840 => "00111110",11841 => "10100010",11842 => "10101010",11843 => "01110100",11844 => "00011101",11845 => "01111011",11846 => "11001001",11847 => "00110101",11848 => "11110011",11849 => "00101010",11850 => "01110100",11851 => "00101110",11852 => "10011100",11853 => "01101110",11854 => "11011100",11855 => "10110101",11856 => "00111110",11857 => "10010010",11858 => "10110011",11859 => "11111000",11860 => "11011011",11861 => "11011010",11862 => "01111100",11863 => "01001101",11864 => "11111011",11865 => "00110011",11866 => "11111000",11867 => "01001110",11868 => "11110101",11869 => "11101101",11870 => "01010011",11871 => "01011101",11872 => "00000000",11873 => "00110001",11874 => "11010001",11875 => "10100100",11876 => "11010111",11877 => "10101000",11878 => "01000001",11879 => "11001000",11880 => "01100010",11881 => "01011100",11882 => "01111010",11883 => "01000101",11884 => "00000001",11885 => "01110101",11886 => "10110001",11887 => "00011011",11888 => "10111001",11889 => "10111100",11890 => "10101010",11891 => "10101010",11892 => "00110010",11893 => "01110010",11894 => "00100110",11895 => "00110000",11896 => "11111110",11897 => "01010111",11898 => "11010110",11899 => "10000000",11900 => "00010111",11901 => "11010000",11902 => "01110110",11903 => "01011000",11904 => "11100100",11905 => "11000011",11906 => "11111000",11907 => "10011101",11908 => "10000010",11909 => "11110001",11910 => "11101000",11911 => "11101010",11912 => "00010011",11913 => "10101010",11914 => "01110001",11915 => "10111001",11916 => "00101010",11917 => "00111011",11918 => "10100100",11919 => "10110101",11920 => "00100001",11921 => "00011111",11922 => "10101001",11923 => "11000100",11924 => "00111111",11925 => "10100001",11926 => "11100110",11927 => "10111010",11928 => "00011010",11929 => "11110110",11930 => "01001001",11931 => "01100010",11932 => "10001010",11933 => "01100011",11934 => "01001110",11935 => "00111001",11936 => "01110111",11937 => "11111100",11938 => "01011100",11939 => "11100101",11940 => "01111000",11941 => "11001111",11942 => "01110110",11943 => "01100011",11944 => "11110010",11945 => "01010010",11946 => "10101011",11947 => "00011010",11948 => "00111111",11949 => "11110010",11950 => "00011111",11951 => "00000110",11952 => "10001110",11953 => "10110100",11954 => "01010011",11955 => "11000111",11956 => "10010111",11957 => "01110010",11958 => "01011101",11959 => "10101001",11960 => "00011001",11961 => "00111100",11962 => "01011001",11963 => "00001100",11964 => "01100110",11965 => "11000001",11966 => "10000100",11967 => "00010000",11968 => "11011111",11969 => "10100001",11970 => "10110010",11971 => "00111001",11972 => "10111100",11973 => "10101000",11974 => "10010101",11975 => "00010000",11976 => "01110111",11977 => "00011011",11978 => "00101001",11979 => "01000011",11980 => "01101001",11981 => "11000101",11982 => "01010010",11983 => "11011100",11984 => "10110100",11985 => "00010001",11986 => "01110101",11987 => "10101101",11988 => "11100110",11989 => "10010001",11990 => "01011110",11991 => "01000111",11992 => "00100010",11993 => "11110101",11994 => "00010110",11995 => "10100101",11996 => "00101110",11997 => "11110011",11998 => "00111101",11999 => "11000111",12000 => "00100111",12001 => "00001010",12002 => "11010001",12003 => "00111100",12004 => "01010011",12005 => "11010111",12006 => "00001010",12007 => "01111110",12008 => "10000101",12009 => "01011100",12010 => "00011111",12011 => "00110010",12012 => "01001100",12013 => "00111110",12014 => "01001101",12015 => "11011100",12016 => "10110101",12017 => "01011001",12018 => "00010010",12019 => "10100111",12020 => "11100100",12021 => "10011110",12022 => "11100111",12023 => "00110101",12024 => "11100111",12025 => "10110110",12026 => "11101110",12027 => "00101010",12028 => "00011101",12029 => "11111100",12030 => "11010110",12031 => "01100011",12032 => "00011000",12033 => "01001101",12034 => "00011101",12035 => "10010011",12036 => "01010001",12037 => "00111111",12038 => "00011010",12039 => "10011000",12040 => "00000101",12041 => "11100000",12042 => "00111100",12043 => "01111100",12044 => "10011001",12045 => "11101110",12046 => "00101010",12047 => "11111001",12048 => "00011101",12049 => "11101000",12050 => "01011011",12051 => "01101000",12052 => "11000010",12053 => "00110010",12054 => "11110001",12055 => "10000100",12056 => "00111100",12057 => "01101011",12058 => "11110011",12059 => "00100110",12060 => "01111010",12061 => "11100011",12062 => "00110101",12063 => "10011001",12064 => "00100000",12065 => "01100111",12066 => "11111001",12067 => "01000010",12068 => "10000101",12069 => "00101001",12070 => "10011100",12071 => "11010011",12072 => "11000101",12073 => "01000111",12074 => "11001000",12075 => "11101000",12076 => "10010010",12077 => "11110000",12078 => "11011011",12079 => "01111011",12080 => "00001111",12081 => "11001100",12082 => "10110001",12083 => "01001011",12084 => "00000110",12085 => "00110101",12086 => "01011101",12087 => "10011001",12088 => "11101111",12089 => "11101011",12090 => "10011100",12091 => "01111100",12092 => "11010110",12093 => "00010111",12094 => "00011110",12095 => "00110001",12096 => "11011111",12097 => "01101000",12098 => "10110011",12099 => "11100010",12100 => "10010010",12101 => "10010001",12102 => "11001000",12103 => "01110101",12104 => "00111100",12105 => "10111101",12106 => "01100010",12107 => "00001111",12108 => "10101111",12109 => "01000110",12110 => "11001111",12111 => "10011111",12112 => "00010011",12113 => "00111100",12114 => "11101110",12115 => "01001111",12116 => "01101111",12117 => "10100001",12118 => "11010001",12119 => "10101101",12120 => "10011011",12121 => "00001100",12122 => "11000010",12123 => "11010100",12124 => "11111100",12125 => "11001001",12126 => "10100010",12127 => "11110101",12128 => "11110101",12129 => "11110101",12130 => "00010101",12131 => "10001101",12132 => "10111100",12133 => "01011101",12134 => "00101101",12135 => "00001011",12136 => "00010000",12137 => "01001110",12138 => "10100011",12139 => "01011111",12140 => "11010011",12141 => "10111010",12142 => "01000101",12143 => "01000000",12144 => "11000110",12145 => "10010001",12146 => "01110001",12147 => "00101101",12148 => "00000100",12149 => "10011010",12150 => "11110110",12151 => "01010100",12152 => "10111011",12153 => "00100010",12154 => "00101111",12155 => "01101100",12156 => "01010011",12157 => "00111010",12158 => "01001111",12159 => "01001010",12160 => "11000111",12161 => "00101110",12162 => "00100010",12163 => "01111001",12164 => "10100110",12165 => "00101101",12166 => "00011011",12167 => "10011101",12168 => "00010011",12169 => "00100111",12170 => "00111010",12171 => "01100000",12172 => "10101100",12173 => "00010011",12174 => "11010001",12175 => "00110101",12176 => "01010000",12177 => "00011001",12178 => "11101100",12179 => "00011001",12180 => "01100110",12181 => "11010110",12182 => "00100110",12183 => "11111010",12184 => "11010000",12185 => "01101010",12186 => "01111010",12187 => "01111110",12188 => "11011010",12189 => "11110101",12190 => "00111010",12191 => "00010110",12192 => "10011110",12193 => "00110011",12194 => "11111111",12195 => "10111011",12196 => "00100111",12197 => "11011111",12198 => "11011100",12199 => "00110011",12200 => "00000011",12201 => "10011111",12202 => "01110110",12203 => "01000110",12204 => "11001100",12205 => "00010011",12206 => "00100100",12207 => "10011111",12208 => "11111001",12209 => "01100000",12210 => "10000111",12211 => "11111001",12212 => "10001010",12213 => "01110001",12214 => "00100100",12215 => "00110000",12216 => "11001110",12217 => "10111001",12218 => "11000000",12219 => "10011010",12220 => "11110000",12221 => "01111010",12222 => "11010110",12223 => "00001100",12224 => "01000010",12225 => "00110001",12226 => "11010010",12227 => "00000100",12228 => "11010100",12229 => "00100110",12230 => "01001111",12231 => "10100001",12232 => "01011001",12233 => "00101001",12234 => "01011100",12235 => "00010111",12236 => "10010101",12237 => "00111100",12238 => "10101100",12239 => "11010011",12240 => "10010011",12241 => "10010010",12242 => "01010011",12243 => "10110010",12244 => "11011010",12245 => "01011111",12246 => "01010010",12247 => "01010000",12248 => "00010100",12249 => "10110000",12250 => "01010010",12251 => "00111111",12252 => "01010001",12253 => "10011010",12254 => "00011011",12255 => "11110010",12256 => "10101100",12257 => "01001111",12258 => "10111011",12259 => "01010101",12260 => "00101000",12261 => "11110001",12262 => "10111101",12263 => "11011101",12264 => "11100101",12265 => "00100111",12266 => "10011111",12267 => "10111010",12268 => "11101011",12269 => "11010101",12270 => "11101000",12271 => "01100110",12272 => "11011000",12273 => "11111111",12274 => "10001000",12275 => "01011011",12276 => "10011101",12277 => "11100110",12278 => "00001001",12279 => "11000101",12280 => "01011101",12281 => "10001110",12282 => "11101110",12283 => "00111011",12284 => "01000001",12285 => "11001000",12286 => "11111001",12287 => "01010010",12288 => "01101110",12289 => "01111110",12290 => "01011110",12291 => "11110000",12292 => "01000011",12293 => "01100011",12294 => "11000000",12295 => "10011000",12296 => "10111010",12297 => "11011000",12298 => "00011111",12299 => "00011011",12300 => "00100011",12301 => "01100000",12302 => "10100001",12303 => "00011000",12304 => "01100011",12305 => "01010001",12306 => "01011110",12307 => "00011110",12308 => "10100100",12309 => "11001100",12310 => "01101100",12311 => "00001100",12312 => "00011011",12313 => "10101000",12314 => "01010111",12315 => "10000000",12316 => "01110110",12317 => "11000000",12318 => "01111110",12319 => "01001011",12320 => "01001001",12321 => "11101110",12322 => "10011110",12323 => "10110001",12324 => "00110011",12325 => "00101010",12326 => "10110101",12327 => "01110011",12328 => "01000101",12329 => "10110001",12330 => "01101000",12331 => "10000001",12332 => "00011110",12333 => "01110010",12334 => "10101101",12335 => "01001100",12336 => "10100101",12337 => "01111001",12338 => "11000111",12339 => "10011110",12340 => "11101001",12341 => "01001001",12342 => "10001110",12343 => "11011100",12344 => "01110001",12345 => "00111011",12346 => "01001010",12347 => "10111000",12348 => "10001111",12349 => "00000000",12350 => "00111011",12351 => "10010000",12352 => "01100100",12353 => "01110110",12354 => "01110010",12355 => "00110110",12356 => "11011101",12357 => "01101111",12358 => "01010011",12359 => "00110010",12360 => "00001101",12361 => "11111000",12362 => "10101001",12363 => "11110011",12364 => "01101100",12365 => "10010001",12366 => "11010110",12367 => "00000100",12368 => "11101100",12369 => "00000001",12370 => "00011101",12371 => "00110101",12372 => "10011100",12373 => "10100001",12374 => "10010101",12375 => "10001000",12376 => "10001000",12377 => "00111110",12378 => "11011101",12379 => "10010111",12380 => "11110011",12381 => "11101101",12382 => "11111010",12383 => "10001100",12384 => "00100011",12385 => "11100111",12386 => "11111000",12387 => "11111001",12388 => "01010100",12389 => "11101100",12390 => "11110100",12391 => "01101000",12392 => "11001010",12393 => "10000111",12394 => "10010110",12395 => "10011111",12396 => "00011101",12397 => "10100111",12398 => "01000101",12399 => "01000010",12400 => "11010011",12401 => "00001100",12402 => "01001001",12403 => "01111101",12404 => "11011000",12405 => "01111111",12406 => "11100011",12407 => "10101110",12408 => "01100111",12409 => "10001111",12410 => "11010110",12411 => "10010001",12412 => "11010100",12413 => "01101100",12414 => "10001001",12415 => "01000100",12416 => "11100111",12417 => "01001110",12418 => "00011000",12419 => "00100010",12420 => "00001001",12421 => "00101101",12422 => "00010101",12423 => "10000010",12424 => "10110100",12425 => "00000100",12426 => "10001111",12427 => "00110111",12428 => "01110000",12429 => "11010111",12430 => "11110101",12431 => "01101111",12432 => "10011111",12433 => "11000110",12434 => "00100101",12435 => "00100011",12436 => "10000111",12437 => "01111001",12438 => "11000101",12439 => "11010010",12440 => "01111100",12441 => "10111011",12442 => "11001000",12443 => "00101010",12444 => "10101011",12445 => "01101010",12446 => "10111100",12447 => "11001110",12448 => "10010111",12449 => "11100010",12450 => "11011000",12451 => "10010101",12452 => "11101010",12453 => "10110111",12454 => "11101110",12455 => "00111100",12456 => "10100101",12457 => "01100000",12458 => "00000011",12459 => "10001101",12460 => "11011111",12461 => "10001000",12462 => "01011110",12463 => "00111100",12464 => "10001111",12465 => "00111010",12466 => "10001110",12467 => "10101011",12468 => "01111000",12469 => "01101111",12470 => "01010100",12471 => "01101110",12472 => "01100010",12473 => "00000100",12474 => "11110111",12475 => "11011010",12476 => "10011111",12477 => "01101100",12478 => "11111000",12479 => "00111101",12480 => "00011101",12481 => "11100010",12482 => "10110110",12483 => "11110010",12484 => "11010001",12485 => "10011100",12486 => "00001011",12487 => "01000000",12488 => "01111110",12489 => "10110010",12490 => "00011100",12491 => "11101101",12492 => "01110010",12493 => "01010111",12494 => "00111100",12495 => "11000000",12496 => "10111001",12497 => "00101111",12498 => "00010000",12499 => "11101001",12500 => "10110111",12501 => "11100100",12502 => "01011111",12503 => "10101101",12504 => "01111111",12505 => "01110111",12506 => "10100001",12507 => "11100011",12508 => "11101110",12509 => "01110111",12510 => "00010101",12511 => "01110101",12512 => "00110111",12513 => "10010000",12514 => "11110100",12515 => "01011110",12516 => "00010000",12517 => "01001100",12518 => "10100101",12519 => "00110110",12520 => "01110001",12521 => "10101101",12522 => "00001000",12523 => "10000111",12524 => "10110010",12525 => "10010011",12526 => "11010011",12527 => "11110000",12528 => "01111000",12529 => "01111110",12530 => "00000101",12531 => "01001011",12532 => "10001010",12533 => "00001000",12534 => "10100101",12535 => "10010100",12536 => "11011101",12537 => "11000000",12538 => "10001010",12539 => "11000011",12540 => "11001010",12541 => "10101110",12542 => "10100100",12543 => "10011010",12544 => "10001010",12545 => "11101011",12546 => "10010100",12547 => "00000111",12548 => "11100011",12549 => "10000111",12550 => "10100011",12551 => "00110011",12552 => "01000110",12553 => "01010101",12554 => "11101010",12555 => "10000010",12556 => "10101110",12557 => "10101010",12558 => "10100100",12559 => "10011111",12560 => "10001000",12561 => "00100111",12562 => "11101001",12563 => "11001111",12564 => "11110000",12565 => "00011101",12566 => "00110100",12567 => "11111110",12568 => "01001011",12569 => "00011101",12570 => "11110110",12571 => "10111001",12572 => "11010101",12573 => "01111011",12574 => "10110110",12575 => "11001101",12576 => "00110001",12577 => "11111000",12578 => "11101010",12579 => "10011101",12580 => "00110101",12581 => "01111010",12582 => "10110101",12583 => "10101010",12584 => "11000111",12585 => "11110000",12586 => "00011011",12587 => "01000101",12588 => "10111111",12589 => "10111000",12590 => "01100101",12591 => "00000100",12592 => "11100011",12593 => "11101110",12594 => "10101001",12595 => "01010001",12596 => "00101011",12597 => "10110111",12598 => "10000101",12599 => "10010111",12600 => "00000000",12601 => "11010000",12602 => "00010100",12603 => "01110000",12604 => "11001001",12605 => "00100111",12606 => "11100111",12607 => "10011000",12608 => "10101111",12609 => "00101010",12610 => "10111001",12611 => "11100010",12612 => "11111011",12613 => "00011101",12614 => "11001000",12615 => "00111110",12616 => "10001100",12617 => "10111000",12618 => "11111111",12619 => "11111101",12620 => "01101011",12621 => "11010100",12622 => "11011110",12623 => "00111000",12624 => "10011110",12625 => "00100000",12626 => "01000110",12627 => "10010010",12628 => "01110000",12629 => "01101100",12630 => "01100011",12631 => "11000110",12632 => "01111011",12633 => "00001110",12634 => "11110100",12635 => "00101010",12636 => "10111111",12637 => "10010001",12638 => "01010110",12639 => "11000011",12640 => "01000011",12641 => "11101110",12642 => "01101100",12643 => "00110010",12644 => "00111000",12645 => "01011110",12646 => "01010111",12647 => "00000010",12648 => "10010110",12649 => "01111100",12650 => "01100101",12651 => "01101101",12652 => "00100000",12653 => "01001000",12654 => "01101010",12655 => "11010000",12656 => "11001000",12657 => "00000111",12658 => "01100111",12659 => "01101111",12660 => "10100011",12661 => "10101010",12662 => "10000101",12663 => "10000101",12664 => "11011001",12665 => "01101001",12666 => "11101010",12667 => "01101000",12668 => "10001111",12669 => "10101010",12670 => "00000111",12671 => "11000111",12672 => "11000111",12673 => "11101101",12674 => "00001000",12675 => "10111100",12676 => "01110010",12677 => "11100111",12678 => "00100111",12679 => "11111111",12680 => "10101111",12681 => "00111100",12682 => "11000001",12683 => "00010001",12684 => "01101011",12685 => "11101011",12686 => "00011101",12687 => "01010111",12688 => "11000010",12689 => "01001001",12690 => "10111001",12691 => "00010011",12692 => "00110011",12693 => "00011110",12694 => "11001101",12695 => "11000001",12696 => "10110111",12697 => "01011111",12698 => "01001110",12699 => "01100011",12700 => "11001101",12701 => "00101110",12702 => "10111110",12703 => "00110111",12704 => "11101010",12705 => "01011011",12706 => "00001110",12707 => "11111000",12708 => "00100100",12709 => "00000011",12710 => "10001010",12711 => "10010001",12712 => "01011100",12713 => "01110000",12714 => "00000001",12715 => "11101011",12716 => "00011101",12717 => "11011110",12718 => "11111111",12719 => "10011000",12720 => "11111010",12721 => "00111010",12722 => "10100001",12723 => "10001101",12724 => "11011001",12725 => "11100000",12726 => "01100101",12727 => "00011010",12728 => "10110010",12729 => "11110110",12730 => "10111011",12731 => "11100101",12732 => "00000010",12733 => "10011110",12734 => "11101000",12735 => "01111100",12736 => "00000101",12737 => "10100010",12738 => "10100000",12739 => "11101100",12740 => "11010101",12741 => "11101101",12742 => "10010101",12743 => "00111001",12744 => "11011000",12745 => "11011001",12746 => "00010100",12747 => "10010101",12748 => "01010100",12749 => "00010111",12750 => "10000110",12751 => "01110000",12752 => "11010001",12753 => "10000111",12754 => "01010100",12755 => "00010110",12756 => "01001100",12757 => "11000000",12758 => "01010010",12759 => "10110110",12760 => "10111000",12761 => "11010101",12762 => "11100101",12763 => "01100100",12764 => "11011000",12765 => "10010100",12766 => "00110110",12767 => "00010010",12768 => "11111110",12769 => "10000101",12770 => "00101100",12771 => "11000101",12772 => "11011101",12773 => "00001100",12774 => "10101110",12775 => "00010110",12776 => "01001110",12777 => "11011010",12778 => "10101101",12779 => "00011001",12780 => "10111111",12781 => "10011001",12782 => "00000111",12783 => "11100100",12784 => "01000000",12785 => "11110100",12786 => "10101011",12787 => "01101000",12788 => "10110101",12789 => "00100011",12790 => "00111111",12791 => "00000010",12792 => "01110000",12793 => "11101011",12794 => "00010001",12795 => "01111000",12796 => "00100100",12797 => "11111000",12798 => "10101110",12799 => "01111011",12800 => "11111001",12801 => "10101101",12802 => "11111011",12803 => "11011100",12804 => "11001111",12805 => "00101010",12806 => "00011101",12807 => "01101101",12808 => "11111100",12809 => "10101111",12810 => "11101000",12811 => "11011100",12812 => "01000100",12813 => "01110110",12814 => "11111111",12815 => "01100110",12816 => "11101111",12817 => "01000110",12818 => "00011011",12819 => "01011000",12820 => "11100010",12821 => "11110111",12822 => "11001001",12823 => "00110011",12824 => "11111111",12825 => "10010001",12826 => "01111101",12827 => "01000111",12828 => "01100011",12829 => "01000110",12830 => "11110001",12831 => "01010001",12832 => "10010010",12833 => "11111000",12834 => "00100000",12835 => "00000010",12836 => "00011001",12837 => "01110101",12838 => "01000010",12839 => "10000000",12840 => "11111111",12841 => "10001011",12842 => "01011001",12843 => "10000010",12844 => "10001110",12845 => "11110010",12846 => "01010111",12847 => "11111101",12848 => "00010000",12849 => "10000001",12850 => "10100001",12851 => "01100100",12852 => "01111111",12853 => "00111010",12854 => "01100010",12855 => "00010110",12856 => "10001011",12857 => "01011111",12858 => "00000100",12859 => "10011101",12860 => "10000001",12861 => "11011000",12862 => "11100111",12863 => "01100001",12864 => "01010010",12865 => "01101001",12866 => "11100001",12867 => "10101011",12868 => "11110111",12869 => "11001101",12870 => "11100101",12871 => "11100100",12872 => "01000100",12873 => "00100101",12874 => "11001010",12875 => "10010101",12876 => "01110011",12877 => "01101001",12878 => "01010010",12879 => "01011001",12880 => "10001010",12881 => "01111111",12882 => "00001001",12883 => "10110100",12884 => "11000010",12885 => "11001011",12886 => "10010000",12887 => "00011111",12888 => "11001101",12889 => "10011101",12890 => "01111001",12891 => "10010000",12892 => "10001111",12893 => "10000111",12894 => "01001110",12895 => "00101011",12896 => "10011010",12897 => "00100111",12898 => "01011111",12899 => "00111001",12900 => "00111101",12901 => "01110010",12902 => "00110100",12903 => "00101100",12904 => "00110000",12905 => "00111000",12906 => "00011011",12907 => "11011011",12908 => "10101101",12909 => "00011000",12910 => "11111011",12911 => "10100110",12912 => "00001000",12913 => "11111011",12914 => "01011010",12915 => "10100001",12916 => "01100001",12917 => "11110100",12918 => "00010101",12919 => "10000011",12920 => "11110001",12921 => "11000100",12922 => "11101100",12923 => "00100001",12924 => "00110101",12925 => "11000010",12926 => "10110010",12927 => "00110010",12928 => "01011010",12929 => "10000010",12930 => "10011000",12931 => "01101000",12932 => "11010000",12933 => "10110111",12934 => "00100010",12935 => "00000111",12936 => "11110000",12937 => "01001010",12938 => "01000111",12939 => "01011010",12940 => "11110101",12941 => "10011010",12942 => "01111011",12943 => "11101101",12944 => "10110110",12945 => "11100110",12946 => "01101001",12947 => "01111010",12948 => "00001001",12949 => "10010011",12950 => "01111000",12951 => "01100001",12952 => "00100011",12953 => "01011000",12954 => "11000110",12955 => "11001100",12956 => "01010000",12957 => "10011101",12958 => "11111001",12959 => "01100100",12960 => "01101111",12961 => "01101100",12962 => "01100010",12963 => "00111100",12964 => "10101100",12965 => "00000000",12966 => "01010011",12967 => "00111111",12968 => "00011001",12969 => "10110100",12970 => "11100001",12971 => "00100001",12972 => "01001000",12973 => "00001110",12974 => "11010110",12975 => "10110111",12976 => "11110110",12977 => "10101110",12978 => "10111100",12979 => "01101001",12980 => "11001110",12981 => "00011011",12982 => "00111110",12983 => "00001101",12984 => "11000100",12985 => "11011010",12986 => "00001010",12987 => "11011101",12988 => "10100100",12989 => "10101011",12990 => "01001010",12991 => "11000111",12992 => "01100001",12993 => "10110011",12994 => "00110001",12995 => "01110011",12996 => "00100000",12997 => "11110000",12998 => "00110100",12999 => "10111110",13000 => "11010001",13001 => "00001001",13002 => "10101111",13003 => "11000011",13004 => "11110110",13005 => "00110010",13006 => "01010110",13007 => "01111011",13008 => "10000010",13009 => "11011110",13010 => "10011001",13011 => "10000000",13012 => "11110011",13013 => "10000111",13014 => "00010100",13015 => "11001110",13016 => "11000110",13017 => "11011101",13018 => "01111111",13019 => "11011010",13020 => "00100111",13021 => "01100111",13022 => "11111110",13023 => "00001101",13024 => "01000011",13025 => "01010001",13026 => "11001000",13027 => "11111110",13028 => "01111011",13029 => "11001101",13030 => "01001101",13031 => "01000111",13032 => "11010001",13033 => "00111001",13034 => "01010011",13035 => "11000000",13036 => "11001000",13037 => "10111101",13038 => "10110000",13039 => "00000001",13040 => "00010111",13041 => "01010110",13042 => "11100101",13043 => "01001011",13044 => "00110100",13045 => "01011110",13046 => "11111101",13047 => "10001100",13048 => "00100001",13049 => "01101100",13050 => "10101010",13051 => "01110010",13052 => "10111111",13053 => "00010100",13054 => "10000001",13055 => "01101100",13056 => "01100011",13057 => "11101110",13058 => "11001001",13059 => "01101010",13060 => "00111000",13061 => "01111010",13062 => "11100011",13063 => "00101111",13064 => "11100110",13065 => "01000010",13066 => "00011111",13067 => "00101001",13068 => "00001111",13069 => "01111110",13070 => "10110000",13071 => "01010001",13072 => "10010110",13073 => "10001110",13074 => "11010111",13075 => "11100010",13076 => "00111010",13077 => "10101110",13078 => "01000100",13079 => "10111000",13080 => "01001000",13081 => "01101110",13082 => "10100000",13083 => "10010101",13084 => "11011111",13085 => "10011011",13086 => "10001101",13087 => "10001100",13088 => "01111100",13089 => "01111001",13090 => "00000001",13091 => "11001111",13092 => "11010001",13093 => "10001100",13094 => "10111100",13095 => "00100001",13096 => "11100000",13097 => "11111101",13098 => "00110111",13099 => "10010010",13100 => "01000000",13101 => "00000110",13102 => "00110101",13103 => "10000111",13104 => "10111000",13105 => "10101100",13106 => "11101010",13107 => "00000101",13108 => "01010001",13109 => "00000010",13110 => "01010001",13111 => "00100011",13112 => "11011111",13113 => "01110100",13114 => "10100110",13115 => "11101111",13116 => "00111011",13117 => "11011000",13118 => "11111111",13119 => "11100010",13120 => "00101000",13121 => "10110000",13122 => "11111101",13123 => "10100001",13124 => "11100100",13125 => "01010111",13126 => "10001000",13127 => "11110011",13128 => "00000110",13129 => "01110011",13130 => "10111111",13131 => "10000000",13132 => "00111110",13133 => "00110000",13134 => "01111010",13135 => "11000000",13136 => "00011100",13137 => "11011100",13138 => "01110011",13139 => "10011101",13140 => "11100101",13141 => "11111111",13142 => "11010000",13143 => "11110011",13144 => "01001101",13145 => "10001010",13146 => "11001010",13147 => "00111100",13148 => "11010110",13149 => "01101111",13150 => "00010000",13151 => "11101000",13152 => "10100110",13153 => "11001110",13154 => "10011110",13155 => "01110110",13156 => "00100011",13157 => "01101110",13158 => "00100100",13159 => "11001010",13160 => "11000111",13161 => "10101101",13162 => "11100011",13163 => "10010001",13164 => "11100111",13165 => "10001100",13166 => "11100100",13167 => "01111111",13168 => "00010100",13169 => "10110001",13170 => "11111011",13171 => "10000100",13172 => "01001100",13173 => "10111101",13174 => "11000111",13175 => "10000000",13176 => "01000101",13177 => "10011110",13178 => "10100010",13179 => "01111101",13180 => "10110000",13181 => "00000101",13182 => "11010101",13183 => "10100111",13184 => "11000001",13185 => "01110000",13186 => "00011101",13187 => "01011010",13188 => "10101001",13189 => "10101000",13190 => "01000111",13191 => "11101000",13192 => "00000001",13193 => "01011111",13194 => "01010010",13195 => "00011110",13196 => "11001010",13197 => "10010100",13198 => "10111011",13199 => "01110110",13200 => "10101010",13201 => "11011101",13202 => "11001001",13203 => "00100110",13204 => "11100001",13205 => "11000000",13206 => "11101010",13207 => "01111010",13208 => "00111100",13209 => "10101010",13210 => "00111111",13211 => "10000000",13212 => "01100101",13213 => "11111100",13214 => "01111111",13215 => "10110101",13216 => "01100001",13217 => "01110111",13218 => "11111001",13219 => "01010111",13220 => "00010010",13221 => "10010100",13222 => "11010010",13223 => "01010101",13224 => "11100110",13225 => "10101111",13226 => "10110000",13227 => "10001111",13228 => "10010010",13229 => "01100000",13230 => "00101110",13231 => "11101011",13232 => "11101001",13233 => "00101101",13234 => "00011100",13235 => "10110101",13236 => "01001000",13237 => "00111100",13238 => "00101111",13239 => "01100010",13240 => "10010110",13241 => "10100001",13242 => "00101101",13243 => "11010101",13244 => "11100101",13245 => "11001100",13246 => "01110111",13247 => "00101010",13248 => "01001001",13249 => "11000101",13250 => "11000011",13251 => "10111011",13252 => "10001110",13253 => "00001111",13254 => "11011110",13255 => "11111010",13256 => "00100111",13257 => "10111101",13258 => "10010000",13259 => "00001010",13260 => "01100110",13261 => "00011111",13262 => "00010001",13263 => "11100000",13264 => "01101011",13265 => "10000111",13266 => "01011111",13267 => "00010001",13268 => "11001001",13269 => "11010100",13270 => "00100010",13271 => "01100101",13272 => "01111011",13273 => "00100011",13274 => "11101010",13275 => "10011010",13276 => "00011110",13277 => "00100001",13278 => "10110001",13279 => "10100101",13280 => "01011110",13281 => "00101100",13282 => "10110101",13283 => "11001001",13284 => "10010110",13285 => "01000110",13286 => "10001101",13287 => "11110111",13288 => "11010000",13289 => "11101011",13290 => "00010011",13291 => "01001111",13292 => "00010010",13293 => "11111010",13294 => "01011110",13295 => "10101010",13296 => "10001001",13297 => "11110010",13298 => "11000101",13299 => "11101001",13300 => "10001101",13301 => "01001000",13302 => "00001111",13303 => "10100010",13304 => "11111111",13305 => "01110011",13306 => "11111100",13307 => "11000011",13308 => "11000011",13309 => "01101101",13310 => "10100111",13311 => "10100011",13312 => "01001110",13313 => "10001101",13314 => "00000000",13315 => "11100111",13316 => "01001101",13317 => "01111101",13318 => "10000001",13319 => "01100001",13320 => "10010100",13321 => "11100100",13322 => "11010010",13323 => "11001100",13324 => "11011000",13325 => "01100001",13326 => "10010010",13327 => "01111100",13328 => "00010011",13329 => "00011111",13330 => "10011110",13331 => "11001010",13332 => "11011111",13333 => "10110001",13334 => "00000101",13335 => "00100101",13336 => "00001001",13337 => "11000001",13338 => "01111110",13339 => "01100101",13340 => "10101000",13341 => "11000110",13342 => "01101110",13343 => "11100111",13344 => "10010111",13345 => "10010010",13346 => "10111011",13347 => "11001011",13348 => "00010010",13349 => "00010000",13350 => "11000000",13351 => "01001010",13352 => "11101010",13353 => "11001011",13354 => "10011111",13355 => "11101110",13356 => "10011110",13357 => "01100110",13358 => "11000011",13359 => "01000001",13360 => "10011000",13361 => "00110011",13362 => "11100111",13363 => "11100111",13364 => "10010100",13365 => "10111111",13366 => "01101011",13367 => "01111100",13368 => "10011110",13369 => "01110000",13370 => "00111111",13371 => "11101001",13372 => "01000010",13373 => "00110011",13374 => "10000011",13375 => "11101101",13376 => "00110011",13377 => "11101010",13378 => "10000010",13379 => "01100001",13380 => "11101100",13381 => "10011001",13382 => "10110110",13383 => "11100101",13384 => "01111110",13385 => "10100111",13386 => "01011111",13387 => "10011101",13388 => "00001110",13389 => "01010001",13390 => "10111101",13391 => "11101101",13392 => "11111110",13393 => "11111001",13394 => "00100100",13395 => "00000011",13396 => "01010110",13397 => "01010111",13398 => "10111110",13399 => "01111110",13400 => "01010111",13401 => "01001010",13402 => "00101111",13403 => "11001100",13404 => "11101000",13405 => "11101111",13406 => "10011010",13407 => "10011101",13408 => "01010010",13409 => "10110110",13410 => "00111010",13411 => "11111110",13412 => "11001111",13413 => "11111101",13414 => "11010001",13415 => "01110101",13416 => "00011100",13417 => "00001111",13418 => "10111100",13419 => "00010100",13420 => "11011100",13421 => "10010111",13422 => "01000101",13423 => "10010011",13424 => "01010110",13425 => "11100111",13426 => "00000001",13427 => "01110110",13428 => "10100110",13429 => "00001011",13430 => "00011111",13431 => "00101100",13432 => "00001011",13433 => "10011000",13434 => "10110000",13435 => "11010000",13436 => "00010011",13437 => "01000010",13438 => "01100111",13439 => "10011011",13440 => "10011000",13441 => "01110011",13442 => "01100101",13443 => "00001100",13444 => "00110011",13445 => "00000100",13446 => "00010111",13447 => "01010101",13448 => "00010100",13449 => "10000110",13450 => "11010111",13451 => "00110010",13452 => "11100011",13453 => "11111000",13454 => "00101010",13455 => "10110001",13456 => "01010000",13457 => "00110101",13458 => "01101101",13459 => "11111001",13460 => "01001011",13461 => "01101111",13462 => "00000010",13463 => "11000100",13464 => "00111111",13465 => "01011001",13466 => "01011010",13467 => "01111111",13468 => "01110000",13469 => "01100111",13470 => "00011010",13471 => "01100011",13472 => "11001110",13473 => "01000110",13474 => "00100010",13475 => "10100010",13476 => "11001111",13477 => "00001111",13478 => "01110111",13479 => "11001101",13480 => "11011101",13481 => "00101000",13482 => "01111111",13483 => "00110000",13484 => "10101001",13485 => "10101101",13486 => "01011110",13487 => "00111001",13488 => "10010110",13489 => "11101011",13490 => "00111110",13491 => "10001101",13492 => "00110011",13493 => "00011101",13494 => "10111011",13495 => "01101011",13496 => "10010111",13497 => "10010111",13498 => "11110100",13499 => "01010011",13500 => "01111001",13501 => "11101101",13502 => "10111000",13503 => "01011111",13504 => "00101100",13505 => "00101010",13506 => "11000011",13507 => "01000100",13508 => "00110000",13509 => "00101001",13510 => "10000000",13511 => "10110101",13512 => "00001000",13513 => "11101101",13514 => "11010110",13515 => "10011101",13516 => "01101100",13517 => "11100110",13518 => "11111011",13519 => "00011110",13520 => "01010101",13521 => "00011000",13522 => "10010111",13523 => "10100100",13524 => "00011011",13525 => "01000101",13526 => "00011110",13527 => "11010110",13528 => "00111110",13529 => "10001111",13530 => "10110000",13531 => "01010000",13532 => "01000101",13533 => "01010000",13534 => "10111101",13535 => "01001010",13536 => "01001000",13537 => "11011010",13538 => "11101111",13539 => "01000101",13540 => "11011001",13541 => "00000010",13542 => "10101000",13543 => "10011011",13544 => "01111111",13545 => "01101000",13546 => "10010000",13547 => "00011100",13548 => "11111111",13549 => "10010101",13550 => "01110000",13551 => "11000101",13552 => "00110110",13553 => "11011101",13554 => "10000111",13555 => "10100011",13556 => "01010111",13557 => "11111111",13558 => "00101110",13559 => "10011011",13560 => "11001011",13561 => "11101001",13562 => "00011111",13563 => "11110100",13564 => "00101011",13565 => "10100001",13566 => "01100101",13567 => "11000110",13568 => "00000100",13569 => "10000011",13570 => "01001100",13571 => "10010001",13572 => "01010001",13573 => "11011110",13574 => "10101001",13575 => "01001001",13576 => "11111010",13577 => "10010001",13578 => "01111100",13579 => "11000110",13580 => "01101010",13581 => "11010001",13582 => "10111110",13583 => "10111011",13584 => "00000001",13585 => "11011011",13586 => "01101111",13587 => "11100101",13588 => "11010001",13589 => "10001010",13590 => "01110100",13591 => "01001001",13592 => "10101111",13593 => "11000000",13594 => "01110110",13595 => "11010110",13596 => "10110111",13597 => "10100010",13598 => "10101110",13599 => "00000001",13600 => "11010000",13601 => "00100101",13602 => "10110000",13603 => "11101001",13604 => "11100001",13605 => "11011001",13606 => "10111011",13607 => "01001111",13608 => "00110010",13609 => "01010011",13610 => "01100101",13611 => "01011101",13612 => "01010001",13613 => "10110100",13614 => "10000001",13615 => "11000001",13616 => "11110001",13617 => "01101011",13618 => "10010101",13619 => "10011000",13620 => "10011001",13621 => "01001100",13622 => "11101011",13623 => "10001011",13624 => "10111010",13625 => "10000000",13626 => "10111010",13627 => "10110111",13628 => "01000111",13629 => "00011011",13630 => "00001001",13631 => "00111000",13632 => "10001110",13633 => "11001100",13634 => "10100100",13635 => "10111111",13636 => "00001101",13637 => "01000111",13638 => "01001011",13639 => "11011100",13640 => "01110000",13641 => "10101010",13642 => "01010100",13643 => "11010011",13644 => "01001000",13645 => "10111000",13646 => "11111110",13647 => "11110011",13648 => "11100000",13649 => "11001101",13650 => "11100010",13651 => "01101101",13652 => "01110010",13653 => "01110001",13654 => "11100101",13655 => "11001010",13656 => "01110101",13657 => "10110011",13658 => "11010111",13659 => "00100110",13660 => "00100000",13661 => "11101001",13662 => "11010011",13663 => "11100001",13664 => "01110001",13665 => "11111000",13666 => "01010100",13667 => "11010011",13668 => "01101000",13669 => "10110111",13670 => "00011010",13671 => "01011110",13672 => "00011110",13673 => "00010011",13674 => "10111100",13675 => "11000000",13676 => "01001011",13677 => "11111100",13678 => "01010000",13679 => "01100000",13680 => "01110111",13681 => "10100010",13682 => "11100011",13683 => "00111110",13684 => "10010011",13685 => "01010011",13686 => "00111110",13687 => "11011000",13688 => "01111110",13689 => "11010010",13690 => "01101101",13691 => "01101010",13692 => "10001110",13693 => "11011011",13694 => "10010001",13695 => "11100010",13696 => "10011010",13697 => "00011000",13698 => "00110101",13699 => "10110111",13700 => "10100010",13701 => "01001111",13702 => "01110100",13703 => "11010010",13704 => "10001000",13705 => "11001100",13706 => "00001010",13707 => "00101101",13708 => "10000011",13709 => "11011100",13710 => "00101110",13711 => "01000100",13712 => "00001011",13713 => "01011100",13714 => "00100010",13715 => "10100000",13716 => "00011110",13717 => "10010111",13718 => "10010101",13719 => "11100001",13720 => "01110111",13721 => "00101101",13722 => "10010010",13723 => "00111011",13724 => "10110110",13725 => "01111111",13726 => "00101101",13727 => "10110101",13728 => "01011001",13729 => "01011010",13730 => "10000111",13731 => "11011110",13732 => "01010010",13733 => "00100011",13734 => "11100000",13735 => "01011001",13736 => "11101110",13737 => "11001101",13738 => "01111001",13739 => "11000010",13740 => "00001010",13741 => "11111100",13742 => "11000000",13743 => "01011110",13744 => "01111100",13745 => "00110101",13746 => "01011100",13747 => "01111011",13748 => "01100000",13749 => "01011101",13750 => "01010100",13751 => "11010010",13752 => "00101000",13753 => "10000110",13754 => "01011111",13755 => "10111100",13756 => "00010011",13757 => "10011010",13758 => "10000001",13759 => "01001101",13760 => "00101100",13761 => "00010101",13762 => "00001011",13763 => "10111000",13764 => "10111110",13765 => "11110110",13766 => "01100110",13767 => "11111001",13768 => "01101111",13769 => "10010110",13770 => "00100101",13771 => "11101100",13772 => "11001011",13773 => "10011011",13774 => "11000100",13775 => "01011010",13776 => "01011101",13777 => "00011011",13778 => "00111111",13779 => "11101111",13780 => "10001011",13781 => "00001000",13782 => "00110000",13783 => "11100111",13784 => "00110111",13785 => "11011000",13786 => "11101111",13787 => "11101001",13788 => "01100010",13789 => "01000110",13790 => "00100101",13791 => "01011100",13792 => "11011101",13793 => "10100100",13794 => "01100111",13795 => "11110000",13796 => "01000111",13797 => "01010010",13798 => "00010100",13799 => "01101110",13800 => "01110000",13801 => "01111111",13802 => "11100000",13803 => "10000111",13804 => "00111110",13805 => "01001101",13806 => "10000111",13807 => "11111010",13808 => "01010011",13809 => "10011011",13810 => "10010101",13811 => "10100010",13812 => "00111011",13813 => "11010011",13814 => "10001000",13815 => "01111110",13816 => "11101101",13817 => "01010011",13818 => "01101000",13819 => "00101000",13820 => "10000110",13821 => "10011011",13822 => "01100010",13823 => "10110010",13824 => "00101110",13825 => "10111101",13826 => "10111111",13827 => "00100100",13828 => "00101001",13829 => "10111001",13830 => "00101001",13831 => "00000000",13832 => "01001011",13833 => "10001000",13834 => "10111010",13835 => "00000111",13836 => "11100010",13837 => "00011000",13838 => "10101111",13839 => "10001001",13840 => "00110000",13841 => "00110111",13842 => "00011110",13843 => "11011101",13844 => "11100000",13845 => "01111110",13846 => "11010010",13847 => "01010010",13848 => "00000100",13849 => "11110101",13850 => "11100111",13851 => "10010100",13852 => "00011110",13853 => "00100000",13854 => "00111000",13855 => "01111001",13856 => "11110100",13857 => "00101000",13858 => "10010111",13859 => "00101011",13860 => "11100000",13861 => "10001111",13862 => "10000110",13863 => "00000101",13864 => "11111001",13865 => "01101101",13866 => "11101011",13867 => "00011111",13868 => "01011100",13869 => "10001110",13870 => "00011101",13871 => "10100110",13872 => "00110100",13873 => "11010110",13874 => "11101011",13875 => "10110101",13876 => "01101001",13877 => "11100111",13878 => "01100001",13879 => "01011010",13880 => "10101011",13881 => "10100110",13882 => "00011011",13883 => "01000011",13884 => "00011101",13885 => "11010111",13886 => "11100100",13887 => "01011101",13888 => "01001110",13889 => "10110011",13890 => "10100110",13891 => "10010100",13892 => "11001000",13893 => "10011110",13894 => "00000011",13895 => "01110000",13896 => "00101001",13897 => "00011111",13898 => "10100111",13899 => "10111000",13900 => "11010111",13901 => "01111101",13902 => "11001101",13903 => "10000011",13904 => "11010101",13905 => "01111100",13906 => "01000100",13907 => "10011101",13908 => "00111000",13909 => "10001000",13910 => "01001101",13911 => "01001101",13912 => "01111101",13913 => "11001111",13914 => "00100110",13915 => "00111110",13916 => "01100100",13917 => "11011111",13918 => "10001000",13919 => "00101010",13920 => "11111011",13921 => "10011100",13922 => "10010110",13923 => "01101101",13924 => "00001000",13925 => "01110110",13926 => "00011000",13927 => "00100101",13928 => "11011001",13929 => "00110011",13930 => "11100101",13931 => "11101000",13932 => "01101010",13933 => "00110011",13934 => "11000011",13935 => "11100110",13936 => "10110011",13937 => "11110000",13938 => "10000101",13939 => "01110110",13940 => "11100111",13941 => "00001010",13942 => "11010111",13943 => "01010011",13944 => "01001010",13945 => "01100101",13946 => "10000100",13947 => "11000001",13948 => "10100000",13949 => "00100100",13950 => "00000111",13951 => "01111001",13952 => "10000100",13953 => "10110001",13954 => "10011011",13955 => "00101111",13956 => "11010001",13957 => "00111010",13958 => "01000101",13959 => "01011101",13960 => "10110110",13961 => "11110101",13962 => "11100111",13963 => "01001001",13964 => "00011111",13965 => "11000001",13966 => "11000001",13967 => "00110000",13968 => "01001001",13969 => "00011101",13970 => "11100000",13971 => "10111000",13972 => "01101110",13973 => "10110001",13974 => "01100000",13975 => "11100010",13976 => "01010011",13977 => "00110010",13978 => "01101101",13979 => "10010110",13980 => "11000110",13981 => "00000100",13982 => "01001001",13983 => "11000000",13984 => "10100111",13985 => "10101001",13986 => "10101010",13987 => "10010001",13988 => "10001100",13989 => "01111010",13990 => "01101011",13991 => "01101110",13992 => "01011111",13993 => "00011001",13994 => "10111000",13995 => "10110000",13996 => "11100010",13997 => "11011011",13998 => "01100100",13999 => "11111001",14000 => "00101010",14001 => "11011011",14002 => "11101101",14003 => "10100010",14004 => "11101110",14005 => "01001010",14006 => "10000111",14007 => "10010011",14008 => "01110101",14009 => "00000110",14010 => "11101110",14011 => "01001001",14012 => "11001000",14013 => "10101101",14014 => "10000101",14015 => "00011001",14016 => "00001101",14017 => "00101100",14018 => "01001111",14019 => "11110001",14020 => "00101110",14021 => "01011110",14022 => "11110100",14023 => "00101110",14024 => "11010100",14025 => "10011011",14026 => "11101100",14027 => "01010110",14028 => "01111011",14029 => "00100111",14030 => "00010010",14031 => "10001111",14032 => "11000000",14033 => "01010100",14034 => "01111010",14035 => "01001100",14036 => "01011011",14037 => "11111101",14038 => "01001001",14039 => "00100110",14040 => "00000001",14041 => "00011011",14042 => "11110110",14043 => "10001010",14044 => "00010011",14045 => "10011011",14046 => "00111111",14047 => "00101100",14048 => "10000000",14049 => "11000100",14050 => "10000011",14051 => "10011100",14052 => "11101100",14053 => "01001100",14054 => "10101011",14055 => "01110101",14056 => "01111011",14057 => "01001110",14058 => "10100100",14059 => "11011111",14060 => "00000000",14061 => "11011010",14062 => "00000001",14063 => "01010001",14064 => "00110111",14065 => "00101101",14066 => "10001001",14067 => "01111100",14068 => "10111000",14069 => "10011101",14070 => "00100011",14071 => "11001010",14072 => "10111110",14073 => "01111001",14074 => "00001100",14075 => "10010110",14076 => "11010010",14077 => "11001000",14078 => "10111001",14079 => "00000010",14080 => "01001001",14081 => "10001000",14082 => "10001011",14083 => "00111100",14084 => "10001010",14085 => "01000101",14086 => "11110110",14087 => "10001100",14088 => "01111010",14089 => "10111110",14090 => "01000000",14091 => "01110101",14092 => "00011110",14093 => "11111011",14094 => "11101001",14095 => "01101000",14096 => "01100001",14097 => "01001011",14098 => "10111001",14099 => "01001111",14100 => "10011000",14101 => "10010011",14102 => "00010010",14103 => "00001010",14104 => "11101001",14105 => "00010011",14106 => "00110001",14107 => "01000010",14108 => "10000100",14109 => "00101010",14110 => "11110110",14111 => "11001000",14112 => "00011100",14113 => "11001111",14114 => "00100001",14115 => "11111011",14116 => "01010111",14117 => "11100000",14118 => "10111110",14119 => "11100011",14120 => "00010100",14121 => "01101101",14122 => "00100111",14123 => "01101001",14124 => "11100000",14125 => "01001101",14126 => "11011001",14127 => "01111001",14128 => "10110110",14129 => "00011101",14130 => "11110001",14131 => "01000000",14132 => "01100111",14133 => "11111111",14134 => "00111000",14135 => "01100010",14136 => "11010000",14137 => "10000110",14138 => "10101001",14139 => "11110010",14140 => "00010100",14141 => "10110011",14142 => "01010111",14143 => "10010101",14144 => "00001111",14145 => "00001000",14146 => "01110111",14147 => "10110111",14148 => "01111000",14149 => "10101000",14150 => "10110010",14151 => "11101100",14152 => "01001111",14153 => "11000011",14154 => "01001010",14155 => "11111101",14156 => "01010010",14157 => "10100111",14158 => "01111000",14159 => "01110100",14160 => "10111011",14161 => "00001101",14162 => "11100111",14163 => "00010001",14164 => "11010010",14165 => "11101101",14166 => "10110011",14167 => "00010100",14168 => "00010100",14169 => "10100001",14170 => "11011100",14171 => "10100100",14172 => "00011000",14173 => "10111110",14174 => "11111110",14175 => "10100010",14176 => "00011001",14177 => "11011101",14178 => "10011000",14179 => "01000101",14180 => "00011101",14181 => "00001010",14182 => "11000111",14183 => "00010010",14184 => "11001110",14185 => "00101001",14186 => "00110110",14187 => "01111111",14188 => "11100011",14189 => "01100001",14190 => "00000110",14191 => "01000001",14192 => "11000001",14193 => "00011001",14194 => "10110001",14195 => "11111010",14196 => "00001000",14197 => "01101011",14198 => "01110000",14199 => "00011100",14200 => "00110111",14201 => "10001000",14202 => "01110111",14203 => "11010001",14204 => "11000101",14205 => "00101000",14206 => "01101001",14207 => "10110011",14208 => "10110110",14209 => "00100111",14210 => "00111110",14211 => "11111111",14212 => "00011111",14213 => "00000011",14214 => "01000001",14215 => "01110011",14216 => "10100000",14217 => "00010010",14218 => "00001100",14219 => "00010111",14220 => "01001100",14221 => "10111100",14222 => "11110111",14223 => "11001010",14224 => "10000011",14225 => "10100110",14226 => "00011000",14227 => "00100001",14228 => "11001010",14229 => "11101010",14230 => "00100100",14231 => "01101101",14232 => "01111001",14233 => "11110101",14234 => "01010111",14235 => "10000101",14236 => "10110001",14237 => "10000100",14238 => "00100111",14239 => "10101100",14240 => "00000111",14241 => "01010110",14242 => "00110000",14243 => "11011110",14244 => "10011111",14245 => "01011001",14246 => "11110000",14247 => "00111001",14248 => "00001100",14249 => "11011001",14250 => "00101101",14251 => "01101100",14252 => "10010111",14253 => "11111001",14254 => "00010100",14255 => "00001001",14256 => "00001011",14257 => "01010010",14258 => "01111101",14259 => "10101111",14260 => "10111010",14261 => "11110110",14262 => "10011000",14263 => "11011010",14264 => "01111110",14265 => "01100111",14266 => "00000011",14267 => "11001011",14268 => "01101011",14269 => "11000101",14270 => "10111101",14271 => "01100011",14272 => "00101010",14273 => "10110010",14274 => "01010010",14275 => "11101010",14276 => "00110001",14277 => "10111100",14278 => "11111000",14279 => "00101101",14280 => "10101010",14281 => "11111110",14282 => "01111001",14283 => "11001011",14284 => "11101000",14285 => "00000001",14286 => "00101011",14287 => "10100000",14288 => "11001100",14289 => "11011101",14290 => "00111111",14291 => "11011000",14292 => "00000111",14293 => "11101010",14294 => "10111010",14295 => "11011101",14296 => "01101001",14297 => "11111000",14298 => "00001010",14299 => "00110110",14300 => "00111110",14301 => "00100101",14302 => "01011001",14303 => "01110001",14304 => "11100001",14305 => "10010001",14306 => "11101100",14307 => "01101001",14308 => "00000000",14309 => "01011101",14310 => "01000111",14311 => "00011010",14312 => "00001101",14313 => "11100001",14314 => "11101000",14315 => "10100100",14316 => "11111001",14317 => "11111010",14318 => "01110010",14319 => "10001000",14320 => "11000100",14321 => "00100011",14322 => "10000101",14323 => "11011101",14324 => "10100001",14325 => "00000000",14326 => "10010111",14327 => "10100001",14328 => "10110001",14329 => "00001001",14330 => "00000111",14331 => "00010000",14332 => "11000000",14333 => "11010100",14334 => "10101001",14335 => "01000100",14336 => "01101001",14337 => "00101010",14338 => "11111100",14339 => "11111010",14340 => "11000001",14341 => "10100011",14342 => "11111010",14343 => "11010111",14344 => "10100100",14345 => "00000101",14346 => "00110001",14347 => "11110001",14348 => "11010101",14349 => "00011000",14350 => "00001000",14351 => "10100100",14352 => "11111110",14353 => "11000110",14354 => "11101000",14355 => "01111100",14356 => "11111111",14357 => "10100110",14358 => "10101110",14359 => "01001111",14360 => "01010011",14361 => "00011101",14362 => "10100010",14363 => "11010101",14364 => "00001011",14365 => "10011011",14366 => "00011101",14367 => "00100010",14368 => "00001011",14369 => "01110110",14370 => "10110101",14371 => "00110001",14372 => "11001011",14373 => "01101100",14374 => "10101011",14375 => "10010001",14376 => "00100110",14377 => "00010000",14378 => "01111110",14379 => "11000111",14380 => "10011001",14381 => "11110001",14382 => "10000111",14383 => "00001100",14384 => "11110000",14385 => "11001000",14386 => "10111000",14387 => "10101000",14388 => "00101111",14389 => "11101001",14390 => "00110110",14391 => "00011011",14392 => "11011110",14393 => "11010101",14394 => "11110111",14395 => "10110010",14396 => "10100001",14397 => "11011110",14398 => "00111010",14399 => "10010001",14400 => "10101111",14401 => "11111011",14402 => "10001001",14403 => "11111100",14404 => "00101101",14405 => "11000100",14406 => "01001111",14407 => "11000101",14408 => "11110011",14409 => "00110110",14410 => "11010010",14411 => "00011100",14412 => "00100101",14413 => "11001110",14414 => "10010101",14415 => "00101101",14416 => "10100000",14417 => "10000100",14418 => "10110000",14419 => "01111001",14420 => "11101001",14421 => "10010001",14422 => "00011000",14423 => "01110110",14424 => "10110011",14425 => "10011111",14426 => "10000010",14427 => "01100101",14428 => "01101100",14429 => "10001011",14430 => "11111100",14431 => "00000100",14432 => "01100001",14433 => "11100101",14434 => "10101001",14435 => "10111101",14436 => "10001010",14437 => "00000100",14438 => "00001110",14439 => "01101110",14440 => "01101000",14441 => "10101001",14442 => "11100100",14443 => "11101101",14444 => "10111111",14445 => "10010100",14446 => "00000110",14447 => "11100010",14448 => "11011110",14449 => "11110011",14450 => "00110010",14451 => "00110001",14452 => "00010111",14453 => "10010001",14454 => "10101111",14455 => "00100000",14456 => "11100110",14457 => "11100001",14458 => "11011111",14459 => "11110010",14460 => "01011000",14461 => "10111011",14462 => "01111111",14463 => "11001000",14464 => "01110001",14465 => "01010110",14466 => "00111000",14467 => "01000101",14468 => "01000110",14469 => "01111100",14470 => "01010001",14471 => "10001100",14472 => "10110111",14473 => "01011111",14474 => "11111100",14475 => "11110101",14476 => "10011100",14477 => "00111111",14478 => "00000001",14479 => "00010001",14480 => "10111011",14481 => "01100101",14482 => "01100101",14483 => "10100100",14484 => "11010111",14485 => "00011111",14486 => "10101110",14487 => "01101000",14488 => "11001100",14489 => "00100111",14490 => "00011101",14491 => "00010101",14492 => "00011110",14493 => "00111110",14494 => "00111001",14495 => "10000011",14496 => "11000110",14497 => "01101001",14498 => "11110111",14499 => "00110011",14500 => "11000011",14501 => "10010011",14502 => "10100110",14503 => "10001101",14504 => "00011011",14505 => "01111010",14506 => "11100100",14507 => "10111011",14508 => "10010001",14509 => "01001011",14510 => "00111010",14511 => "00110111",14512 => "11111111",14513 => "00111101",14514 => "10001100",14515 => "10110000",14516 => "01010100",14517 => "10101100",14518 => "11010011",14519 => "10101011",14520 => "00111100",14521 => "10000111",14522 => "11110110",14523 => "00011111",14524 => "01001011",14525 => "00011100",14526 => "01100111",14527 => "11111001",14528 => "00101111",14529 => "01110100",14530 => "10101110",14531 => "00110000",14532 => "11100011",14533 => "00110010",14534 => "10001001",14535 => "00011000",14536 => "10001100",14537 => "11111011",14538 => "10111100",14539 => "00101101",14540 => "11101100",14541 => "01000101",14542 => "00110011",14543 => "01111011",14544 => "00100010",14545 => "11101011",14546 => "10011100",14547 => "01001101",14548 => "00011101",14549 => "10001001",14550 => "10101000",14551 => "11101010",14552 => "01100110",14553 => "01101100",14554 => "10100111",14555 => "10001111",14556 => "01010011",14557 => "01111111",14558 => "10110100",14559 => "00111100",14560 => "11100110",14561 => "00011111",14562 => "00111000",14563 => "00010000",14564 => "01000101",14565 => "00100101",14566 => "10101100",14567 => "10000101",14568 => "00111101",14569 => "00011001",14570 => "01101011",14571 => "11101100",14572 => "11000110",14573 => "01100010",14574 => "11010100",14575 => "01001010",14576 => "01000110",14577 => "11100011",14578 => "00001111",14579 => "01111000",14580 => "01110111",14581 => "10110001",14582 => "01001011",14583 => "10110101",14584 => "00000110",14585 => "00111100",14586 => "01011000",14587 => "01110000",14588 => "00101011",14589 => "10000101",14590 => "00010001",14591 => "00110100",14592 => "10100011",14593 => "10110101",14594 => "01001000",14595 => "01100101",14596 => "11101100",14597 => "01000100",14598 => "00001010",14599 => "11010110",14600 => "10100010",14601 => "01100010",14602 => "10100100",14603 => "10100010",14604 => "10110000",14605 => "11010001",14606 => "01001010",14607 => "11111110",14608 => "11101110",14609 => "10111111",14610 => "00010001",14611 => "00000001",14612 => "00100101",14613 => "11110011",14614 => "10110000",14615 => "01101100",14616 => "00011101",14617 => "11100100",14618 => "10010110",14619 => "01011111",14620 => "10001100",14621 => "01110100",14622 => "11111100",14623 => "01101101",14624 => "11001010",14625 => "00100101",14626 => "10010110",14627 => "01110110",14628 => "11010100",14629 => "11010100",14630 => "11111100",14631 => "11000000",14632 => "01011111",14633 => "11110000",14634 => "00111000",14635 => "10010001",14636 => "10111011",14637 => "01010000",14638 => "11110010",14639 => "11101011",14640 => "00111010",14641 => "00110101",14642 => "01110111",14643 => "11110101",14644 => "01001000",14645 => "01001111",14646 => "01000111",14647 => "01000100",14648 => "11010011",14649 => "10001110",14650 => "10100000",14651 => "00101110",14652 => "01101011",14653 => "01100001",14654 => "10001011",14655 => "10001010",14656 => "10001010",14657 => "10111101",14658 => "01000000",14659 => "10001110",14660 => "01011000",14661 => "01010101",14662 => "01110000",14663 => "00110100",14664 => "01001010",14665 => "11111100",14666 => "00001000",14667 => "01000100",14668 => "01111010",14669 => "01010010",14670 => "00111111",14671 => "00011100",14672 => "00011001",14673 => "10111010",14674 => "11011001",14675 => "00110110",14676 => "10100000",14677 => "01010001",14678 => "00000010",14679 => "11110011",14680 => "11110001",14681 => "10111100",14682 => "11011111",14683 => "00001010",14684 => "10111010",14685 => "10010010",14686 => "01111000",14687 => "01011000",14688 => "11111011",14689 => "01100000",14690 => "10111100",14691 => "00110110",14692 => "10100100",14693 => "11001101",14694 => "10010110",14695 => "11110010",14696 => "10111111",14697 => "00110011",14698 => "00101110",14699 => "11000011",14700 => "00001001",14701 => "11101101",14702 => "00001001",14703 => "01011000",14704 => "00101011",14705 => "01001100",14706 => "11010111",14707 => "01111101",14708 => "00100010",14709 => "01111001",14710 => "00100000",14711 => "01110010",14712 => "10010000",14713 => "01111100",14714 => "10111001",14715 => "00110000",14716 => "10001001",14717 => "01111001",14718 => "11110111",14719 => "10101110",14720 => "11100100",14721 => "00010000",14722 => "00110111",14723 => "01001010",14724 => "10011100",14725 => "10110110",14726 => "11101010",14727 => "10011101",14728 => "10010010",14729 => "00110110",14730 => "11001101",14731 => "11001101",14732 => "11000100",14733 => "01010111",14734 => "11100100",14735 => "00001110",14736 => "11011110",14737 => "10000011",14738 => "01001001",14739 => "11001110",14740 => "10001111",14741 => "01110100",14742 => "11110101",14743 => "10110101",14744 => "11101001",14745 => "11100110",14746 => "00110001",14747 => "11101000",14748 => "01011011",14749 => "11101111",14750 => "10011010",14751 => "00100101",14752 => "10100000",14753 => "10101001",14754 => "00111010",14755 => "01110101",14756 => "00000001",14757 => "00110011",14758 => "11100111",14759 => "01110001",14760 => "00111010",14761 => "11111111",14762 => "00001110",14763 => "10011010",14764 => "11011011",14765 => "11111111",14766 => "10100010",14767 => "00011110",14768 => "10101101",14769 => "11001001",14770 => "00000101",14771 => "00110110",14772 => "00010100",14773 => "10010001",14774 => "01000011",14775 => "01111010",14776 => "11000000",14777 => "10001010",14778 => "11110100",14779 => "01001011",14780 => "10110100",14781 => "11101000",14782 => "10101110",14783 => "10110101",14784 => "01010111",14785 => "11010101",14786 => "11110110",14787 => "00110111",14788 => "10001111",14789 => "01011101",14790 => "00101101",14791 => "01101111",14792 => "11111100",14793 => "00101110",14794 => "00110110",14795 => "11011110",14796 => "00101111",14797 => "11011110",14798 => "10010001",14799 => "01111001",14800 => "10110001",14801 => "01010100",14802 => "11101011",14803 => "11001011",14804 => "01011111",14805 => "01110001",14806 => "00100111",14807 => "10111011",14808 => "01000100",14809 => "00100000",14810 => "10011000",14811 => "10100100",14812 => "10100110",14813 => "11001001",14814 => "10000000",14815 => "00011110",14816 => "10010111",14817 => "10101111",14818 => "00110010",14819 => "11010011",14820 => "00111111",14821 => "00111001",14822 => "10101101",14823 => "10110110",14824 => "00001100",14825 => "10000001",14826 => "11100000",14827 => "11010101",14828 => "10111110",14829 => "11011101",14830 => "10100001",14831 => "00110101",14832 => "01010000",14833 => "00110101",14834 => "01111000",14835 => "01010100",14836 => "11111111",14837 => "00000011",14838 => "10011111",14839 => "01100101",14840 => "11000111",14841 => "00000011",14842 => "00011000",14843 => "01000001",14844 => "00000000",14845 => "11100001",14846 => "11011001",14847 => "01000101",14848 => "00100010",14849 => "00100100",14850 => "00100101",14851 => "11001111",14852 => "01110111",14853 => "01010001",14854 => "10001010",14855 => "10101110",14856 => "11001111",14857 => "11110011",14858 => "11000000",14859 => "11010111",14860 => "01110001",14861 => "01101101",14862 => "01000111",14863 => "00011111",14864 => "10011101",14865 => "01000100",14866 => "00010111",14867 => "00101111",14868 => "00001110",14869 => "11010010",14870 => "10010000",14871 => "11011011",14872 => "00110110",14873 => "11010110",14874 => "11011010",14875 => "10000111",14876 => "01010001",14877 => "01011110",14878 => "10101111",14879 => "00110011",14880 => "11110100",14881 => "10001011",14882 => "10011110",14883 => "00101011",14884 => "01010001",14885 => "00001011",14886 => "10001010",14887 => "11110000",14888 => "11100011",14889 => "00011111",14890 => "10011000",14891 => "00101111",14892 => "00111101",14893 => "01100001",14894 => "01110111",14895 => "00100100",14896 => "10110010",14897 => "10000011",14898 => "10110000",14899 => "01111111",14900 => "00011100",14901 => "00010011",14902 => "11101110",14903 => "00000011",14904 => "00100110",14905 => "01101111",14906 => "01011101",14907 => "10010000",14908 => "11000011",14909 => "00101000",14910 => "11000010",14911 => "11111101",14912 => "00101111",14913 => "01101100",14914 => "11000001",14915 => "10110101",14916 => "00110101",14917 => "00111111",14918 => "11111111",14919 => "01101001",14920 => "01010010",14921 => "10111101",14922 => "01001111",14923 => "10111110",14924 => "10011100",14925 => "10101000",14926 => "00000001",14927 => "01011010",14928 => "00011110",14929 => "10001011",14930 => "11001100",14931 => "00101101",14932 => "00111111",14933 => "01010000",14934 => "01000100",14935 => "11000100",14936 => "01111011",14937 => "11001010",14938 => "00001010",14939 => "00110111",14940 => "11111110",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00111010" report "FAIL high bits" severity failure;
assert RAM(0) = "01011100" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
