 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "10011000",3 => "01100100",4 => "11001110",5 => "00111110",6 => "01101010",7 => "00110110",8 => "10110111",9 => "01010000",10 => "10001100",11 => "11111101",12 => "11011000",13 => "01011011",14 => "11110110",15 => "11100010",16 => "01011011",17 => "11110000",18 => "10000001",19 => "10001100",20 => "00000010",21 => "11100010",22 => "10011010",23 => "10011101",24 => "01001101",25 => "01100101",26 => "00100101",27 => "00111010",28 => "10101010",29 => "10110101",30 => "10111001",31 => "11111110",32 => "10010111",33 => "10010000",34 => "00110111",35 => "00110100",36 => "11110111",37 => "01101000",38 => "01010000",39 => "00000100",40 => "10110110",41 => "00111001",42 => "00100111",43 => "11110001",44 => "00111100",45 => "11001101",46 => "11001010",47 => "11010110",48 => "01011101",49 => "00000101",50 => "00110110",51 => "00011011",52 => "11000111",53 => "11100011",54 => "01000101",55 => "11111000",56 => "01110100",57 => "10111100",58 => "00111001",59 => "01111111",60 => "01001011",61 => "00100010",62 => "10110111",63 => "00010100",64 => "11001100",65 => "10001111",66 => "11101110",67 => "00010000",68 => "11100000",69 => "10000111",70 => "10100100",71 => "00101111",72 => "00101011",73 => "11001111",74 => "10100110",75 => "10001000",76 => "00010100",77 => "11000000",78 => "01101001",79 => "00101111",80 => "11101010",81 => "00010001",82 => "11111001",83 => "01111111",84 => "11000000",85 => "11000000",86 => "10011101",87 => "01111110",88 => "11001110",89 => "10100101",90 => "01011101",91 => "00100000",92 => "11111110",93 => "01010001",94 => "11101010",95 => "01010101",96 => "00011100",97 => "01101111",98 => "01111000",99 => "10100011",100 => "00010010",101 => "10111111",102 => "01010010",103 => "01100000",104 => "01001110",105 => "00101110",106 => "01000101",107 => "10010100",108 => "00101101",109 => "01101001",110 => "11000101",111 => "10111110",112 => "10100011",113 => "11010111",114 => "11100100",115 => "11101100",116 => "00110000",117 => "10001101",118 => "01010011",119 => "01110110",120 => "01100010",121 => "10111001",122 => "01000001",123 => "11111111",124 => "10011110",125 => "10100011",126 => "11010000",127 => "10111011",128 => "11000000",129 => "10110011",130 => "01000011",131 => "00000010",132 => "11010011",133 => "01010100",134 => "00100111",135 => "00000000",136 => "10011111",137 => "11011111",138 => "00000111",139 => "00010111",140 => "11001001",141 => "11110010",142 => "11111001",143 => "10011110",144 => "10010101",145 => "10110100",146 => "00000011",147 => "01011011",148 => "10101010",149 => "10110010",150 => "10100010",151 => "01101101",152 => "11001100",153 => "11000101",154 => "10101111",155 => "11100010",156 => "00110011",157 => "11111011",158 => "10111001",159 => "00110101",160 => "10101010",161 => "11100010",162 => "01010101",163 => "00101010",164 => "11100101",165 => "11110100",166 => "00010111",167 => "00101001",168 => "00111011",169 => "00011001",170 => "11101010",171 => "11101101",172 => "01000000",173 => "10100011",174 => "10100101",175 => "10101110",176 => "10101011",177 => "00111110",178 => "10011101",179 => "00011000",180 => "11011111",181 => "00011000",182 => "01100110",183 => "01111111",184 => "00011010",185 => "00100001",186 => "10111001",187 => "10111001",188 => "00111000",189 => "01000000",190 => "01100000",191 => "11111111",192 => "01100100",193 => "00111111",194 => "01010110",195 => "11010101",196 => "10110110",197 => "11000110",198 => "10101010",199 => "00011111",200 => "11001010",201 => "00110110",202 => "01010101",203 => "11000010",204 => "00011101",205 => "01101011",206 => "10110100",207 => "11011001",208 => "11011001",209 => "01110001",210 => "10001001",211 => "01110100",212 => "11100111",213 => "10001100",214 => "00100110",215 => "01111101",216 => "10100011",217 => "11011101",218 => "01001110",219 => "01000111",220 => "01100110",221 => "00100110",222 => "11101000",223 => "11011100",224 => "10011011",225 => "11101111",226 => "10000001",227 => "00101011",228 => "10111101",229 => "10011110",230 => "11011011",231 => "01110010",232 => "00101101",233 => "11011001",234 => "11111111",235 => "00100010",236 => "11111101",237 => "11101001",238 => "01010100",239 => "11101101",240 => "01001111",241 => "10010001",242 => "11101100",243 => "00111100",244 => "00001100",245 => "11111001",246 => "01101111",247 => "10101001",248 => "01101110",249 => "01000110",250 => "10010100",251 => "00011011",252 => "00100111",253 => "01101111",254 => "00101010",255 => "00101100",256 => "01111000",257 => "01110111",258 => "11000110",259 => "00100000",260 => "00110101",261 => "11000011",262 => "10011101",263 => "01001001",264 => "01100110",265 => "00100011",266 => "11111100",267 => "01101000",268 => "10101100",269 => "01100101",270 => "11111111",271 => "00011101",272 => "11110110",273 => "01001100",274 => "01111010",275 => "10101110",276 => "11100001",277 => "11011101",278 => "00100100",279 => "01110101",280 => "00110000",281 => "01100101",282 => "10101001",283 => "10110111",284 => "00010011",285 => "01000010",286 => "11000010",287 => "11110100",288 => "11001000",289 => "11001111",290 => "11011010",291 => "00011010",292 => "01110000",293 => "00010110",294 => "00001000",295 => "01011011",296 => "00101000",297 => "01001011",298 => "00111011",299 => "01001010",300 => "01001101",301 => "00111111",302 => "01000100",303 => "11100111",304 => "01110001",305 => "00010001",306 => "11110111",307 => "01010000",308 => "10010111",309 => "10000010",310 => "10011101",311 => "01011000",312 => "10000110",313 => "11110111",314 => "11101101",315 => "10101001",316 => "01011100",317 => "00100100",318 => "10010000",319 => "01011111",320 => "10100100",321 => "00001000",322 => "11010000",323 => "00000110",324 => "11000101",325 => "01111010",326 => "11110011",327 => "01110001",328 => "01010110",329 => "10100100",330 => "00101001",331 => "00100000",332 => "10101000",333 => "11110001",334 => "01111000",335 => "10001001",336 => "11111110",337 => "00110011",338 => "00010101",339 => "01011001",340 => "01100101",341 => "01110111",342 => "11000111",343 => "10001110",344 => "11100101",345 => "00001110",346 => "00110001",347 => "11011110",348 => "10110000",349 => "00000110",350 => "10100100",351 => "01101100",352 => "00001011",353 => "01000101",354 => "11110011",355 => "01011110",356 => "00001110",357 => "00101000",358 => "01100111",359 => "01101011",360 => "11110010",361 => "10001001",362 => "01001100",363 => "10101101",364 => "11010111",365 => "11111011",366 => "10100100",367 => "11111010",368 => "01001100",369 => "11101100",370 => "11110011",371 => "00111111",372 => "11111000",373 => "00000010",374 => "10000010",375 => "10101001",376 => "00000100",377 => "11010001",378 => "00110101",379 => "00101111",380 => "11001101",381 => "00010011",382 => "10010101",383 => "11110001",384 => "01110001",385 => "01010011",386 => "01110111",387 => "10111001",388 => "11010011",389 => "10010010",390 => "11100110",391 => "11110111",392 => "01111011",393 => "01100111",394 => "00000011",395 => "11010001",396 => "10010110",397 => "10010001",398 => "00011110",399 => "01010010",400 => "11111111",401 => "01011100",402 => "10010000",403 => "11110101",404 => "11100010",405 => "00100011",406 => "11100011",407 => "11111100",408 => "01011111",409 => "00110110",410 => "00111000",411 => "01010011",412 => "11110011",413 => "01001100",414 => "11001001",415 => "11010000",416 => "01100000",417 => "11111010",418 => "10111101",419 => "00100010",420 => "10111011",421 => "11011011",422 => "11011101",423 => "00111110",424 => "00000110",425 => "10011001",426 => "00110101",427 => "00110000",428 => "00011000",429 => "01011110",430 => "10100111",431 => "11001100",432 => "10010110",433 => "11010101",434 => "11000010",435 => "00110110",436 => "00110111",437 => "10001111",438 => "10000111",439 => "11110101",440 => "00010101",441 => "10100000",442 => "11110111",443 => "10101100",444 => "01110101",445 => "01010011",446 => "00001110",447 => "00010110",448 => "11101101",449 => "00111001",450 => "01000100",451 => "00101101",452 => "11001101",453 => "01001110",454 => "00101101",455 => "00101100",456 => "11101010",457 => "11101010",458 => "01111001",459 => "01100101",460 => "11100111",461 => "11011101",462 => "01011000",463 => "01100110",464 => "00000011",465 => "11010100",466 => "10111010",467 => "00100100",468 => "01110011",469 => "00000101",470 => "10001100",471 => "10100001",472 => "01111000",473 => "11111110",474 => "11001100",475 => "01010101",476 => "10111111",477 => "10111001",478 => "10110000",479 => "00001110",480 => "11001000",481 => "00000010",482 => "10101110",483 => "10011100",484 => "00100110",485 => "10110110",486 => "01000000",487 => "00011101",488 => "00101010",489 => "01100010",490 => "00111101",491 => "01100010",492 => "10101001",493 => "10000100",494 => "10100001",495 => "10111100",496 => "00010100",497 => "10100111",498 => "00110100",499 => "11001111",500 => "11111110",501 => "10101111",502 => "10111100",503 => "01010001",504 => "10100111",505 => "01110011",506 => "01101110",507 => "11001011",508 => "01000101",509 => "01001100",510 => "11010100",511 => "01011010",512 => "10000110",513 => "01001000",514 => "01010000",515 => "00001010",516 => "00100101",517 => "10110011",518 => "00010101",519 => "11111101",520 => "10010000",521 => "00001000",522 => "11100111",523 => "01101001",524 => "10111010",525 => "01000001",526 => "00011110",527 => "11010111",528 => "11110010",529 => "10011111",530 => "01101110",531 => "10011010",532 => "10011011",533 => "10010011",534 => "01101010",535 => "11110101",536 => "11101100",537 => "11010100",538 => "10011101",539 => "10110110",540 => "01110100",541 => "10010011",542 => "01101110",543 => "00000101",544 => "10101000",545 => "11111101",546 => "10010001",547 => "10010011",548 => "00001011",549 => "10110101",550 => "10111000",551 => "11010100",552 => "10111110",553 => "11100001",554 => "10000010",555 => "01010110",556 => "10111010",557 => "11100000",558 => "11100001",559 => "10001100",560 => "11101111",561 => "00001101",562 => "10001110",563 => "10001101",564 => "00100011",565 => "01000101",566 => "01100001",567 => "01001100",568 => "00001110",569 => "01110011",570 => "00101100",571 => "01101101",572 => "11100000",573 => "01001101",574 => "00000010",575 => "01100110",576 => "01010000",577 => "00111101",578 => "11111001",579 => "11001111",580 => "10111111",581 => "11111000",582 => "11101011",583 => "11010100",584 => "11010111",585 => "10101110",586 => "10010001",587 => "00100011",588 => "01100110",589 => "01110111",590 => "01011101",591 => "01110001",592 => "01101010",593 => "00010110",594 => "00001001",595 => "10111010",596 => "00000001",597 => "10100101",598 => "01010101",599 => "10000100",600 => "10111100",601 => "01111111",602 => "00011001",603 => "10011000",604 => "00111100",605 => "10111110",606 => "11100000",607 => "11111101",608 => "00011000",609 => "10110101",610 => "00101111",611 => "10010000",612 => "00000000",613 => "00000111",614 => "00001000",615 => "00111010",616 => "00001010",617 => "10101000",618 => "11010001",619 => "00101111",620 => "11101101",621 => "00010000",622 => "11100101",623 => "11010010",624 => "10101000",625 => "01111101",626 => "01000001",627 => "10110100",628 => "11110101",629 => "01111110",630 => "01001111",631 => "00000001",632 => "10011111",633 => "10110110",634 => "01001101",635 => "01001111",636 => "00110001",637 => "01011001",638 => "01011101",639 => "11101101",640 => "10101010",641 => "01001000",642 => "10110010",643 => "00101111",644 => "00001000",645 => "01011010",646 => "11001010",647 => "01011011",648 => "10111110",649 => "10010111",650 => "01111111",651 => "11010110",652 => "00100011",653 => "11111000",654 => "10000100",655 => "01101110",656 => "11110101",657 => "01000011",658 => "11001101",659 => "11111111",660 => "10001111",661 => "00101111",662 => "00101010",663 => "01101100",664 => "11010101",665 => "11010011",666 => "10011000",667 => "11011111",668 => "01011110",669 => "11001001",670 => "01001010",671 => "11010111",672 => "11111000",673 => "01000010",674 => "00011101",675 => "01101000",676 => "00100100",677 => "11100010",678 => "01101100",679 => "10111101",680 => "01010111",681 => "00001100",682 => "10001101",683 => "10110010",684 => "10010111",685 => "01111011",686 => "00101111",687 => "11110001",688 => "00100011",689 => "01001010",690 => "01110011",691 => "01111110",692 => "10110001",693 => "00011100",694 => "10100100",695 => "00111011",696 => "10000100",697 => "00110000",698 => "01110111",699 => "10010101",700 => "01001001",701 => "11110010",702 => "11101001",703 => "01110011",704 => "00010010",705 => "10110100",706 => "11110110",707 => "00001100",708 => "10110110",709 => "01010010",710 => "00110101",711 => "00001110",712 => "10011111",713 => "00100111",714 => "01110001",715 => "11101111",716 => "01100110",717 => "11110110",718 => "01101101",719 => "10000101",720 => "00011110",721 => "00010011",722 => "01101010",723 => "11100110",724 => "00010111",725 => "10000010",726 => "10101100",727 => "01010110",728 => "10001011",729 => "01100111",730 => "00110000",731 => "00010000",732 => "00010101",733 => "01010100",734 => "00100011",735 => "10110100",736 => "11011011",737 => "10001010",738 => "11000001",739 => "11011111",740 => "01111000",741 => "00010101",742 => "01110001",743 => "11000101",744 => "00001111",745 => "00101111",746 => "00100100",747 => "00100110",748 => "00010001",749 => "00110110",750 => "10101011",751 => "11011111",752 => "10011010",753 => "10110111",754 => "00101100",755 => "10101111",756 => "00111101",757 => "10000100",758 => "11111000",759 => "11011110",760 => "10101000",761 => "00010011",762 => "10100011",763 => "00110010",764 => "01011101",765 => "01001011",766 => "10101111",767 => "10110111",768 => "01100110",769 => "10001011",770 => "00001110",771 => "10101001",772 => "10100000",773 => "00101001",774 => "00001000",775 => "00000100",776 => "10001011",777 => "00100101",778 => "00111010",779 => "11111101",780 => "11100011",781 => "00100110",782 => "10011100",783 => "01100111",784 => "00110101",785 => "00110000",786 => "11011001",787 => "00111110",788 => "10011101",789 => "11110100",790 => "10011101",791 => "00111100",792 => "10101011",793 => "10101110",794 => "10101100",795 => "11010001",796 => "00101101",797 => "11000111",798 => "01001010",799 => "01001001",800 => "01001010",801 => "11101101",802 => "00000110",803 => "11011110",804 => "11111101",805 => "01100110",806 => "11100001",807 => "00000010",808 => "10011100",809 => "11100011",810 => "00011111",811 => "01010111",812 => "10010010",813 => "11011010",814 => "00001011",815 => "10100111",816 => "11100001",817 => "11101011",818 => "11111001",819 => "11101000",820 => "11000011",821 => "10110110",822 => "00010111",823 => "01110000",824 => "11001010",825 => "11101101",826 => "11000000",827 => "00010000",828 => "10111100",829 => "00011001",830 => "11011000",831 => "10100110",832 => "01111000",833 => "00011101",834 => "00011100",835 => "10100110",836 => "10011111",837 => "01101101",838 => "11110100",839 => "01011010",840 => "00000100",841 => "01011000",842 => "11110101",843 => "01010101",844 => "10110100",845 => "00001110",846 => "11011010",847 => "00100010",848 => "11111000",849 => "00110010",850 => "11010101",851 => "10110111",852 => "10011101",853 => "01101001",854 => "00011110",855 => "00000001",856 => "11111000",857 => "01100000",858 => "10000011",859 => "10001010",860 => "01010001",861 => "00100111",862 => "11011101",863 => "10010011",864 => "01111001",865 => "11011101",866 => "10111101",867 => "11111001",868 => "00111111",869 => "01001110",870 => "11110111",871 => "11001101",872 => "01110010",873 => "10101000",874 => "01101101",875 => "01001100",876 => "11000101",877 => "10011110",878 => "00011101",879 => "01111101",880 => "10111111",881 => "10001010",882 => "10001100",883 => "01000010",884 => "11101100",885 => "00101111",886 => "01110000",887 => "11100111",888 => "00000010",889 => "00000001",890 => "10110111",891 => "00110111",892 => "00000010",893 => "01000011",894 => "11011000",895 => "00101100",896 => "10011011",897 => "00010011",898 => "11101100",899 => "01000101",900 => "11011100",901 => "10100011",902 => "00101110",903 => "11010110",904 => "11011010",905 => "00010101",906 => "11000011",907 => "11111010",908 => "10000100",909 => "11010101",910 => "11010001",911 => "01100000",912 => "10111001",913 => "10010111",914 => "10101110",915 => "00100100",916 => "11001011",917 => "01111110",918 => "00100100",919 => "10110110",920 => "10111001",921 => "11000000",922 => "10011010",923 => "01010011",924 => "10000101",925 => "00111110",926 => "11000001",927 => "10100110",928 => "10010110",929 => "10101101",930 => "11000110",931 => "01011111",932 => "10111001",933 => "01110001",934 => "00100010",935 => "01010101",936 => "10011000",937 => "10101110",938 => "00001001",939 => "01100000",940 => "11001110",941 => "10000101",942 => "10001000",943 => "11010000",944 => "10010001",945 => "11011000",946 => "00010010",947 => "00101101",948 => "00111111",949 => "10011011",950 => "01101001",951 => "10110100",952 => "01000010",953 => "10010111",954 => "11010000",955 => "01110111",956 => "01111010",957 => "01110010",958 => "00011110",959 => "10111111",960 => "11101010",961 => "11000011",962 => "00000011",963 => "11111000",964 => "10101010",965 => "10100111",966 => "10100110",967 => "01111110",968 => "01111011",969 => "11111100",970 => "10110110",971 => "11110000",972 => "01101111",973 => "00000000",974 => "11011000",975 => "00000010",976 => "01110011",977 => "10100100",978 => "01110110",979 => "01101011",980 => "10010100",981 => "01101001",982 => "11110011",983 => "11100010",984 => "00110101",985 => "11001101",986 => "11110010",987 => "11011011",988 => "01001100",989 => "00000101",990 => "00111010",991 => "01110110",992 => "01101011",993 => "00100111",994 => "00000100",995 => "00001001",996 => "00000001",997 => "00001110",998 => "00110011",999 => "00010010",1000 => "00011100",1001 => "01001010",1002 => "00111010",1003 => "00011011",1004 => "01010100",1005 => "11100101",1006 => "11101001",1007 => "10110011",1008 => "11001101",1009 => "11111001",1010 => "01001101",1011 => "01010111",1012 => "10111010",1013 => "00101000",1014 => "00011000",1015 => "11001100",1016 => "01100001",1017 => "10111111",1018 => "01111100",1019 => "01010100",1020 => "00010111",1021 => "00100111",1022 => "00101110",1023 => "10011100",1024 => "11100110",1025 => "11100100",1026 => "10001101",1027 => "01110110",1028 => "10011000",1029 => "11110010",1030 => "01001100",1031 => "10101101",1032 => "01101110",1033 => "11011000",1034 => "01011010",1035 => "11010011",1036 => "01010100",1037 => "01010110",1038 => "11110000",1039 => "01110110",1040 => "01001111",1041 => "11101011",1042 => "10111001",1043 => "10010000",1044 => "00000110",1045 => "00100111",1046 => "00100111",1047 => "00101000",1048 => "01110111",1049 => "01110010",1050 => "01100111",1051 => "01000010",1052 => "00010111",1053 => "01110100",1054 => "01000011",1055 => "10000101",1056 => "11010000",1057 => "00101011",1058 => "10101010",1059 => "00101100",1060 => "00000010",1061 => "10100110",1062 => "00101111",1063 => "01111000",1064 => "10010001",1065 => "00110100",1066 => "00010010",1067 => "10101110",1068 => "10001111",1069 => "01110100",1070 => "10011101",1071 => "01000111",1072 => "01000100",1073 => "10111101",1074 => "11001010",1075 => "01001100",1076 => "10011100",1077 => "01111010",1078 => "01111111",1079 => "10100100",1080 => "00100011",1081 => "00111110",1082 => "11001010",1083 => "00000110",1084 => "01110101",1085 => "01110001",1086 => "11001111",1087 => "11110100",1088 => "10011100",1089 => "00110101",1090 => "00010110",1091 => "01101110",1092 => "00111100",1093 => "10000101",1094 => "00010010",1095 => "00100010",1096 => "10000100",1097 => "01101000",1098 => "00110110",1099 => "00011001",1100 => "00110101",1101 => "01110001",1102 => "11011000",1103 => "11111110",1104 => "11000100",1105 => "01000011",1106 => "00011011",1107 => "10010011",1108 => "01010011",1109 => "01001000",1110 => "11000000",1111 => "11110100",1112 => "00111101",1113 => "10101110",1114 => "00001110",1115 => "10100001",1116 => "10110111",1117 => "10100000",1118 => "00101001",1119 => "11010010",1120 => "00011000",1121 => "00000001",1122 => "11111100",1123 => "10111100",1124 => "10111110",1125 => "00000011",1126 => "00110101",1127 => "00001010",1128 => "10011000",1129 => "01100111",1130 => "11000011",1131 => "00111101",1132 => "01100011",1133 => "00001111",1134 => "10111011",1135 => "10110011",1136 => "01000010",1137 => "00111010",1138 => "10110011",1139 => "11111111",1140 => "00110001",1141 => "11100010",1142 => "01000011",1143 => "11110110",1144 => "10001010",1145 => "11101111",1146 => "10010100",1147 => "00010110",1148 => "11000110",1149 => "10111110",1150 => "01000001",1151 => "01111001",1152 => "00001011",1153 => "10011101",1154 => "00101011",1155 => "11101011",1156 => "10110000",1157 => "01011111",1158 => "11011010",1159 => "01100001",1160 => "00110001",1161 => "01000111",1162 => "00010010",1163 => "10000000",1164 => "11101110",1165 => "10100010",1166 => "01101111",1167 => "00010110",1168 => "01001100",1169 => "00101110",1170 => "01111001",1171 => "01000101",1172 => "01000111",1173 => "11001110",1174 => "10010110",1175 => "11010000",1176 => "11101100",1177 => "00001110",1178 => "11111101",1179 => "01110000",1180 => "00101011",1181 => "10011000",1182 => "11110010",1183 => "01110010",1184 => "00111011",1185 => "01100111",1186 => "10010101",1187 => "10111111",1188 => "00110001",1189 => "11010010",1190 => "00010111",1191 => "10111000",1192 => "10110011",1193 => "11100000",1194 => "10111110",1195 => "11001001",1196 => "00010101",1197 => "00011000",1198 => "10010100",1199 => "01101011",1200 => "11101011",1201 => "10110010",1202 => "11111010",1203 => "11001011",1204 => "11110011",1205 => "10011010",1206 => "10000001",1207 => "10011111",1208 => "01000000",1209 => "11100011",1210 => "10000101",1211 => "00111010",1212 => "11010000",1213 => "10101001",1214 => "11011010",1215 => "00101100",1216 => "00010110",1217 => "00010001",1218 => "01001110",1219 => "00000110",1220 => "00110001",1221 => "00001011",1222 => "11010110",1223 => "00001101",1224 => "00011011",1225 => "01111110",1226 => "10100110",1227 => "00011111",1228 => "00011101",1229 => "11100100",1230 => "01010110",1231 => "00001001",1232 => "01110100",1233 => "11110010",1234 => "10011100",1235 => "10011000",1236 => "01100100",1237 => "00011001",1238 => "10001100",1239 => "01110001",1240 => "00010110",1241 => "11110001",1242 => "10100100",1243 => "11010010",1244 => "11000000",1245 => "01010101",1246 => "01010000",1247 => "01011000",1248 => "11110001",1249 => "10101011",1250 => "00000110",1251 => "00010011",1252 => "11100100",1253 => "10110001",1254 => "10010000",1255 => "11100101",1256 => "01100101",1257 => "11111001",1258 => "11100101",1259 => "00001100",1260 => "11010101",1261 => "11100011",1262 => "11001010",1263 => "01001111",1264 => "11111001",1265 => "11101110",1266 => "01100101",1267 => "11100111",1268 => "11000000",1269 => "11011010",1270 => "10101010",1271 => "11001000",1272 => "01111011",1273 => "11111111",1274 => "10111111",1275 => "00100101",1276 => "10100011",1277 => "00010100",1278 => "10101100",1279 => "10001111",1280 => "01100000",1281 => "10011100",1282 => "10011001",1283 => "10000011",1284 => "10010101",1285 => "01010101",1286 => "10011011",1287 => "11011000",1288 => "01110001",1289 => "11010111",1290 => "11100000",1291 => "11001100",1292 => "00010011",1293 => "00010110",1294 => "01100111",1295 => "01110101",1296 => "00101111",1297 => "10111111",1298 => "00010111",1299 => "01100110",1300 => "00011011",1301 => "01101110",1302 => "11101001",1303 => "00110001",1304 => "01100110",1305 => "01011011",1306 => "00000111",1307 => "01000110",1308 => "10110011",1309 => "00100011",1310 => "11101001",1311 => "01011100",1312 => "01111111",1313 => "10010011",1314 => "11001011",1315 => "10000100",1316 => "10000111",1317 => "01001010",1318 => "11011000",1319 => "11110001",1320 => "11110000",1321 => "01101100",1322 => "01101100",1323 => "00010000",1324 => "11011110",1325 => "10100111",1326 => "01000101",1327 => "10011110",1328 => "00010010",1329 => "10110000",1330 => "00000001",1331 => "11110111",1332 => "01111001",1333 => "11011101",1334 => "10100110",1335 => "00110001",1336 => "11011011",1337 => "10100010",1338 => "10001101",1339 => "10101000",1340 => "01010101",1341 => "10111100",1342 => "00000001",1343 => "10101011",1344 => "00110100",1345 => "01100010",1346 => "01010101",1347 => "11110011",1348 => "11111101",1349 => "10011001",1350 => "11011111",1351 => "10101110",1352 => "01110100",1353 => "11100110",1354 => "10100010",1355 => "00110101",1356 => "11100001",1357 => "01000100",1358 => "01000100",1359 => "10101100",1360 => "01110100",1361 => "01111010",1362 => "11101011",1363 => "00010010",1364 => "10110101",1365 => "01111101",1366 => "11101010",1367 => "11100011",1368 => "01010100",1369 => "11000011",1370 => "10001010",1371 => "00000100",1372 => "11111101",1373 => "01101011",1374 => "01001001",1375 => "00100011",1376 => "11110100",1377 => "00010100",1378 => "11011110",1379 => "00000011",1380 => "01100000",1381 => "11110001",1382 => "01000111",1383 => "11010010",1384 => "10000001",1385 => "10110010",1386 => "11111101",1387 => "11000100",1388 => "10100011",1389 => "10111010",1390 => "11000111",1391 => "10100101",1392 => "01101110",1393 => "00110100",1394 => "10100101",1395 => "01001001",1396 => "00101110",1397 => "00011000",1398 => "00110000",1399 => "11001110",1400 => "01000001",1401 => "11110011",1402 => "00101010",1403 => "11100110",1404 => "00000000",1405 => "11111011",1406 => "10000100",1407 => "00011110",1408 => "00110000",1409 => "01101111",1410 => "00010110",1411 => "00001010",1412 => "10011000",1413 => "11010110",1414 => "10010000",1415 => "10110101",1416 => "10100011",1417 => "01000010",1418 => "11101110",1419 => "10111101",1420 => "01110010",1421 => "11000100",1422 => "01011101",1423 => "00010101",1424 => "01101011",1425 => "11110101",1426 => "01000011",1427 => "11011101",1428 => "01010001",1429 => "10001010",1430 => "10001001",1431 => "01000001",1432 => "11000010",1433 => "11010101",1434 => "01010100",1435 => "01010011",1436 => "10111100",1437 => "00010010",1438 => "10110000",1439 => "00000000",1440 => "01011000",1441 => "01010001",1442 => "00110101",1443 => "11011101",1444 => "00101001",1445 => "00000101",1446 => "01001000",1447 => "10011011",1448 => "10001111",1449 => "00010100",1450 => "10010110",1451 => "00011000",1452 => "01010100",1453 => "01000101",1454 => "11100010",1455 => "10111110",1456 => "01001100",1457 => "11101101",1458 => "00001010",1459 => "01110000",1460 => "01011100",1461 => "01001111",1462 => "10101010",1463 => "10000000",1464 => "00100001",1465 => "00010010",1466 => "10010111",1467 => "10000010",1468 => "00110101",1469 => "10100101",1470 => "01100110",1471 => "11110101",1472 => "01010011",1473 => "01100011",1474 => "11110010",1475 => "11001001",1476 => "01011000",1477 => "01111001",1478 => "00101110",1479 => "10011100",1480 => "11101000",1481 => "11101100",1482 => "01110001",1483 => "10011000",1484 => "01001100",1485 => "11100011",1486 => "00110011",1487 => "10101000",1488 => "01100001",1489 => "11111011",1490 => "11000011",1491 => "10101010",1492 => "01111011",1493 => "10101000",1494 => "11010010",1495 => "00001101",1496 => "00101110",1497 => "01100001",1498 => "01100110",1499 => "10000011",1500 => "01011101",1501 => "11111110",1502 => "11001110",1503 => "10101000",1504 => "10110000",1505 => "00001001",1506 => "01000001",1507 => "01110010",1508 => "01100010",1509 => "01101111",1510 => "01000101",1511 => "01100001",1512 => "11101100",1513 => "11000011",1514 => "11010010",1515 => "01101110",1516 => "01000000",1517 => "00000011",1518 => "10101101",1519 => "11010111",1520 => "10000100",1521 => "11100011",1522 => "01000001",1523 => "10111010",1524 => "10001011",1525 => "11101001",1526 => "00101111",1527 => "11011101",1528 => "11100101",1529 => "11000110",1530 => "10101000",1531 => "01110010",1532 => "00100011",1533 => "10010010",1534 => "01100000",1535 => "11110011",1536 => "01010011",1537 => "01010110",1538 => "01111111",1539 => "10110110",1540 => "10000001",1541 => "01010100",1542 => "00101100",1543 => "11010000",1544 => "00110001",1545 => "11000110",1546 => "00101001",1547 => "10000100",1548 => "11000011",1549 => "01010110",1550 => "01100110",1551 => "01000001",1552 => "10111111",1553 => "10010101",1554 => "10100000",1555 => "10111001",1556 => "11110101",1557 => "00001111",1558 => "11000111",1559 => "01111111",1560 => "10111010",1561 => "10011010",1562 => "01010101",1563 => "11010010",1564 => "10100111",1565 => "10101111",1566 => "00000111",1567 => "01001010",1568 => "01001001",1569 => "00110000",1570 => "10000001",1571 => "11101100",1572 => "10010110",1573 => "11111100",1574 => "10110011",1575 => "10110001",1576 => "01001100",1577 => "10111011",1578 => "00101111",1579 => "11011011",1580 => "11100100",1581 => "10101001",1582 => "10010110",1583 => "00101101",1584 => "00011011",1585 => "10100001",1586 => "00101010",1587 => "11001111",1588 => "01111111",1589 => "01010000",1590 => "00110000",1591 => "01011000",1592 => "00011101",1593 => "10100100",1594 => "01001101",1595 => "00110011",1596 => "01010100",1597 => "01100001",1598 => "01110111",1599 => "11111101",1600 => "11100000",1601 => "11000010",1602 => "11000001",1603 => "11001011",1604 => "11100111",1605 => "10011010",1606 => "10000010",1607 => "00010111",1608 => "00010111",1609 => "11111001",1610 => "10101011",1611 => "01000000",1612 => "01111001",1613 => "00001101",1614 => "11110110",1615 => "01000101",1616 => "11110110",1617 => "11011111",1618 => "01111110",1619 => "00101101",1620 => "01010011",1621 => "00100001",1622 => "00111101",1623 => "10011000",1624 => "00000110",1625 => "11001000",1626 => "00001110",1627 => "11111000",1628 => "01000011",1629 => "00001010",1630 => "01110110",1631 => "01000000",1632 => "00011011",1633 => "10011011",1634 => "00101000",1635 => "00100000",1636 => "01001100",1637 => "01000100",1638 => "11001101",1639 => "00001110",1640 => "01101001",1641 => "10111110",1642 => "01101001",1643 => "01111010",1644 => "10000101",1645 => "11010111",1646 => "10000111",1647 => "00000010",1648 => "10001101",1649 => "11100011",1650 => "00110111",1651 => "11100101",1652 => "01001100",1653 => "01110001",1654 => "10111001",1655 => "00010110",1656 => "00010111",1657 => "10100001",1658 => "01101111",1659 => "11100000",1660 => "01000111",1661 => "01101101",1662 => "10101111",1663 => "10001010",1664 => "01001100",1665 => "11100111",1666 => "10011001",1667 => "10001111",1668 => "00111110",1669 => "01100111",1670 => "00000101",1671 => "10010001",1672 => "11001101",1673 => "01101001",1674 => "01100001",1675 => "00000111",1676 => "01000110",1677 => "10110111",1678 => "00110100",1679 => "01011111",1680 => "10100100",1681 => "10001001",1682 => "10010110",1683 => "01111011",1684 => "00100101",1685 => "11100010",1686 => "10100001",1687 => "00111101",1688 => "11100110",1689 => "11011001",1690 => "11011001",1691 => "01010100",1692 => "11010001",1693 => "11100000",1694 => "10101110",1695 => "11101010",1696 => "11001011",1697 => "01101111",1698 => "11000001",1699 => "01101111",1700 => "00100011",1701 => "01001001",1702 => "00010101",1703 => "11110100",1704 => "10000100",1705 => "11000100",1706 => "00111010",1707 => "10010110",1708 => "01100100",1709 => "01001110",1710 => "11111111",1711 => "01110011",1712 => "10011111",1713 => "11001010",1714 => "10110110",1715 => "10000011",1716 => "10001100",1717 => "01110110",1718 => "11001000",1719 => "11010011",1720 => "10011111",1721 => "01100101",1722 => "10101010",1723 => "11000111",1724 => "10101000",1725 => "10000011",1726 => "01100100",1727 => "10110010",1728 => "00110110",1729 => "11100000",1730 => "01100111",1731 => "01011001",1732 => "10001001",1733 => "01100110",1734 => "11011111",1735 => "10100101",1736 => "00000000",1737 => "11100111",1738 => "00111111",1739 => "10101100",1740 => "10000000",1741 => "00001100",1742 => "01000111",1743 => "01011011",1744 => "11111110",1745 => "01000011",1746 => "00111110",1747 => "01010111",1748 => "01101010",1749 => "01101010",1750 => "11000000",1751 => "01011110",1752 => "00100010",1753 => "10001101",1754 => "10100100",1755 => "00001000",1756 => "01111101",1757 => "10111011",1758 => "11000110",1759 => "11001010",1760 => "11111001",1761 => "01001001",1762 => "00110011",1763 => "10000110",1764 => "01100000",1765 => "11110100",1766 => "00010001",1767 => "10101101",1768 => "01110001",1769 => "01010111",1770 => "11001000",1771 => "01101001",1772 => "10011110",1773 => "10011110",1774 => "01011001",1775 => "01100010",1776 => "00000111",1777 => "11000001",1778 => "10010011",1779 => "00111001",1780 => "11000110",1781 => "11101111",1782 => "01101110",1783 => "01010111",1784 => "11000011",1785 => "11011010",1786 => "10101101",1787 => "10110001",1788 => "10101001",1789 => "11011110",1790 => "01111110",1791 => "01110110",1792 => "10101001",1793 => "11000000",1794 => "01110010",1795 => "11101001",1796 => "01100101",1797 => "10011001",1798 => "01011001",1799 => "10100010",1800 => "00010011",1801 => "10110000",1802 => "00010110",1803 => "01001111",1804 => "10110100",1805 => "10110011",1806 => "01000010",1807 => "10011001",1808 => "01000101",1809 => "00010101",1810 => "11010011",1811 => "00100011",1812 => "10100101",1813 => "10110101",1814 => "00001100",1815 => "00110100",1816 => "01111111",1817 => "00110010",1818 => "11001000",1819 => "00001001",1820 => "00111000",1821 => "00111001",1822 => "01011111",1823 => "01000110",1824 => "10011110",1825 => "01111011",1826 => "01110000",1827 => "01111000",1828 => "11000001",1829 => "10110011",1830 => "10100111",1831 => "11111101",1832 => "01011101",1833 => "01111111",1834 => "10001011",1835 => "10011110",1836 => "11111101",1837 => "00010111",1838 => "11011101",1839 => "00100001",1840 => "01100010",1841 => "11001111",1842 => "01110111",1843 => "10001110",1844 => "01101110",1845 => "10110110",1846 => "01011100",1847 => "10100100",1848 => "10011000",1849 => "10000010",1850 => "11010001",1851 => "11001100",1852 => "01011000",1853 => "01111011",1854 => "00001100",1855 => "00100111",1856 => "00110011",1857 => "00100100",1858 => "11111001",1859 => "10000000",1860 => "10101001",1861 => "11001111",1862 => "01001000",1863 => "01011111",1864 => "11000101",1865 => "11010011",1866 => "01100110",1867 => "00011000",1868 => "01111010",1869 => "01011101",1870 => "10010101",1871 => "00000100",1872 => "11000100",1873 => "10010001",1874 => "01100100",1875 => "11001000",1876 => "11110111",1877 => "01100110",1878 => "01111011",1879 => "11100101",1880 => "10000000",1881 => "01110111",1882 => "00010001",1883 => "01011000",1884 => "01000100",1885 => "10000001",1886 => "10111011",1887 => "11111110",1888 => "01011111",1889 => "11101001",1890 => "01011010",1891 => "11111101",1892 => "11101010",1893 => "01010000",1894 => "11011101",1895 => "00000110",1896 => "10001011",1897 => "11000001",1898 => "10101000",1899 => "10000100",1900 => "10101111",1901 => "01001010",1902 => "01110010",1903 => "01111001",1904 => "11110110",1905 => "10100101",1906 => "01101110",1907 => "00001001",1908 => "11011011",1909 => "11010011",1910 => "11111010",1911 => "00101001",1912 => "01110010",1913 => "10000101",1914 => "11101001",1915 => "01001110",1916 => "01101000",1917 => "01111010",1918 => "01101000",1919 => "10110001",1920 => "10011010",1921 => "10101000",1922 => "00000101",1923 => "10100100",1924 => "10010010",1925 => "11101010",1926 => "10010000",1927 => "11110100",1928 => "01010001",1929 => "00101111",1930 => "10100001",1931 => "10100101",1932 => "00011110",1933 => "00110000",1934 => "11101111",1935 => "01000111",1936 => "00101101",1937 => "11010010",1938 => "00001101",1939 => "11110111",1940 => "00011100",1941 => "10010001",1942 => "00001110",1943 => "00000101",1944 => "01000010",1945 => "00000101",1946 => "11001001",1947 => "01010110",1948 => "01010000",1949 => "01001011",1950 => "00001001",1951 => "01001100",1952 => "10001101",1953 => "11111101",1954 => "01100011",1955 => "10011101",1956 => "00001100",1957 => "10111101",1958 => "01100111",1959 => "10100111",1960 => "11110100",1961 => "10001010",1962 => "00100110",1963 => "01011010",1964 => "01111111",1965 => "10011011",1966 => "01010010",1967 => "01111110",1968 => "00001111",1969 => "11110100",1970 => "11111110",1971 => "00101000",1972 => "11011000",1973 => "00101101",1974 => "11011001",1975 => "10100011",1976 => "11101101",1977 => "00100011",1978 => "11010011",1979 => "01100111",1980 => "00111011",1981 => "11010000",1982 => "01011100",1983 => "11000001",1984 => "00011100",1985 => "10001000",1986 => "11100111",1987 => "01001110",1988 => "11000010",1989 => "01001111",1990 => "00011011",1991 => "01001111",1992 => "01110110",1993 => "10100110",1994 => "10010101",1995 => "00010101",1996 => "01011001",1997 => "11111100",1998 => "01000110",1999 => "11110110",2000 => "00100000",2001 => "01000110",2002 => "10100010",2003 => "01101111",2004 => "11010000",2005 => "00000011",2006 => "10010001",2007 => "10001001",2008 => "01001001",2009 => "00010011",2010 => "11010011",2011 => "00111111",2012 => "01001011",2013 => "00000110",2014 => "01001011",2015 => "10100100",2016 => "01100111",2017 => "11000111",2018 => "11100101",2019 => "10001101",2020 => "00100100",2021 => "10011100",2022 => "10101010",2023 => "00111110",2024 => "01111110",2025 => "11010100",2026 => "00000111",2027 => "01000000",2028 => "01111000",2029 => "11010001",2030 => "10110010",2031 => "00010110",2032 => "00011101",2033 => "01011010",2034 => "11001111",2035 => "01000010",2036 => "11010100",2037 => "01100101",2038 => "00110100",2039 => "01001111",2040 => "01110010",2041 => "01101001",2042 => "11011110",2043 => "11111000",2044 => "11011101",2045 => "10010000",2046 => "01111001",2047 => "10011000",2048 => "11001000",2049 => "01101000",2050 => "01111111",2051 => "01000101",2052 => "01100101",2053 => "10001010",2054 => "00011001",2055 => "10001110",2056 => "01100010",2057 => "01110110",2058 => "11001010",2059 => "11001111",2060 => "01101011",2061 => "11010101",2062 => "01001100",2063 => "11011100",2064 => "01011010",2065 => "10000110",2066 => "10101000",2067 => "10100100",2068 => "10001010",2069 => "11010000",2070 => "11110101",2071 => "10100001",2072 => "00101011",2073 => "10011101",2074 => "01001100",2075 => "00111010",2076 => "11110010",2077 => "01100011",2078 => "01101010",2079 => "01110101",2080 => "00011000",2081 => "11110111",2082 => "11011111",2083 => "01111000",2084 => "01011100",2085 => "10011011",2086 => "01011001",2087 => "10001001",2088 => "11001000",2089 => "01011101",2090 => "00001110",2091 => "00001010",2092 => "01010100",2093 => "00011100",2094 => "11100110",2095 => "01010110",2096 => "00110101",2097 => "00011001",2098 => "10010000",2099 => "01001010",2100 => "01100100",2101 => "11111010",2102 => "11101001",2103 => "10101011",2104 => "00100011",2105 => "11110111",2106 => "11101100",2107 => "00011000",2108 => "00011100",2109 => "00100001",2110 => "10101110",2111 => "10001011",2112 => "00110111",2113 => "00110101",2114 => "01010001",2115 => "11011101",2116 => "10001000",2117 => "10101100",2118 => "11001111",2119 => "11011000",2120 => "00100011",2121 => "11101000",2122 => "10110110",2123 => "11101111",2124 => "11011110",2125 => "10000100",2126 => "00100010",2127 => "00001011",2128 => "01001000",2129 => "01111101",2130 => "01100110",2131 => "10001101",2132 => "01001000",2133 => "00001000",2134 => "00110000",2135 => "01101000",2136 => "00101010",2137 => "01011100",2138 => "10111000",2139 => "11011100",2140 => "01100011",2141 => "11111010",2142 => "11111100",2143 => "01110110",2144 => "00010100",2145 => "00111111",2146 => "11110111",2147 => "00110100",2148 => "01100011",2149 => "11111101",2150 => "10010000",2151 => "00001101",2152 => "01110001",2153 => "01000000",2154 => "00000100",2155 => "11001001",2156 => "00101110",2157 => "10111110",2158 => "01101110",2159 => "00100011",2160 => "00100001",2161 => "01001001",2162 => "01101100",2163 => "01101011",2164 => "01000001",2165 => "10101000",2166 => "00110010",2167 => "10100101",2168 => "00101100",2169 => "00101100",2170 => "00101010",2171 => "00010100",2172 => "10011000",2173 => "11101010",2174 => "01000100",2175 => "10001101",2176 => "10111011",2177 => "01001010",2178 => "01001101",2179 => "11001100",2180 => "10010010",2181 => "11001100",2182 => "00010011",2183 => "10101111",2184 => "11010010",2185 => "01111110",2186 => "11001101",2187 => "00011000",2188 => "11000100",2189 => "00010000",2190 => "00001100",2191 => "11011010",2192 => "10101000",2193 => "10000000",2194 => "01111011",2195 => "11010110",2196 => "00010100",2197 => "01111111",2198 => "01011000",2199 => "10000000",2200 => "11000010",2201 => "10001100",2202 => "01100001",2203 => "10001100",2204 => "01001111",2205 => "11110010",2206 => "11111010",2207 => "01010100",2208 => "10100011",2209 => "10111110",2210 => "11011110",2211 => "11111111",2212 => "11110001",2213 => "11100111",2214 => "01001011",2215 => "01000001",2216 => "00100110",2217 => "11100010",2218 => "10100010",2219 => "10000001",2220 => "11010111",2221 => "00110000",2222 => "10001101",2223 => "11010011",2224 => "10010000",2225 => "11011011",2226 => "01111110",2227 => "11001010",2228 => "11010101",2229 => "10110011",2230 => "10010011",2231 => "10111101",2232 => "11110011",2233 => "10000100",2234 => "11100100",2235 => "10101010",2236 => "01100100",2237 => "11101100",2238 => "11110011",2239 => "10000000",2240 => "01010001",2241 => "11100111",2242 => "11011001",2243 => "11001000",2244 => "11100100",2245 => "00001111",2246 => "01101100",2247 => "11110110",2248 => "00101111",2249 => "01001110",2250 => "10101111",2251 => "00000000",2252 => "01011111",2253 => "01101001",2254 => "11101011",2255 => "00111110",2256 => "11101011",2257 => "11010110",2258 => "11100101",2259 => "01001101",2260 => "11101101",2261 => "11101000",2262 => "10100011",2263 => "11111001",2264 => "00011000",2265 => "01111100",2266 => "01000100",2267 => "01111001",2268 => "10101001",2269 => "01100110",2270 => "01010101",2271 => "01101000",2272 => "11110010",2273 => "10000000",2274 => "00110011",2275 => "00000001",2276 => "00000010",2277 => "11100110",2278 => "01011101",2279 => "11111111",2280 => "01011011",2281 => "11100111",2282 => "01110111",2283 => "00101011",2284 => "11111100",2285 => "01001000",2286 => "01011010",2287 => "11111101",2288 => "11001100",2289 => "10000111",2290 => "11011010",2291 => "11011111",2292 => "00011111",2293 => "00100000",2294 => "01010000",2295 => "00101000",2296 => "10010000",2297 => "01111001",2298 => "10011001",2299 => "00101000",2300 => "11110000",2301 => "10001110",2302 => "11100011",2303 => "01011101",2304 => "01000100",2305 => "11001011",2306 => "11111001",2307 => "10100010",2308 => "00000000",2309 => "11111101",2310 => "01011001",2311 => "10011000",2312 => "11011011",2313 => "00101011",2314 => "01110100",2315 => "00010110",2316 => "11101000",2317 => "01011110",2318 => "01001001",2319 => "11110111",2320 => "00110000",2321 => "00000000",2322 => "01000000",2323 => "00101011",2324 => "10110011",2325 => "10001100",2326 => "10101110",2327 => "00000110",2328 => "00001111",2329 => "11100000",2330 => "10110011",2331 => "11010011",2332 => "11111010",2333 => "01111010",2334 => "10101111",2335 => "00011011",2336 => "10110000",2337 => "11100000",2338 => "10010110",2339 => "01000111",2340 => "11010101",2341 => "01011011",2342 => "01101111",2343 => "10010101",2344 => "00001111",2345 => "01110011",2346 => "10001110",2347 => "10001000",2348 => "01001001",2349 => "01111111",2350 => "01110110",2351 => "10011010",2352 => "11001010",2353 => "00110111",2354 => "10001110",2355 => "01011101",2356 => "00000111",2357 => "11101010",2358 => "01101111",2359 => "01011111",2360 => "11011101",2361 => "10101001",2362 => "00111110",2363 => "10010001",2364 => "01101111",2365 => "11011010",2366 => "01100001",2367 => "01100010",2368 => "01010000",2369 => "11110001",2370 => "00111001",2371 => "11100001",2372 => "10000011",2373 => "10010100",2374 => "11111001",2375 => "00000110",2376 => "11111111",2377 => "01111100",2378 => "10101100",2379 => "10101011",2380 => "10111110",2381 => "11010011",2382 => "11000100",2383 => "10000110",2384 => "00000010",2385 => "00110000",2386 => "10111100",2387 => "11101010",2388 => "01001101",2389 => "11100101",2390 => "10100101",2391 => "00110111",2392 => "00001001",2393 => "01000011",2394 => "11111001",2395 => "11010011",2396 => "01000011",2397 => "01101010",2398 => "11100101",2399 => "11101010",2400 => "01101100",2401 => "11100011",2402 => "11101000",2403 => "00101010",2404 => "01101010",2405 => "01011101",2406 => "01101101",2407 => "00000000",2408 => "00000101",2409 => "11101000",2410 => "01001110",2411 => "01111101",2412 => "11101111",2413 => "11001001",2414 => "00000110",2415 => "01011110",2416 => "11101011",2417 => "11100001",2418 => "01000010",2419 => "11100010",2420 => "00000101",2421 => "10010001",2422 => "01101010",2423 => "10101011",2424 => "00011001",2425 => "01001110",2426 => "01111010",2427 => "00110010",2428 => "00110100",2429 => "00001111",2430 => "11000110",2431 => "10110011",2432 => "01000010",2433 => "11001110",2434 => "01001011",2435 => "01111100",2436 => "00011000",2437 => "01100100",2438 => "11010101",2439 => "00101110",2440 => "00011110",2441 => "01001101",2442 => "01110011",2443 => "00111110",2444 => "10011000",2445 => "10111010",2446 => "11001110",2447 => "11011100",2448 => "00100111",2449 => "00110101",2450 => "11111011",2451 => "00111110",2452 => "11011000",2453 => "11001010",2454 => "11101110",2455 => "01111101",2456 => "00101001",2457 => "10000010",2458 => "00001010",2459 => "10010100",2460 => "00000101",2461 => "10100100",2462 => "00101010",2463 => "00111110",2464 => "01011010",2465 => "01010000",2466 => "01000010",2467 => "11100011",2468 => "00011011",2469 => "01110100",2470 => "11110101",2471 => "10111000",2472 => "11110101",2473 => "01010000",2474 => "11100111",2475 => "11100011",2476 => "00001100",2477 => "11011011",2478 => "00001110",2479 => "10001010",2480 => "11101100",2481 => "11100001",2482 => "01010100",2483 => "10100101",2484 => "10010100",2485 => "11010111",2486 => "11110000",2487 => "01010100",2488 => "01110100",2489 => "10111100",2490 => "11101011",2491 => "10000110",2492 => "01101011",2493 => "00100000",2494 => "00111110",2495 => "01011011",2496 => "01101100",2497 => "10111110",2498 => "01000111",2499 => "00001001",2500 => "10110110",2501 => "10111111",2502 => "10110010",2503 => "11101101",2504 => "01000011",2505 => "11111011",2506 => "01001101",2507 => "01001101",2508 => "11001101",2509 => "10000111",2510 => "00110010",2511 => "01111000",2512 => "10111110",2513 => "11100001",2514 => "00110101",2515 => "00111100",2516 => "00000010",2517 => "10100001",2518 => "00001000",2519 => "11010011",2520 => "01111111",2521 => "10000110",2522 => "11110011",2523 => "10000100",2524 => "11111010",2525 => "11011111",2526 => "01110101",2527 => "00011101",2528 => "11000101",2529 => "00101110",2530 => "00111000",2531 => "10100010",2532 => "01011000",2533 => "00101110",2534 => "00000111",2535 => "01111111",2536 => "01111111",2537 => "00110110",2538 => "11111001",2539 => "10001111",2540 => "01011001",2541 => "11000100",2542 => "10110011",2543 => "10110100",2544 => "00010111",2545 => "01110011",2546 => "01101001",2547 => "10100110",2548 => "01100010",2549 => "10010011",2550 => "01001110",2551 => "01100101",2552 => "11110010",2553 => "01110110",2554 => "11101111",2555 => "10111011",2556 => "10001010",2557 => "01011001",2558 => "00001011",2559 => "01101000",2560 => "10001111",2561 => "00000111",2562 => "10001111",2563 => "00101101",2564 => "00001011",2565 => "00011011",2566 => "11101100",2567 => "10000001",2568 => "10111111",2569 => "00010000",2570 => "00110101",2571 => "00000011",2572 => "00000110",2573 => "10110001",2574 => "11001110",2575 => "11110100",2576 => "00111000",2577 => "01111101",2578 => "01101100",2579 => "10011001",2580 => "00101100",2581 => "10100100",2582 => "01111000",2583 => "01110000",2584 => "00101110",2585 => "11110100",2586 => "01111001",2587 => "00111000",2588 => "01111010",2589 => "01000000",2590 => "01101101",2591 => "10001001",2592 => "11001000",2593 => "00011001",2594 => "00110011",2595 => "01101111",2596 => "10010010",2597 => "00010111",2598 => "01110100",2599 => "00111011",2600 => "11100111",2601 => "01111101",2602 => "10001101",2603 => "11111101",2604 => "11000111",2605 => "10100001",2606 => "00111101",2607 => "00111111",2608 => "10010101",2609 => "10011100",2610 => "11010110",2611 => "00011010",2612 => "00000000",2613 => "11100100",2614 => "00101111",2615 => "00010101",2616 => "01101011",2617 => "10101011",2618 => "01001101",2619 => "01011000",2620 => "10011001",2621 => "10111011",2622 => "01000100",2623 => "11101101",2624 => "01100010",2625 => "00100001",2626 => "10000011",2627 => "00100010",2628 => "00011110",2629 => "01001000",2630 => "01110011",2631 => "10000101",2632 => "10110111",2633 => "01110000",2634 => "11110011",2635 => "11100100",2636 => "00000110",2637 => "11111010",2638 => "01000010",2639 => "11100010",2640 => "11001010",2641 => "11100111",2642 => "10010001",2643 => "00101110",2644 => "01011000",2645 => "01100101",2646 => "11011110",2647 => "11111010",2648 => "11101101",2649 => "00011111",2650 => "10010100",2651 => "01000011",2652 => "10001111",2653 => "10011010",2654 => "10101011",2655 => "10010111",2656 => "11110000",2657 => "10001110",2658 => "11110100",2659 => "01101011",2660 => "00101011",2661 => "11011000",2662 => "01111000",2663 => "11001010",2664 => "11111000",2665 => "00011101",2666 => "11010100",2667 => "10000000",2668 => "10001011",2669 => "00101001",2670 => "01100101",2671 => "11100101",2672 => "10001101",2673 => "00011100",2674 => "01000101",2675 => "10010110",2676 => "01100011",2677 => "01101011",2678 => "10001011",2679 => "00001101",2680 => "10111010",2681 => "00010001",2682 => "00000011",2683 => "00111001",2684 => "00101011",2685 => "10001010",2686 => "11000111",2687 => "10101111",2688 => "01010110",2689 => "11001010",2690 => "00100001",2691 => "11101100",2692 => "00101111",2693 => "01110011",2694 => "10100100",2695 => "01011010",2696 => "10011010",2697 => "00000111",2698 => "10111101",2699 => "10001100",2700 => "11100010",2701 => "11101111",2702 => "01001001",2703 => "01011000",2704 => "00000011",2705 => "10101000",2706 => "01010000",2707 => "10001100",2708 => "00111001",2709 => "10010110",2710 => "01001110",2711 => "11111000",2712 => "10111010",2713 => "10011001",2714 => "11000110",2715 => "11100100",2716 => "00101011",2717 => "01101001",2718 => "00010100",2719 => "01001110",2720 => "00001100",2721 => "10011111",2722 => "11000100",2723 => "11010101",2724 => "01110001",2725 => "01101101",2726 => "01010110",2727 => "00011101",2728 => "01011010",2729 => "10000010",2730 => "00010110",2731 => "00011010",2732 => "00001011",2733 => "11110110",2734 => "01101010",2735 => "00101001",2736 => "01010000",2737 => "11010001",2738 => "01000000",2739 => "10100010",2740 => "00011001",2741 => "01001100",2742 => "01011111",2743 => "10110100",2744 => "01111000",2745 => "00101101",2746 => "01011010",2747 => "00001101",2748 => "10111110",2749 => "01000011",2750 => "01100010",2751 => "11001001",2752 => "10000000",2753 => "10100100",2754 => "10111100",2755 => "11000110",2756 => "11111101",2757 => "10110001",2758 => "01010100",2759 => "10111001",2760 => "11100111",2761 => "01000001",2762 => "01010010",2763 => "00101011",2764 => "11110110",2765 => "10111001",2766 => "01011010",2767 => "01110101",2768 => "10100101",2769 => "01110101",2770 => "10110110",2771 => "00101111",2772 => "01101010",2773 => "01110101",2774 => "01000111",2775 => "01111111",2776 => "01000000",2777 => "01001001",2778 => "01000001",2779 => "01110101",2780 => "10111001",2781 => "11111110",2782 => "00101110",2783 => "11100101",2784 => "11111000",2785 => "01010101",2786 => "01111010",2787 => "00011010",2788 => "10010111",2789 => "10011001",2790 => "11111010",2791 => "11110110",2792 => "11101000",2793 => "01101010",2794 => "00111010",2795 => "01011000",2796 => "01011111",2797 => "01111101",2798 => "00010010",2799 => "10110101",2800 => "00011011",2801 => "10111100",2802 => "10001000",2803 => "10001010",2804 => "11110100",2805 => "00111100",2806 => "10001010",2807 => "00111100",2808 => "00000000",2809 => "10010011",2810 => "11001101",2811 => "00100111",2812 => "00110001",2813 => "10100101",2814 => "00001000",2815 => "10100100",2816 => "00100111",2817 => "10101010",2818 => "00001010",2819 => "00010110",2820 => "10001101",2821 => "00010001",2822 => "10110010",2823 => "10010000",2824 => "00010000",2825 => "10011011",2826 => "10111101",2827 => "10110011",2828 => "10001010",2829 => "00100111",2830 => "10001000",2831 => "01000001",2832 => "10011111",2833 => "00001100",2834 => "01101000",2835 => "00011011",2836 => "11001101",2837 => "01100100",2838 => "11110100",2839 => "11011100",2840 => "11101001",2841 => "00101101",2842 => "11010101",2843 => "10011011",2844 => "10100101",2845 => "00110011",2846 => "00011010",2847 => "11110100",2848 => "10011100",2849 => "11110001",2850 => "11110010",2851 => "10010011",2852 => "00101001",2853 => "11111001",2854 => "00100101",2855 => "00011110",2856 => "01011100",2857 => "01110000",2858 => "11100100",2859 => "11000010",2860 => "10000101",2861 => "11100100",2862 => "11001100",2863 => "01110100",2864 => "11000000",2865 => "10111000",2866 => "10100111",2867 => "11010110",2868 => "11011111",2869 => "01100011",2870 => "01111100",2871 => "11010000",2872 => "11101100",2873 => "10110011",2874 => "11100010",2875 => "00101010",2876 => "11111110",2877 => "11111110",2878 => "00000011",2879 => "11111101",2880 => "11000001",2881 => "00001101",2882 => "11100001",2883 => "00111101",2884 => "11000110",2885 => "01111101",2886 => "01100111",2887 => "10100001",2888 => "01010000",2889 => "11011110",2890 => "01100010",2891 => "10001110",2892 => "00011100",2893 => "11100101",2894 => "01100000",2895 => "10000011",2896 => "01101001",2897 => "11111111",2898 => "01001001",2899 => "00110101",2900 => "01100000",2901 => "10111000",2902 => "00000110",2903 => "00100010",2904 => "00100101",2905 => "10110000",2906 => "10001001",2907 => "10011101",2908 => "10110110",2909 => "11011100",2910 => "00010011",2911 => "11100101",2912 => "00011110",2913 => "11100000",2914 => "01001000",2915 => "00101110",2916 => "10100101",2917 => "11010000",2918 => "01010100",2919 => "11001101",2920 => "01011000",2921 => "10111101",2922 => "11001000",2923 => "11011010",2924 => "11011000",2925 => "00010101",2926 => "10000101",2927 => "01011100",2928 => "11111111",2929 => "11011001",2930 => "11100000",2931 => "11111001",2932 => "10101111",2933 => "01110111",2934 => "01011000",2935 => "10000100",2936 => "10100101",2937 => "00001100",2938 => "01100011",2939 => "00110111",2940 => "11001101",2941 => "00101110",2942 => "01111101",2943 => "11101111",2944 => "11011000",2945 => "11000010",2946 => "10100111",2947 => "10100110",2948 => "01100011",2949 => "00001110",2950 => "01000110",2951 => "01011000",2952 => "10101110",2953 => "00100010",2954 => "01110100",2955 => "11011100",2956 => "11110100",2957 => "01011110",2958 => "10011001",2959 => "11010011",2960 => "10010010",2961 => "11110100",2962 => "00101010",2963 => "11011010",2964 => "11110101",2965 => "10111010",2966 => "11101011",2967 => "01110011",2968 => "10100101",2969 => "00111001",2970 => "11001000",2971 => "00001100",2972 => "01101000",2973 => "11101111",2974 => "01110011",2975 => "10011011",2976 => "10111100",2977 => "00110100",2978 => "11101000",2979 => "01101110",2980 => "11010100",2981 => "10001100",2982 => "00100011",2983 => "11101101",2984 => "01100111",2985 => "11001110",2986 => "01011011",2987 => "10001110",2988 => "01101001",2989 => "00010110",2990 => "10101101",2991 => "01110011",2992 => "01110000",2993 => "11101010",2994 => "00010111",2995 => "11110111",2996 => "00000011",2997 => "01110011",2998 => "11010111",2999 => "01110001",3000 => "01111011",3001 => "11101100",3002 => "00110111",3003 => "10110100",3004 => "00100011",3005 => "01111111",3006 => "01101000",3007 => "01011100",3008 => "00101010",3009 => "10111010",3010 => "11111100",3011 => "01010010",3012 => "01001101",3013 => "01001110",3014 => "11001100",3015 => "11101001",3016 => "10111000",3017 => "10111110",3018 => "01010110",3019 => "10001111",3020 => "01101010",3021 => "11011100",3022 => "00101110",3023 => "10010111",3024 => "11110101",3025 => "00111100",3026 => "10100001",3027 => "11110000",3028 => "00011101",3029 => "11111110",3030 => "11100110",3031 => "10001110",3032 => "01001001",3033 => "00011111",3034 => "00011101",3035 => "01111011",3036 => "01010001",3037 => "10111010",3038 => "01011101",3039 => "11100100",3040 => "01110010",3041 => "10100000",3042 => "11001110",3043 => "11001000",3044 => "00010000",3045 => "11001011",3046 => "00010110",3047 => "10000001",3048 => "10110010",3049 => "10100101",3050 => "00001011",3051 => "01111010",3052 => "00111000",3053 => "01011001",3054 => "00000100",3055 => "01000011",3056 => "11111100",3057 => "10101110",3058 => "01110011",3059 => "00101111",3060 => "01001011",3061 => "10110001",3062 => "10111000",3063 => "10010101",3064 => "01111010",3065 => "10111100",3066 => "11011101",3067 => "00110100",3068 => "11100000",3069 => "10000001",3070 => "01100001",3071 => "00011110",3072 => "10100010",3073 => "10110110",3074 => "00101110",3075 => "01101010",3076 => "00001101",3077 => "11110110",3078 => "10001010",3079 => "01010101",3080 => "10000010",3081 => "10011000",3082 => "11100011",3083 => "00010111",3084 => "00001000",3085 => "01100010",3086 => "01100101",3087 => "10110011",3088 => "11000010",3089 => "10011101",3090 => "10101110",3091 => "00110111",3092 => "11010101",3093 => "10111111",3094 => "01101010",3095 => "11111111",3096 => "00011000",3097 => "00110011",3098 => "00111100",3099 => "10101010",3100 => "10101000",3101 => "01100001",3102 => "01100101",3103 => "01111011",3104 => "00101101",3105 => "10111101",3106 => "11000101",3107 => "10000010",3108 => "00010001",3109 => "00100010",3110 => "01011100",3111 => "01110001",3112 => "01000011",3113 => "10101011",3114 => "11100010",3115 => "10010001",3116 => "11100010",3117 => "01000001",3118 => "11010000",3119 => "11101110",3120 => "01011100",3121 => "11010110",3122 => "10111111",3123 => "00111000",3124 => "10011101",3125 => "10000111",3126 => "01000101",3127 => "11111100",3128 => "00000111",3129 => "00011000",3130 => "11110111",3131 => "11101100",3132 => "11111100",3133 => "01001100",3134 => "11010000",3135 => "10110111",3136 => "10000101",3137 => "01101110",3138 => "01011011",3139 => "01100100",3140 => "11011000",3141 => "10111000",3142 => "00010110",3143 => "10000011",3144 => "01010000",3145 => "01000101",3146 => "00011010",3147 => "11110000",3148 => "00100011",3149 => "11001010",3150 => "11000010",3151 => "00111000",3152 => "10010100",3153 => "11100111",3154 => "10101001",3155 => "01000001",3156 => "00110000",3157 => "01011111",3158 => "10101011",3159 => "11110100",3160 => "11111000",3161 => "00101001",3162 => "10110010",3163 => "10110011",3164 => "11100100",3165 => "10101001",3166 => "10111011",3167 => "11111010",3168 => "11001111",3169 => "11111111",3170 => "01011100",3171 => "01001010",3172 => "00111111",3173 => "00100101",3174 => "10010000",3175 => "01101011",3176 => "00111010",3177 => "10000111",3178 => "10001111",3179 => "01000011",3180 => "01111110",3181 => "10111010",3182 => "11010110",3183 => "01100011",3184 => "11101011",3185 => "10011011",3186 => "01011010",3187 => "10110010",3188 => "01010110",3189 => "01010110",3190 => "00100110",3191 => "10100100",3192 => "01010110",3193 => "10101100",3194 => "01111001",3195 => "11000101",3196 => "10000010",3197 => "01001100",3198 => "11010000",3199 => "01111111",3200 => "00001110",3201 => "11001010",3202 => "01101011",3203 => "01001001",3204 => "10101110",3205 => "10001011",3206 => "00110100",3207 => "10111110",3208 => "10011101",3209 => "10101100",3210 => "10000000",3211 => "11001001",3212 => "11000101",3213 => "11011110",3214 => "01011000",3215 => "11101111",3216 => "10010001",3217 => "00100111",3218 => "10010111",3219 => "01010111",3220 => "11001000",3221 => "11011001",3222 => "11100110",3223 => "01101001",3224 => "10100110",3225 => "10100110",3226 => "11110110",3227 => "01000011",3228 => "00100011",3229 => "11011100",3230 => "00010101",3231 => "01100011",3232 => "00101011",3233 => "10010000",3234 => "11001111",3235 => "11110110",3236 => "11011010",3237 => "00111001",3238 => "00001000",3239 => "10101000",3240 => "00000011",3241 => "01100000",3242 => "01111001",3243 => "00101111",3244 => "01100001",3245 => "11011100",3246 => "01100100",3247 => "01010011",3248 => "11010100",3249 => "01110100",3250 => "10111011",3251 => "11000101",3252 => "11111110",3253 => "00101010",3254 => "11110011",3255 => "10010111",3256 => "01010010",3257 => "10001100",3258 => "10100100",3259 => "11100100",3260 => "00100100",3261 => "01111011",3262 => "01010110",3263 => "10100011",3264 => "10001000",3265 => "11001000",3266 => "01011011",3267 => "01010110",3268 => "00110000",3269 => "11100100",3270 => "10100000",3271 => "01110011",3272 => "01000101",3273 => "01001101",3274 => "11000110",3275 => "11001011",3276 => "10100001",3277 => "00001011",3278 => "10000011",3279 => "10011111",3280 => "00000110",3281 => "10100011",3282 => "01001111",3283 => "01100110",3284 => "01111101",3285 => "10111011",3286 => "01011001",3287 => "10010000",3288 => "00110110",3289 => "00011110",3290 => "10000000",3291 => "10000000",3292 => "10100001",3293 => "10011000",3294 => "10100100",3295 => "00001111",3296 => "01010100",3297 => "11010101",3298 => "10000100",3299 => "00111010",3300 => "11000101",3301 => "11001000",3302 => "00101100",3303 => "00111111",3304 => "01010111",3305 => "11100001",3306 => "00001011",3307 => "01101011",3308 => "11001000",3309 => "01101110",3310 => "01100011",3311 => "01010010",3312 => "00100011",3313 => "00110010",3314 => "01011101",3315 => "10010101",3316 => "11001010",3317 => "11000110",3318 => "10011011",3319 => "00000111",3320 => "00111010",3321 => "01110010",3322 => "00110001",3323 => "10111010",3324 => "11101010",3325 => "01001001",3326 => "01001000",3327 => "10111001",3328 => "00010011",3329 => "00111110",3330 => "11110001",3331 => "11101110",3332 => "11010001",3333 => "01010101",3334 => "10111110",3335 => "10101110",3336 => "10111101",3337 => "11000011",3338 => "10011111",3339 => "10010111",3340 => "00010110",3341 => "00001010",3342 => "00101111",3343 => "11010001",3344 => "11001000",3345 => "00000100",3346 => "00000001",3347 => "01111000",3348 => "11010001",3349 => "10111011",3350 => "01111010",3351 => "10110000",3352 => "00011010",3353 => "01110010",3354 => "01011110",3355 => "11101100",3356 => "11111000",3357 => "10011110",3358 => "01011011",3359 => "00100010",3360 => "00110111",3361 => "11111101",3362 => "01000101",3363 => "11001011",3364 => "01010000",3365 => "00011101",3366 => "01111000",3367 => "10100011",3368 => "10111111",3369 => "00111011",3370 => "10001001",3371 => "10000110",3372 => "00101000",3373 => "01001111",3374 => "01001100",3375 => "01101001",3376 => "11010000",3377 => "10101101",3378 => "10000001",3379 => "11101010",3380 => "01001010",3381 => "11100010",3382 => "11001011",3383 => "01100010",3384 => "00010001",3385 => "10001010",3386 => "00000001",3387 => "11000111",3388 => "01010100",3389 => "11010001",3390 => "00000111",3391 => "11111101",3392 => "01001100",3393 => "00010111",3394 => "01100100",3395 => "01001011",3396 => "10011101",3397 => "01101011",3398 => "01101111",3399 => "01000010",3400 => "00000011",3401 => "11101010",3402 => "10011100",3403 => "11100000",3404 => "01101010",3405 => "00011001",3406 => "00001101",3407 => "10110111",3408 => "11011110",3409 => "01010011",3410 => "10101001",3411 => "11010100",3412 => "00100001",3413 => "01011111",3414 => "01111011",3415 => "10000010",3416 => "10011010",3417 => "01101101",3418 => "11001101",3419 => "11010010",3420 => "00101000",3421 => "00111110",3422 => "01111011",3423 => "01010010",3424 => "11000000",3425 => "01100001",3426 => "10100110",3427 => "00011001",3428 => "01010011",3429 => "01000101",3430 => "10000101",3431 => "11010000",3432 => "11110110",3433 => "00110101",3434 => "10000001",3435 => "00001101",3436 => "01100111",3437 => "00011110",3438 => "00011100",3439 => "01001101",3440 => "11101100",3441 => "10000011",3442 => "01110101",3443 => "11000011",3444 => "01111100",3445 => "00101001",3446 => "00100100",3447 => "00000000",3448 => "11101011",3449 => "01101000",3450 => "11011101",3451 => "10001001",3452 => "11000001",3453 => "01111111",3454 => "00011010",3455 => "00100100",3456 => "00111010",3457 => "10011011",3458 => "01100001",3459 => "01111011",3460 => "10001010",3461 => "11110110",3462 => "10011111",3463 => "10110100",3464 => "01100100",3465 => "11111100",3466 => "00100110",3467 => "11100101",3468 => "10010001",3469 => "11110010",3470 => "01110111",3471 => "00011010",3472 => "10011110",3473 => "00011100",3474 => "00011011",3475 => "10011101",3476 => "11000110",3477 => "01110111",3478 => "11011111",3479 => "00000000",3480 => "11010100",3481 => "10101100",3482 => "10100011",3483 => "00111001",3484 => "10100100",3485 => "01011001",3486 => "01101000",3487 => "10000110",3488 => "11100000",3489 => "01001111",3490 => "01000110",3491 => "10001110",3492 => "10000111",3493 => "11010011",3494 => "11110001",3495 => "10101000",3496 => "00101110",3497 => "00100011",3498 => "10000000",3499 => "01011011",3500 => "00001110",3501 => "00101111",3502 => "00011001",3503 => "11111001",3504 => "10011100",3505 => "01111000",3506 => "11111100",3507 => "00111111",3508 => "11011100",3509 => "00001010",3510 => "01011110",3511 => "00101000",3512 => "01100010",3513 => "10100111",3514 => "00010110",3515 => "10100101",3516 => "11100100",3517 => "10110100",3518 => "00111010",3519 => "01010001",3520 => "00011000",3521 => "00111110",3522 => "11101010",3523 => "01010001",3524 => "11101011",3525 => "11000010",3526 => "11110100",3527 => "01000000",3528 => "00011011",3529 => "11101100",3530 => "11010000",3531 => "01101111",3532 => "01111010",3533 => "11111111",3534 => "00100101",3535 => "10100011",3536 => "11111101",3537 => "01011010",3538 => "10100011",3539 => "00101101",3540 => "01001111",3541 => "11100000",3542 => "11000000",3543 => "11111010",3544 => "11100110",3545 => "00010100",3546 => "11010111",3547 => "10010000",3548 => "10011100",3549 => "11111101",3550 => "10110110",3551 => "11000111",3552 => "10000101",3553 => "01111010",3554 => "01100001",3555 => "01001001",3556 => "10101100",3557 => "01010000",3558 => "00100000",3559 => "01110001",3560 => "10111101",3561 => "01010100",3562 => "01100010",3563 => "00111010",3564 => "00101101",3565 => "11110011",3566 => "11100011",3567 => "11101101",3568 => "10010110",3569 => "00010010",3570 => "01000110",3571 => "10101011",3572 => "10101100",3573 => "00101101",3574 => "10001101",3575 => "11011011",3576 => "10110111",3577 => "00000001",3578 => "10001010",3579 => "01001101",3580 => "00011011",3581 => "00000010",3582 => "00000010",3583 => "10000101",3584 => "00110000",3585 => "10010101",3586 => "10001001",3587 => "00001010",3588 => "10110111",3589 => "10001110",3590 => "10111010",3591 => "01100100",3592 => "01110011",3593 => "01101100",3594 => "10100110",3595 => "10101110",3596 => "11101011",3597 => "11000101",3598 => "10000000",3599 => "11101010",3600 => "00100010",3601 => "11001110",3602 => "11001111",3603 => "11000000",3604 => "01110110",3605 => "00111111",3606 => "01111111",3607 => "01110011",3608 => "01110100",3609 => "01101111",3610 => "10111011",3611 => "10111100",3612 => "00010110",3613 => "11101011",3614 => "00111111",3615 => "01000111",3616 => "01101111",3617 => "11101110",3618 => "01101000",3619 => "10110011",3620 => "11110001",3621 => "10011011",3622 => "10111001",3623 => "01010100",3624 => "10101111",3625 => "11100010",3626 => "01011010",3627 => "10111111",3628 => "00101001",3629 => "01111101",3630 => "01110101",3631 => "01010000",3632 => "00010010",3633 => "01101001",3634 => "10100011",3635 => "11011001",3636 => "10010100",3637 => "11100011",3638 => "00001010",3639 => "11000001",3640 => "01111001",3641 => "10001101",3642 => "11111000",3643 => "00100011",3644 => "01000100",3645 => "10101000",3646 => "00001011",3647 => "00000011",3648 => "00111010",3649 => "00010101",3650 => "10010101",3651 => "01000101",3652 => "01000001",3653 => "11011011",3654 => "11101010",3655 => "01110101",3656 => "11000000",3657 => "11001100",3658 => "11101111",3659 => "11111111",3660 => "01001010",3661 => "00101101",3662 => "10111110",3663 => "10000110",3664 => "10110100",3665 => "11010001",3666 => "10000111",3667 => "10111001",3668 => "00001010",3669 => "01011011",3670 => "01010100",3671 => "10010000",3672 => "10101011",3673 => "10100001",3674 => "01011000",3675 => "10010100",3676 => "00101011",3677 => "01100010",3678 => "11100101",3679 => "11100010",3680 => "00010110",3681 => "10101110",3682 => "10001100",3683 => "00001111",3684 => "10101111",3685 => "11011000",3686 => "00111101",3687 => "00011101",3688 => "01000100",3689 => "00111110",3690 => "00011011",3691 => "11101011",3692 => "00011111",3693 => "01100110",3694 => "00111101",3695 => "01111010",3696 => "01100110",3697 => "00011101",3698 => "11101011",3699 => "01111110",3700 => "00010000",3701 => "00110000",3702 => "10010101",3703 => "01010100",3704 => "00111111",3705 => "00110010",3706 => "11110011",3707 => "01101101",3708 => "01111100",3709 => "10111001",3710 => "00111110",3711 => "01001101",3712 => "01110000",3713 => "10110000",3714 => "00100011",3715 => "11011001",3716 => "00000010",3717 => "01111111",3718 => "01010101",3719 => "01001010",3720 => "00100010",3721 => "10111010",3722 => "10010101",3723 => "00001111",3724 => "11011000",3725 => "00101111",3726 => "00011101",3727 => "11000010",3728 => "11100100",3729 => "01111010",3730 => "01100011",3731 => "11111111",3732 => "11000110",3733 => "01000010",3734 => "11100000",3735 => "10111000",3736 => "00011010",3737 => "00010110",3738 => "00111011",3739 => "11111001",3740 => "00100101",3741 => "01100101",3742 => "10001000",3743 => "01001100",3744 => "10110100",3745 => "00011101",3746 => "00011010",3747 => "01110100",3748 => "10110011",3749 => "11011110",3750 => "11001110",3751 => "10001100",3752 => "01100000",3753 => "00111111",3754 => "01101100",3755 => "00101011",3756 => "01010110",3757 => "00011001",3758 => "01010101",3759 => "01000001",3760 => "11010110",3761 => "00111011",3762 => "10110011",3763 => "11111010",3764 => "00100100",3765 => "10111011",3766 => "01101111",3767 => "11111101",3768 => "01001110",3769 => "10111101",3770 => "00100001",3771 => "11001000",3772 => "11001110",3773 => "10111001",3774 => "00110100",3775 => "01111101",3776 => "00111111",3777 => "11100010",3778 => "01111110",3779 => "01100100",3780 => "10011010",3781 => "00110001",3782 => "10100111",3783 => "10010101",3784 => "11111111",3785 => "00100011",3786 => "10111011",3787 => "10111001",3788 => "11001011",3789 => "01010000",3790 => "11000001",3791 => "01100110",3792 => "10010000",3793 => "10011000",3794 => "00110010",3795 => "11111111",3796 => "01100110",3797 => "00100001",3798 => "01000111",3799 => "10010011",3800 => "01100101",3801 => "00010010",3802 => "11110000",3803 => "01011101",3804 => "01011111",3805 => "11000001",3806 => "10011100",3807 => "11101110",3808 => "11000001",3809 => "10010100",3810 => "11111000",3811 => "00010000",3812 => "10011101",3813 => "11111011",3814 => "11001011",3815 => "10111101",3816 => "10110110",3817 => "00000011",3818 => "10001011",3819 => "10000100",3820 => "10100100",3821 => "01000000",3822 => "01111001",3823 => "01011100",3824 => "11010111",3825 => "01001011",3826 => "10111111",3827 => "10110110",3828 => "01110011",3829 => "11110000",3830 => "10000101",3831 => "00110001",3832 => "11000101",3833 => "11101001",3834 => "01111010",3835 => "11001111",3836 => "00110010",3837 => "10101100",3838 => "01111110",3839 => "01011001",3840 => "10101100",3841 => "11011011",3842 => "01000010",3843 => "11101010",3844 => "10110000",3845 => "11001011",3846 => "01110011",3847 => "11000001",3848 => "01001101",3849 => "11110010",3850 => "01110010",3851 => "01111011",3852 => "00011111",3853 => "01011111",3854 => "11101000",3855 => "11101001",3856 => "10010101",3857 => "11001000",3858 => "10001110",3859 => "01111101",3860 => "00001111",3861 => "00100101",3862 => "00110101",3863 => "00111001",3864 => "10010010",3865 => "01000110",3866 => "10101000",3867 => "01111101",3868 => "00011001",3869 => "00111011",3870 => "01101110",3871 => "01000101",3872 => "00110011",3873 => "11010100",3874 => "10111000",3875 => "11110110",3876 => "00101000",3877 => "00101110",3878 => "00110000",3879 => "10011101",3880 => "01101111",3881 => "11101110",3882 => "10101001",3883 => "10011111",3884 => "00011111",3885 => "00010110",3886 => "10101100",3887 => "00110111",3888 => "00011000",3889 => "11111111",3890 => "01100111",3891 => "01100111",3892 => "00000111",3893 => "00110101",3894 => "00111101",3895 => "00111101",3896 => "11011101",3897 => "10110111",3898 => "00010100",3899 => "01011110",3900 => "01010011",3901 => "11101100",3902 => "01010001",3903 => "01001111",3904 => "10011000",3905 => "10101100",3906 => "10111110",3907 => "01101001",3908 => "01001111",3909 => "01001110",3910 => "00110000",3911 => "01100110",3912 => "10110100",3913 => "11001001",3914 => "00011001",3915 => "01011000",3916 => "00010101",3917 => "11110010",3918 => "01010101",3919 => "00101111",3920 => "01100001",3921 => "01100100",3922 => "00011000",3923 => "00000000",3924 => "10111001",3925 => "00010011",3926 => "10111010",3927 => "01001010",3928 => "11000110",3929 => "10111111",3930 => "11100001",3931 => "01000010",3932 => "11000110",3933 => "01010111",3934 => "10000000",3935 => "10001111",3936 => "00101100",3937 => "10001101",3938 => "11101011",3939 => "10001011",3940 => "00010010",3941 => "11111010",3942 => "01100100",3943 => "11001001",3944 => "10101010",3945 => "00100101",3946 => "10111101",3947 => "01011001",3948 => "01111001",3949 => "01000100",3950 => "11010000",3951 => "01011111",3952 => "11010010",3953 => "01011011",3954 => "11100101",3955 => "11110010",3956 => "11101000",3957 => "01000011",3958 => "11011111",3959 => "01111110",3960 => "11111111",3961 => "11110011",3962 => "01111101",3963 => "00000110",3964 => "10000100",3965 => "11001110",3966 => "00111111",3967 => "01111111",3968 => "10101010",3969 => "10001011",3970 => "00111000",3971 => "00011001",3972 => "01000000",3973 => "00011110",3974 => "01001100",3975 => "00100111",3976 => "00001001",3977 => "11111111",3978 => "00100110",3979 => "11011101",3980 => "00000100",3981 => "10110111",3982 => "11001100",3983 => "11001010",3984 => "10101011",3985 => "11000101",3986 => "11100010",3987 => "00100101",3988 => "01110001",3989 => "01100111",3990 => "10011110",3991 => "10111001",3992 => "01000101",3993 => "10001010",3994 => "10001110",3995 => "01100001",3996 => "10010010",3997 => "11110100",3998 => "11110110",3999 => "10101010",4000 => "11101101",4001 => "00000100",4002 => "11110100",4003 => "11011111",4004 => "10011000",4005 => "10011111",4006 => "00101110",4007 => "00011011",4008 => "01101101",4009 => "00010000",4010 => "11001100",4011 => "01111101",4012 => "00100111",4013 => "11001011",4014 => "11100101",4015 => "00100100",4016 => "00001101",4017 => "01110110",4018 => "10110100",4019 => "11001100",4020 => "00101010",4021 => "11000010",4022 => "10011000",4023 => "10000111",4024 => "11001000",4025 => "10100111",4026 => "01011100",4027 => "10001111",4028 => "00000101",4029 => "01110100",4030 => "00000100",4031 => "11010100",4032 => "11011100",4033 => "00101000",4034 => "01110101",4035 => "10010101",4036 => "10000101",4037 => "11111001",4038 => "11110011",4039 => "01011110",4040 => "00101011",4041 => "00011000",4042 => "00011011",4043 => "11100001",4044 => "10001001",4045 => "00101111",4046 => "11000110",4047 => "00011010",4048 => "10111100",4049 => "10100110",4050 => "01110010",4051 => "00110100",4052 => "00100110",4053 => "10011010",4054 => "01100101",4055 => "01010001",4056 => "10001011",4057 => "11111101",4058 => "01100011",4059 => "11000001",4060 => "10111001",4061 => "11111001",4062 => "11011011",4063 => "10100110",4064 => "11100011",4065 => "10010001",4066 => "10110110",4067 => "11100001",4068 => "11001111",4069 => "10000010",4070 => "01011010",4071 => "00010010",4072 => "10000010",4073 => "11101000",4074 => "10000000",4075 => "11100111",4076 => "01010101",4077 => "10101101",4078 => "00111111",4079 => "00111000",4080 => "01110011",4081 => "11010101",4082 => "11101011",4083 => "10100110",4084 => "01000001",4085 => "00100111",4086 => "00100100",4087 => "00110101",4088 => "11011001",4089 => "00111101",4090 => "10000001",4091 => "01000110",4092 => "01110110",4093 => "01100011",4094 => "10100001",4095 => "11011110",4096 => "01111010",4097 => "00111100",4098 => "11010000",4099 => "00000110",4100 => "11110001",4101 => "11100100",4102 => "00011011",4103 => "11111101",4104 => "10100011",4105 => "01111100",4106 => "11011010",4107 => "01110010",4108 => "11101000",4109 => "01011111",4110 => "10100010",4111 => "11011010",4112 => "10000111",4113 => "00110011",4114 => "01011010",4115 => "00001011",4116 => "11001100",4117 => "00110010",4118 => "11100101",4119 => "10100101",4120 => "01011111",4121 => "01011101",4122 => "00000111",4123 => "00001000",4124 => "11000101",4125 => "10011000",4126 => "11010001",4127 => "00000110",4128 => "01101000",4129 => "00011111",4130 => "01110000",4131 => "10100100",4132 => "01101100",4133 => "10011011",4134 => "11110100",4135 => "10100011",4136 => "11101001",4137 => "11010010",4138 => "01111111",4139 => "10010001",4140 => "10111100",4141 => "11100110",4142 => "00000111",4143 => "10000100",4144 => "00111110",4145 => "11010101",4146 => "01111011",4147 => "11011110",4148 => "01001110",4149 => "11010111",4150 => "10101001",4151 => "10000011",4152 => "01010111",4153 => "00000000",4154 => "01101011",4155 => "01011001",4156 => "00100110",4157 => "00011011",4158 => "01001000",4159 => "11111101",4160 => "11000110",4161 => "10101001",4162 => "10011011",4163 => "10111111",4164 => "11101011",4165 => "00101001",4166 => "00001011",4167 => "11110011",4168 => "01011001",4169 => "01111000",4170 => "01001001",4171 => "10011111",4172 => "11011001",4173 => "11011001",4174 => "01101011",4175 => "01011001",4176 => "01100110",4177 => "00011100",4178 => "00110011",4179 => "00100011",4180 => "00000101",4181 => "00001110",4182 => "00101111",4183 => "00011110",4184 => "10101110",4185 => "01010110",4186 => "00111101",4187 => "10000010",4188 => "00001010",4189 => "11001000",4190 => "01000111",4191 => "00110000",4192 => "11011000",4193 => "11100101",4194 => "11010001",4195 => "01110110",4196 => "00110111",4197 => "00101000",4198 => "01011001",4199 => "10111101",4200 => "11011100",4201 => "01011000",4202 => "11101010",4203 => "00011011",4204 => "11011000",4205 => "10101111",4206 => "00110110",4207 => "00001110",4208 => "10001000",4209 => "01001000",4210 => "00110010",4211 => "01011000",4212 => "10001011",4213 => "10101001",4214 => "01101110",4215 => "00001000",4216 => "00101010",4217 => "11110101",4218 => "00110000",4219 => "00010111",4220 => "10100001",4221 => "11010110",4222 => "11011011",4223 => "00000011",4224 => "10011001",4225 => "11101011",4226 => "11111011",4227 => "10110000",4228 => "00101101",4229 => "10000011",4230 => "01101000",4231 => "11101010",4232 => "10011100",4233 => "01010011",4234 => "00111111",4235 => "00101101",4236 => "01001011",4237 => "10111111",4238 => "11000110",4239 => "10001001",4240 => "01000000",4241 => "10110011",4242 => "00010101",4243 => "11100111",4244 => "00101100",4245 => "10011111",4246 => "01011001",4247 => "10110001",4248 => "00111010",4249 => "01100110",4250 => "00100100",4251 => "01101001",4252 => "00011110",4253 => "01110010",4254 => "01010110",4255 => "10111100",4256 => "10100100",4257 => "01001101",4258 => "11011111",4259 => "01010011",4260 => "11011001",4261 => "11100110",4262 => "00001111",4263 => "00000001",4264 => "01011111",4265 => "01100010",4266 => "10001010",4267 => "00010110",4268 => "01000001",4269 => "11010001",4270 => "10011100",4271 => "00100101",4272 => "00001100",4273 => "11011100",4274 => "11011100",4275 => "10010011",4276 => "00000100",4277 => "10000110",4278 => "00101101",4279 => "10111111",4280 => "01000101",4281 => "01101100",4282 => "11011110",4283 => "01011110",4284 => "11111111",4285 => "01010011",4286 => "11000011",4287 => "00111010",4288 => "01000000",4289 => "00011111",4290 => "00101011",4291 => "01110100",4292 => "10010100",4293 => "10000011",4294 => "00101010",4295 => "00101101",4296 => "00110110",4297 => "10010011",4298 => "10011011",4299 => "01011101",4300 => "10011011",4301 => "00110000",4302 => "01100010",4303 => "10100001",4304 => "00101110",4305 => "11111001",4306 => "01110000",4307 => "10001001",4308 => "11111101",4309 => "11111001",4310 => "10001010",4311 => "10001110",4312 => "11100100",4313 => "10110010",4314 => "11111010",4315 => "01101010",4316 => "11111110",4317 => "00010110",4318 => "10001101",4319 => "11011101",4320 => "00110001",4321 => "10010101",4322 => "01100111",4323 => "01001111",4324 => "00100011",4325 => "11110000",4326 => "10100101",4327 => "00111100",4328 => "00100000",4329 => "11011100",4330 => "11001100",4331 => "10010111",4332 => "10011110",4333 => "01000110",4334 => "01000110",4335 => "11001110",4336 => "01101111",4337 => "00101110",4338 => "00000001",4339 => "00011100",4340 => "10000111",4341 => "11101100",4342 => "01101011",4343 => "11001100",4344 => "10011100",4345 => "10001110",4346 => "00110111",4347 => "11101101",4348 => "00110111",4349 => "11000011",4350 => "01101100",4351 => "10000110",4352 => "00000001",4353 => "11100110",4354 => "11101110",4355 => "11110010",4356 => "10001010",4357 => "01001100",4358 => "11001000",4359 => "11010110",4360 => "00000111",4361 => "10001110",4362 => "11101000",4363 => "00111000",4364 => "10010100",4365 => "10100010",4366 => "01001111",4367 => "10111101",4368 => "00000110",4369 => "10100010",4370 => "00010010",4371 => "00110111",4372 => "00100011",4373 => "00101111",4374 => "10001111",4375 => "00111111",4376 => "01001101",4377 => "00011001",4378 => "00111110",4379 => "11111010",4380 => "11111100",4381 => "01110111",4382 => "00110011",4383 => "01100011",4384 => "11010000",4385 => "11101111",4386 => "01011110",4387 => "10010110",4388 => "11000000",4389 => "01111100",4390 => "11001110",4391 => "00111000",4392 => "01011101",4393 => "11111100",4394 => "10001000",4395 => "10111111",4396 => "10011011",4397 => "01111101",4398 => "11101110",4399 => "10101110",4400 => "00010011",4401 => "01110000",4402 => "01000111",4403 => "10110000",4404 => "11101101",4405 => "00100000",4406 => "01000100",4407 => "11111011",4408 => "01101011",4409 => "00111100",4410 => "00101011",4411 => "11000101",4412 => "11000110",4413 => "01110100",4414 => "11011011",4415 => "00101000",4416 => "10000000",4417 => "10110010",4418 => "00001100",4419 => "11101001",4420 => "11010100",4421 => "10110110",4422 => "10110000",4423 => "01110011",4424 => "01001010",4425 => "10101001",4426 => "01011101",4427 => "10111001",4428 => "00010101",4429 => "01010000",4430 => "00001010",4431 => "10100000",4432 => "00111110",4433 => "11010010",4434 => "10011011",4435 => "00000110",4436 => "00101111",4437 => "10000000",4438 => "00111100",4439 => "01111010",4440 => "00100011",4441 => "10010000",4442 => "11011001",4443 => "01001001",4444 => "11111111",4445 => "10000111",4446 => "10101001",4447 => "11010101",4448 => "11000100",4449 => "10000110",4450 => "11010101",4451 => "10010111",4452 => "01100100",4453 => "01110011",4454 => "01011010",4455 => "11001110",4456 => "11010111",4457 => "11010101",4458 => "11111000",4459 => "11110001",4460 => "10100101",4461 => "00110111",4462 => "00110110",4463 => "01110011",4464 => "00000000",4465 => "11010001",4466 => "11100011",4467 => "01001010",4468 => "00001100",4469 => "01110011",4470 => "01011000",4471 => "01100111",4472 => "00110111",4473 => "11111001",4474 => "11110011",4475 => "01101011",4476 => "10001110",4477 => "10101001",4478 => "11001101",4479 => "01011010",4480 => "11000101",4481 => "11011000",4482 => "00010011",4483 => "11000111",4484 => "10001110",4485 => "00101010",4486 => "11000001",4487 => "01000011",4488 => "01100100",4489 => "00100000",4490 => "10110111",4491 => "10110000",4492 => "11001001",4493 => "11111010",4494 => "00101100",4495 => "10111011",4496 => "11101111",4497 => "00000011",4498 => "10001101",4499 => "10011000",4500 => "01011100",4501 => "10110100",4502 => "01100111",4503 => "00010001",4504 => "01000011",4505 => "10101011",4506 => "01010011",4507 => "01101011",4508 => "10010000",4509 => "11100011",4510 => "10011001",4511 => "11010010",4512 => "11101011",4513 => "01011010",4514 => "00000011",4515 => "00110011",4516 => "11010011",4517 => "00010001",4518 => "11100110",4519 => "11000111",4520 => "11100110",4521 => "01000011",4522 => "10000010",4523 => "10001110",4524 => "01100100",4525 => "00010000",4526 => "10011110",4527 => "01111110",4528 => "10000101",4529 => "01100010",4530 => "11010000",4531 => "01000110",4532 => "00001010",4533 => "00011001",4534 => "11001111",4535 => "11011111",4536 => "00101001",4537 => "10101111",4538 => "00000101",4539 => "01010101",4540 => "11011010",4541 => "11000011",4542 => "01111000",4543 => "00101100",4544 => "11100001",4545 => "10110000",4546 => "00010100",4547 => "11001101",4548 => "00111010",4549 => "11100100",4550 => "01000111",4551 => "00000010",4552 => "11110000",4553 => "11010101",4554 => "01001101",4555 => "00011000",4556 => "00111011",4557 => "10110011",4558 => "01011111",4559 => "00000010",4560 => "01100101",4561 => "10011010",4562 => "10111110",4563 => "10001111",4564 => "11100110",4565 => "00010011",4566 => "01100100",4567 => "10001010",4568 => "11010111",4569 => "11001100",4570 => "11011010",4571 => "11100011",4572 => "10101000",4573 => "11101010",4574 => "01010011",4575 => "11111111",4576 => "11001011",4577 => "00001101",4578 => "10001011",4579 => "00100101",4580 => "10100110",4581 => "11000001",4582 => "10000010",4583 => "10101001",4584 => "10010010",4585 => "11010100",4586 => "11011000",4587 => "00101000",4588 => "10010110",4589 => "01000100",4590 => "00110000",4591 => "01100111",4592 => "01101000",4593 => "01011011",4594 => "11010001",4595 => "11111101",4596 => "10010000",4597 => "00100111",4598 => "01110000",4599 => "01100100",4600 => "01110010",4601 => "11000001",4602 => "10111010",4603 => "10011111",4604 => "11010011",4605 => "10011100",4606 => "01001100",4607 => "10011101",4608 => "01110111",4609 => "00010100",4610 => "01010011",4611 => "00111111",4612 => "00110001",4613 => "01101111",4614 => "10001100",4615 => "00100001",4616 => "11111000",4617 => "00010100",4618 => "11111000",4619 => "01111101",4620 => "01010001",4621 => "10100111",4622 => "11010110",4623 => "10111000",4624 => "01110111",4625 => "11001000",4626 => "01001101",4627 => "01111101",4628 => "01010111",4629 => "10110101",4630 => "11000000",4631 => "11001111",4632 => "11011000",4633 => "01010100",4634 => "00101100",4635 => "10010001",4636 => "11000011",4637 => "11101110",4638 => "01110110",4639 => "01000011",4640 => "10011100",4641 => "11010010",4642 => "11100010",4643 => "01111101",4644 => "10011110",4645 => "10110000",4646 => "11101100",4647 => "10101100",4648 => "11111111",4649 => "10010011",4650 => "11001101",4651 => "10011111",4652 => "10101110",4653 => "01100000",4654 => "00101001",4655 => "00010101",4656 => "10011001",4657 => "01001001",4658 => "10010010",4659 => "10011101",4660 => "00100011",4661 => "01101010",4662 => "10100000",4663 => "10101010",4664 => "11010011",4665 => "01100100",4666 => "01010101",4667 => "01111100",4668 => "00001000",4669 => "10100000",4670 => "01111011",4671 => "00011101",4672 => "01111110",4673 => "01000110",4674 => "00111010",4675 => "00110101",4676 => "10001011",4677 => "11011010",4678 => "00100101",4679 => "00101011",4680 => "10001101",4681 => "11001001",4682 => "11001101",4683 => "01111100",4684 => "01000101",4685 => "10001001",4686 => "11001101",4687 => "00000000",4688 => "11010101",4689 => "01011001",4690 => "11100110",4691 => "10110000",4692 => "11011010",4693 => "01111000",4694 => "10010100",4695 => "01000001",4696 => "01110000",4697 => "11011101",4698 => "11010010",4699 => "00110110",4700 => "00010011",4701 => "10001001",4702 => "01101101",4703 => "11010100",4704 => "11100101",4705 => "01001100",4706 => "00010010",4707 => "11111001",4708 => "01110111",4709 => "01000111",4710 => "10010100",4711 => "11011110",4712 => "01101001",4713 => "11110111",4714 => "11110110",4715 => "10111111",4716 => "10101011",4717 => "10101010",4718 => "01010011",4719 => "01110011",4720 => "11111000",4721 => "11101100",4722 => "10000011",4723 => "11111011",4724 => "10110010",4725 => "00010110",4726 => "11010010",4727 => "01110111",4728 => "00001011",4729 => "01001111",4730 => "00000000",4731 => "11100001",4732 => "00011100",4733 => "11011000",4734 => "01110011",4735 => "01111000",4736 => "11001100",4737 => "11111011",4738 => "01100011",4739 => "00110110",4740 => "10001001",4741 => "00101010",4742 => "11011010",4743 => "11010011",4744 => "00100010",4745 => "00011000",4746 => "11011001",4747 => "10110000",4748 => "10111111",4749 => "01001100",4750 => "10011110",4751 => "00111101",4752 => "11101000",4753 => "10110000",4754 => "01111010",4755 => "00100100",4756 => "01111110",4757 => "00111010",4758 => "00010001",4759 => "00010011",4760 => "11010001",4761 => "01010111",4762 => "10000010",4763 => "00000001",4764 => "10001111",4765 => "01000000",4766 => "00010001",4767 => "01010010",4768 => "00110011",4769 => "00000111",4770 => "00000101",4771 => "11001111",4772 => "01100011",4773 => "01000100",4774 => "00111100",4775 => "11111010",4776 => "00101000",4777 => "01101101",4778 => "11000010",4779 => "00101100",4780 => "01000000",4781 => "10111010",4782 => "00110111",4783 => "11110011",4784 => "00110001",4785 => "11101000",4786 => "00001011",4787 => "11010010",4788 => "11010010",4789 => "11101000",4790 => "10111011",4791 => "10010000",4792 => "01110000",4793 => "01100001",4794 => "11111010",4795 => "00011101",4796 => "01010011",4797 => "00110110",4798 => "11011111",4799 => "11110111",4800 => "00011010",4801 => "01011000",4802 => "11011010",4803 => "01100110",4804 => "11000111",4805 => "00000001",4806 => "00101001",4807 => "01010111",4808 => "01011011",4809 => "00010111",4810 => "10111101",4811 => "10100010",4812 => "11010100",4813 => "11001100",4814 => "10000011",4815 => "10100001",4816 => "00101111",4817 => "00001010",4818 => "01100010",4819 => "01011000",4820 => "10101110",4821 => "00011001",4822 => "00001001",4823 => "01001011",4824 => "11111100",4825 => "11010100",4826 => "10100010",4827 => "11100110",4828 => "11010001",4829 => "00000100",4830 => "00000110",4831 => "01110011",4832 => "11010101",4833 => "10010101",4834 => "00100011",4835 => "11001111",4836 => "10010001",4837 => "11001001",4838 => "11010000",4839 => "00111010",4840 => "00100111",4841 => "11000100",4842 => "10111101",4843 => "01100111",4844 => "01101011",4845 => "10101111",4846 => "00011110",4847 => "01010101",4848 => "11111111",4849 => "00001001",4850 => "01010010",4851 => "00000001",4852 => "01000111",4853 => "11001100",4854 => "01001010",4855 => "00011111",4856 => "11010101",4857 => "10111000",4858 => "10111111",4859 => "00011011",4860 => "10100100",4861 => "11010100",4862 => "11000110",4863 => "01011001",4864 => "11110110",4865 => "10000000",4866 => "11100000",4867 => "00010000",4868 => "01001100",4869 => "10110100",4870 => "10110001",4871 => "11101111",4872 => "01111110",4873 => "10011010",4874 => "10101110",4875 => "10011010",4876 => "10000011",4877 => "10001011",4878 => "00111110",4879 => "01011001",4880 => "00101101",4881 => "01000110",4882 => "11100101",4883 => "01111100",4884 => "00010010",4885 => "11011101",4886 => "01110101",4887 => "11111100",4888 => "10110101",4889 => "01111011",4890 => "01001011",4891 => "00010011",4892 => "00111001",4893 => "01101101",4894 => "10110001",4895 => "01000001",4896 => "01110101",4897 => "01111100",4898 => "01000000",4899 => "01100010",4900 => "11000101",4901 => "10111011",4902 => "10011100",4903 => "11111011",4904 => "11110001",4905 => "00011001",4906 => "01010110",4907 => "10001010",4908 => "00010011",4909 => "00010111",4910 => "01010111",4911 => "11000000",4912 => "00110100",4913 => "01000001",4914 => "01000011",4915 => "01011101",4916 => "01111101",4917 => "01101001",4918 => "01110110",4919 => "01101000",4920 => "10001001",4921 => "01101100",4922 => "10010011",4923 => "11100010",4924 => "11000100",4925 => "01110101",4926 => "11001100",4927 => "00110101",4928 => "11001000",4929 => "00101100",4930 => "00000001",4931 => "10011001",4932 => "11101000",4933 => "11101010",4934 => "11110100",4935 => "00010111",4936 => "01110011",4937 => "10110100",4938 => "11011011",4939 => "01001011",4940 => "10001011",4941 => "01110101",4942 => "01000111",4943 => "11100001",4944 => "11110101",4945 => "10000111",4946 => "11001010",4947 => "10110110",4948 => "11100101",4949 => "00101001",4950 => "11110111",4951 => "00010101",4952 => "10000000",4953 => "11111011",4954 => "01001100",4955 => "00110011",4956 => "11010001",4957 => "00101010",4958 => "01110001",4959 => "01010100",4960 => "11000011",4961 => "11101110",4962 => "00010001",4963 => "10001110",4964 => "00101001",4965 => "01111001",4966 => "11101010",4967 => "01000010",4968 => "10111011",4969 => "11101101",4970 => "01100101",4971 => "11100011",4972 => "10110100",4973 => "00111011",4974 => "11101011",4975 => "10001000",4976 => "10000111",4977 => "11110110",4978 => "11111101",4979 => "10100000",4980 => "00111001",4981 => "11110111",4982 => "10111110",4983 => "10000110",4984 => "00010011",4985 => "01100010",4986 => "00000001",4987 => "00010001",4988 => "10100011",4989 => "01101101",4990 => "01100100",4991 => "01110111",4992 => "00100011",4993 => "10011000",4994 => "11001101",4995 => "00111011",4996 => "11100001",4997 => "11111110",4998 => "00101101",4999 => "11110100",5000 => "10001101",5001 => "10100110",5002 => "10111011",5003 => "01010101",5004 => "01111101",5005 => "00000100",5006 => "01001010",5007 => "00100010",5008 => "10101000",5009 => "10100100",5010 => "11111101",5011 => "00110000",5012 => "10011101",5013 => "10001101",5014 => "11111000",5015 => "01111001",5016 => "10001111",5017 => "11000001",5018 => "10001001",5019 => "01100010",5020 => "00011111",5021 => "10101001",5022 => "00001010",5023 => "11111110",5024 => "11000000",5025 => "10000110",5026 => "01111000",5027 => "11110100",5028 => "10101011",5029 => "00100101",5030 => "00100111",5031 => "10100010",5032 => "10100001",5033 => "11110101",5034 => "10011000",5035 => "01000011",5036 => "10101011",5037 => "01010100",5038 => "01110001",5039 => "00100100",5040 => "11111011",5041 => "10110101",5042 => "11101010",5043 => "00000010",5044 => "01001100",5045 => "00010111",5046 => "00000011",5047 => "01100110",5048 => "10000111",5049 => "11010010",5050 => "11110111",5051 => "01010110",5052 => "10000000",5053 => "11110000",5054 => "11011100",5055 => "10010001",5056 => "00011110",5057 => "11001010",5058 => "00101000",5059 => "00100001",5060 => "11100100",5061 => "01111000",5062 => "00011001",5063 => "10000001",5064 => "10110000",5065 => "11011100",5066 => "00111011",5067 => "11101011",5068 => "10011111",5069 => "00011000",5070 => "01110000",5071 => "11010110",5072 => "10111101",5073 => "11010110",5074 => "00110011",5075 => "00110110",5076 => "01000010",5077 => "00000110",5078 => "10000000",5079 => "00010001",5080 => "01001101",5081 => "11000001",5082 => "10010111",5083 => "10101110",5084 => "11010110",5085 => "01001101",5086 => "01010111",5087 => "10001111",5088 => "10001111",5089 => "11010100",5090 => "01000111",5091 => "11100010",5092 => "01010111",5093 => "00110010",5094 => "01001110",5095 => "11000010",5096 => "11011011",5097 => "00111111",5098 => "11110011",5099 => "01100001",5100 => "01110101",5101 => "11001010",5102 => "01111100",5103 => "00011110",5104 => "11011001",5105 => "00111101",5106 => "01100110",5107 => "11110010",5108 => "00011101",5109 => "00000001",5110 => "01001010",5111 => "00101100",5112 => "00111101",5113 => "00001111",5114 => "00010000",5115 => "11010111",5116 => "01010101",5117 => "01000111",5118 => "10011100",5119 => "10010000",5120 => "11100101",5121 => "01001000",5122 => "00001000",5123 => "11011010",5124 => "10101111",5125 => "11000110",5126 => "11011001",5127 => "00110000",5128 => "10110010",5129 => "11000001",5130 => "11010101",5131 => "10101110",5132 => "10110111",5133 => "00001101",5134 => "01111111",5135 => "01110101",5136 => "01000100",5137 => "11001010",5138 => "01011011",5139 => "10100001",5140 => "10011111",5141 => "00110101",5142 => "01101011",5143 => "01100100",5144 => "11001110",5145 => "00101100",5146 => "10101101",5147 => "01100001",5148 => "00010101",5149 => "01110010",5150 => "01110111",5151 => "11010100",5152 => "10001110",5153 => "01101101",5154 => "00001100",5155 => "00001101",5156 => "00010000",5157 => "10101101",5158 => "11011101",5159 => "01011110",5160 => "00110111",5161 => "10001001",5162 => "00111001",5163 => "10101100",5164 => "01111101",5165 => "10110000",5166 => "10111001",5167 => "10100101",5168 => "11010001",5169 => "00010000",5170 => "11011100",5171 => "11111001",5172 => "01010001",5173 => "00101100",5174 => "01101100",5175 => "11111101",5176 => "10100110",5177 => "01111011",5178 => "11101111",5179 => "01111100",5180 => "11010111",5181 => "10101010",5182 => "00110000",5183 => "00101101",5184 => "01000100",5185 => "10001000",5186 => "10110001",5187 => "11001000",5188 => "11100001",5189 => "00111100",5190 => "01110110",5191 => "01000100",5192 => "00001000",5193 => "10110101",5194 => "00011011",5195 => "10110001",5196 => "01100010",5197 => "10111100",5198 => "10000001",5199 => "10001110",5200 => "11001010",5201 => "11010010",5202 => "11101110",5203 => "00011111",5204 => "01100001",5205 => "10111101",5206 => "10101111",5207 => "10111000",5208 => "10011110",5209 => "10000111",5210 => "10111001",5211 => "01111011",5212 => "10110100",5213 => "10001010",5214 => "11110111",5215 => "01110010",5216 => "00000000",5217 => "10011101",5218 => "11001001",5219 => "00001010",5220 => "11111110",5221 => "01000110",5222 => "01101100",5223 => "11100010",5224 => "01010101",5225 => "11010001",5226 => "01011000",5227 => "10110101",5228 => "11001011",5229 => "01000011",5230 => "01111011",5231 => "11000000",5232 => "10000001",5233 => "00111011",5234 => "10101111",5235 => "11111011",5236 => "10100101",5237 => "01001000",5238 => "00101011",5239 => "01100100",5240 => "11010010",5241 => "00001100",5242 => "10000100",5243 => "01110011",5244 => "11000100",5245 => "01000101",5246 => "11001000",5247 => "00111110",5248 => "11100111",5249 => "10001001",5250 => "11101001",5251 => "10000001",5252 => "01111100",5253 => "01000011",5254 => "00100010",5255 => "11100100",5256 => "01110100",5257 => "00000101",5258 => "11100111",5259 => "00100010",5260 => "01001101",5261 => "00101000",5262 => "10100010",5263 => "01111110",5264 => "11101101",5265 => "11010111",5266 => "01000100",5267 => "11000111",5268 => "10111001",5269 => "00101010",5270 => "10100000",5271 => "10001001",5272 => "01011001",5273 => "00010011",5274 => "11101110",5275 => "10111000",5276 => "11100001",5277 => "10001101",5278 => "11101101",5279 => "00101001",5280 => "10111010",5281 => "11111100",5282 => "11101001",5283 => "11010001",5284 => "01110010",5285 => "11111000",5286 => "00001100",5287 => "00000111",5288 => "11101111",5289 => "10011100",5290 => "11010110",5291 => "10110111",5292 => "00110000",5293 => "01100010",5294 => "11011001",5295 => "10111000",5296 => "11101000",5297 => "11101001",5298 => "10100000",5299 => "11110111",5300 => "10000010",5301 => "01010111",5302 => "01000110",5303 => "00000110",5304 => "11111111",5305 => "01011101",5306 => "00000100",5307 => "10110110",5308 => "10011010",5309 => "00110011",5310 => "11001111",5311 => "11110100",5312 => "00101111",5313 => "00100111",5314 => "10100000",5315 => "00000001",5316 => "00100110",5317 => "10100010",5318 => "01011000",5319 => "00111000",5320 => "01101000",5321 => "01001111",5322 => "11010000",5323 => "10000010",5324 => "00010100",5325 => "11101000",5326 => "11011001",5327 => "00111100",5328 => "00110110",5329 => "00000101",5330 => "01000001",5331 => "11011110",5332 => "10011010",5333 => "01000001",5334 => "00101101",5335 => "11010010",5336 => "00011010",5337 => "10010001",5338 => "00101011",5339 => "00001101",5340 => "01111100",5341 => "00000101",5342 => "00011010",5343 => "01010111",5344 => "11010001",5345 => "00111001",5346 => "11100111",5347 => "01110110",5348 => "00101101",5349 => "10001110",5350 => "00001000",5351 => "01001110",5352 => "00000001",5353 => "01001100",5354 => "11001011",5355 => "10110100",5356 => "10001100",5357 => "01111111",5358 => "10001010",5359 => "00000111",5360 => "11111110",5361 => "10110010",5362 => "11100110",5363 => "10001001",5364 => "00010011",5365 => "10101100",5366 => "10010001",5367 => "10010001",5368 => "10100011",5369 => "10111001",5370 => "11010100",5371 => "01011110",5372 => "01001000",5373 => "10010010",5374 => "10001011",5375 => "11110111",5376 => "01111110",5377 => "01001001",5378 => "01111101",5379 => "00010000",5380 => "11101111",5381 => "11110111",5382 => "11111001",5383 => "10111101",5384 => "01101001",5385 => "01100100",5386 => "11110000",5387 => "10101010",5388 => "11100001",5389 => "10100100",5390 => "00011110",5391 => "11011000",5392 => "00100000",5393 => "01000110",5394 => "00001111",5395 => "01001100",5396 => "00110000",5397 => "11010010",5398 => "00100011",5399 => "11000100",5400 => "11101000",5401 => "01001010",5402 => "00000100",5403 => "01001111",5404 => "00011110",5405 => "00011101",5406 => "01010100",5407 => "10011000",5408 => "01101011",5409 => "00101000",5410 => "10100101",5411 => "00011011",5412 => "00000101",5413 => "11011010",5414 => "11011100",5415 => "01010100",5416 => "00101011",5417 => "01010010",5418 => "11010010",5419 => "00111001",5420 => "01000101",5421 => "00001010",5422 => "01100010",5423 => "10111111",5424 => "01110000",5425 => "11111001",5426 => "01001010",5427 => "00010000",5428 => "10110100",5429 => "10110010",5430 => "00000001",5431 => "10001110",5432 => "11011111",5433 => "10100001",5434 => "00011111",5435 => "11111110",5436 => "11110010",5437 => "01100110",5438 => "01111000",5439 => "01100111",5440 => "01111101",5441 => "01010001",5442 => "10100100",5443 => "01110101",5444 => "11100100",5445 => "10111011",5446 => "00100100",5447 => "01010000",5448 => "10100000",5449 => "11010000",5450 => "01100010",5451 => "10110110",5452 => "11101110",5453 => "10100001",5454 => "00101010",5455 => "01110010",5456 => "01110010",5457 => "11001011",5458 => "10011101",5459 => "00111010",5460 => "10000011",5461 => "10010000",5462 => "10101101",5463 => "10111010",5464 => "10001000",5465 => "10011110",5466 => "10000001",5467 => "01111011",5468 => "01101110",5469 => "00111011",5470 => "10000001",5471 => "01111101",5472 => "01000011",5473 => "00101100",5474 => "01011100",5475 => "01111110",5476 => "10101101",5477 => "10000101",5478 => "00000010",5479 => "11111011",5480 => "00001010",5481 => "10001000",5482 => "00001101",5483 => "01101110",5484 => "10000000",5485 => "11011101",5486 => "10100111",5487 => "10010111",5488 => "11110111",5489 => "11001101",5490 => "10011000",5491 => "10010000",5492 => "11001111",5493 => "01001111",5494 => "01100100",5495 => "11101100",5496 => "00001100",5497 => "10100100",5498 => "10011000",5499 => "11011000",5500 => "01110111",5501 => "10011111",5502 => "11101001",5503 => "01010010",5504 => "11100001",5505 => "01001111",5506 => "01000000",5507 => "11101001",5508 => "00100001",5509 => "00101101",5510 => "10001100",5511 => "11001010",5512 => "10101000",5513 => "01011000",5514 => "11010101",5515 => "10001101",5516 => "10011010",5517 => "10010111",5518 => "11110111",5519 => "10011000",5520 => "11011011",5521 => "11100011",5522 => "01000010",5523 => "11010101",5524 => "00111101",5525 => "01111110",5526 => "00001001",5527 => "00101011",5528 => "00010110",5529 => "11001001",5530 => "10010100",5531 => "11010101",5532 => "01100000",5533 => "11010110",5534 => "00000101",5535 => "11000011",5536 => "01001000",5537 => "01001101",5538 => "11011010",5539 => "11100010",5540 => "01111010",5541 => "11110001",5542 => "01010011",5543 => "11010110",5544 => "10010000",5545 => "10110011",5546 => "10001001",5547 => "00010000",5548 => "11011001",5549 => "10010010",5550 => "11100011",5551 => "00010110",5552 => "01100010",5553 => "00011111",5554 => "00100110",5555 => "11001011",5556 => "11101011",5557 => "01010011",5558 => "00111011",5559 => "11110010",5560 => "01110011",5561 => "11101000",5562 => "00001111",5563 => "01110111",5564 => "11010110",5565 => "00111101",5566 => "11011001",5567 => "00010011",5568 => "10000101",5569 => "01001101",5570 => "00011111",5571 => "11001101",5572 => "00101110",5573 => "11101110",5574 => "00011101",5575 => "11110001",5576 => "10010010",5577 => "01001001",5578 => "01100001",5579 => "01110000",5580 => "00100011",5581 => "01110011",5582 => "00100010",5583 => "10010011",5584 => "10110111",5585 => "00110000",5586 => "01011000",5587 => "01000011",5588 => "10000001",5589 => "00111000",5590 => "10010011",5591 => "00010011",5592 => "10101000",5593 => "01110000",5594 => "01001100",5595 => "11101011",5596 => "11111101",5597 => "00001010",5598 => "11101011",5599 => "01101110",5600 => "10011101",5601 => "01110010",5602 => "10110101",5603 => "11111011",5604 => "00000101",5605 => "00011000",5606 => "00111000",5607 => "11000000",5608 => "11101111",5609 => "10001100",5610 => "01100111",5611 => "11101011",5612 => "01000011",5613 => "10001101",5614 => "10011100",5615 => "10101001",5616 => "11001101",5617 => "00111011",5618 => "11101001",5619 => "00111011",5620 => "01001011",5621 => "11100100",5622 => "01100110",5623 => "10001101",5624 => "11010101",5625 => "00101100",5626 => "11111001",5627 => "10011111",5628 => "00011110",5629 => "00000001",5630 => "00010010",5631 => "11011001",5632 => "01101011",5633 => "10101001",5634 => "01101100",5635 => "01111111",5636 => "11100100",5637 => "01010011",5638 => "01110011",5639 => "11110111",5640 => "11110001",5641 => "00010111",5642 => "01010001",5643 => "01001110",5644 => "10000101",5645 => "01010001",5646 => "10011010",5647 => "10100001",5648 => "11010000",5649 => "11000001",5650 => "01011110",5651 => "01011100",5652 => "01011001",5653 => "01100101",5654 => "00010101",5655 => "01101101",5656 => "01111000",5657 => "10111100",5658 => "11010001",5659 => "10011001",5660 => "11000000",5661 => "01111101",5662 => "01100101",5663 => "10101110",5664 => "10101010",5665 => "11100000",5666 => "10100110",5667 => "10111001",5668 => "00000001",5669 => "11101110",5670 => "10110111",5671 => "10011001",5672 => "11001100",5673 => "00111110",5674 => "10001110",5675 => "00001000",5676 => "00111101",5677 => "00011000",5678 => "11011011",5679 => "00011000",5680 => "10110110",5681 => "10011011",5682 => "00011100",5683 => "01010100",5684 => "00000000",5685 => "10101101",5686 => "00010110",5687 => "10011000",5688 => "10001101",5689 => "10000100",5690 => "11101001",5691 => "01001010",5692 => "01000110",5693 => "10001010",5694 => "10010101",5695 => "01110101",5696 => "10010010",5697 => "11100011",5698 => "01100111",5699 => "00101000",5700 => "00000100",5701 => "00101101",5702 => "10111001",5703 => "10100010",5704 => "10111100",5705 => "00111101",5706 => "01101111",5707 => "01110101",5708 => "01111001",5709 => "11011101",5710 => "00111010",5711 => "10101111",5712 => "01110111",5713 => "00110110",5714 => "10011111",5715 => "10001000",5716 => "01001000",5717 => "11000010",5718 => "10010101",5719 => "11101001",5720 => "10100110",5721 => "11011110",5722 => "11110110",5723 => "01101001",5724 => "00100101",5725 => "00011011",5726 => "00101001",5727 => "01110010",5728 => "11111001",5729 => "00100110",5730 => "01001100",5731 => "00101010",5732 => "11001101",5733 => "11001011",5734 => "10101010",5735 => "11111000",5736 => "00000001",5737 => "01100100",5738 => "10100101",5739 => "01001111",5740 => "10001101",5741 => "00111010",5742 => "00000100",5743 => "11100001",5744 => "11101100",5745 => "01000111",5746 => "01100100",5747 => "10111000",5748 => "00010000",5749 => "01111010",5750 => "00111110",5751 => "10101011",5752 => "00111001",5753 => "10000011",5754 => "01110110",5755 => "11000111",5756 => "00110100",5757 => "00011100",5758 => "11110110",5759 => "11000001",5760 => "00011100",5761 => "10110101",5762 => "00000010",5763 => "10110001",5764 => "01011011",5765 => "10011110",5766 => "10100111",5767 => "10100010",5768 => "00101110",5769 => "00101010",5770 => "10001110",5771 => "11010111",5772 => "10111011",5773 => "10100101",5774 => "01101101",5775 => "11101100",5776 => "11110011",5777 => "01110101",5778 => "11001000",5779 => "00010100",5780 => "11000011",5781 => "11011101",5782 => "11111011",5783 => "00011101",5784 => "00110011",5785 => "10101001",5786 => "11000001",5787 => "11101011",5788 => "01011101",5789 => "00110110",5790 => "10111000",5791 => "11101100",5792 => "00110010",5793 => "01001011",5794 => "10111100",5795 => "11110111",5796 => "10001001",5797 => "11001111",5798 => "11000000",5799 => "10001101",5800 => "01000010",5801 => "00101110",5802 => "11000111",5803 => "11011111",5804 => "00110000",5805 => "10011101",5806 => "11111100",5807 => "10101100",5808 => "10001010",5809 => "00000110",5810 => "00111001",5811 => "11110010",5812 => "11110101",5813 => "11010001",5814 => "11001111",5815 => "01010100",5816 => "00000101",5817 => "01011011",5818 => "00110100",5819 => "10101111",5820 => "10101110",5821 => "10111011",5822 => "10101011",5823 => "00000111",5824 => "00101011",5825 => "00100001",5826 => "11111001",5827 => "01001001",5828 => "11100101",5829 => "00011000",5830 => "00111110",5831 => "00110001",5832 => "10011000",5833 => "00110100",5834 => "01011111",5835 => "00110001",5836 => "01011111",5837 => "00101011",5838 => "00010001",5839 => "11010111",5840 => "00001011",5841 => "11101101",5842 => "11101011",5843 => "10011001",5844 => "11100101",5845 => "11101100",5846 => "11101100",5847 => "01001101",5848 => "10111110",5849 => "01011010",5850 => "10001110",5851 => "10100000",5852 => "01111110",5853 => "00110111",5854 => "01000111",5855 => "10110001",5856 => "10011011",5857 => "01100111",5858 => "11100001",5859 => "00000000",5860 => "10000011",5861 => "11010011",5862 => "10000001",5863 => "00101101",5864 => "01000101",5865 => "10101110",5866 => "01101100",5867 => "00110100",5868 => "11001000",5869 => "10010001",5870 => "11111011",5871 => "00100111",5872 => "00111010",5873 => "10111100",5874 => "11001001",5875 => "10100111",5876 => "00010101",5877 => "00100011",5878 => "10011010",5879 => "00100011",5880 => "00100110",5881 => "00001010",5882 => "11100001",5883 => "10110111",5884 => "00010110",5885 => "01111000",5886 => "11101011",5887 => "01000111",5888 => "00100010",5889 => "10011110",5890 => "00001101",5891 => "10110111",5892 => "11000000",5893 => "11000101",5894 => "11110100",5895 => "01011110",5896 => "01000101",5897 => "01111011",5898 => "00110001",5899 => "10110110",5900 => "10001111",5901 => "00100111",5902 => "01100000",5903 => "11111110",5904 => "10011010",5905 => "10011011",5906 => "10011100",5907 => "11010000",5908 => "10000000",5909 => "01100000",5910 => "00101111",5911 => "01110001",5912 => "00000010",5913 => "11010101",5914 => "11000001",5915 => "10101010",5916 => "00010010",5917 => "01001111",5918 => "10001001",5919 => "01011100",5920 => "11111000",5921 => "11001011",5922 => "11010100",5923 => "01001101",5924 => "11010111",5925 => "10001010",5926 => "11000001",5927 => "11101100",5928 => "00010000",5929 => "01010110",5930 => "00001011",5931 => "01011000",5932 => "01000101",5933 => "00000010",5934 => "00001010",5935 => "11110000",5936 => "00111010",5937 => "10110011",5938 => "10101001",5939 => "01011100",5940 => "01010100",5941 => "01111101",5942 => "00100011",5943 => "00101011",5944 => "11110100",5945 => "11111111",5946 => "00100001",5947 => "11010001",5948 => "00000001",5949 => "00111010",5950 => "01000110",5951 => "00111000",5952 => "10000110",5953 => "11000110",5954 => "01001110",5955 => "00101000",5956 => "01111001",5957 => "00011001",5958 => "01111000",5959 => "11100111",5960 => "01001011",5961 => "00000101",5962 => "00010010",5963 => "01101000",5964 => "00110001",5965 => "00001110",5966 => "00101010",5967 => "00100101",5968 => "00100110",5969 => "00011011",5970 => "11110101",5971 => "11000110",5972 => "01000000",5973 => "00011110",5974 => "00111110",5975 => "10010110",5976 => "00100101",5977 => "11010110",5978 => "11000000",5979 => "00011110",5980 => "01011011",5981 => "00101111",5982 => "10100111",5983 => "10001100",5984 => "10001100",5985 => "10110110",5986 => "01111100",5987 => "11011001",5988 => "01100111",5989 => "00001111",5990 => "10101000",5991 => "00011111",5992 => "00100011",5993 => "11010101",5994 => "00100000",5995 => "00001111",5996 => "10001010",5997 => "10101010",5998 => "00001100",5999 => "00101101",6000 => "00111110",6001 => "00011000",6002 => "11100001",6003 => "10101000",6004 => "11110010",6005 => "01010111",6006 => "01110001",6007 => "11110001",6008 => "00011110",6009 => "01110001",6010 => "11011101",6011 => "00111010",6012 => "01010111",6013 => "01100001",6014 => "10111001",6015 => "01011001",6016 => "11001000",6017 => "00010010",6018 => "00011001",6019 => "00001110",6020 => "10110110",6021 => "10000111",6022 => "01010001",6023 => "01010101",6024 => "10111011",6025 => "11101111",6026 => "11001111",6027 => "11111011",6028 => "00101010",6029 => "11000111",6030 => "10101101",6031 => "00101110",6032 => "00011010",6033 => "11101010",6034 => "00111110",6035 => "10101101",6036 => "00101100",6037 => "10010010",6038 => "10001011",6039 => "10011110",6040 => "01001010",6041 => "00010111",6042 => "11111100",6043 => "01001001",6044 => "00011000",6045 => "11001110",6046 => "11001010",6047 => "11000100",6048 => "01000011",6049 => "11101001",6050 => "01001010",6051 => "11000110",6052 => "01111111",6053 => "10100100",6054 => "10011111",6055 => "11010001",6056 => "01011101",6057 => "10011000",6058 => "00010110",6059 => "10101010",6060 => "10101011",6061 => "01111110",6062 => "10011111",6063 => "01000000",6064 => "01111010",6065 => "00100111",6066 => "01001001",6067 => "00110000",6068 => "11010110",6069 => "01001000",6070 => "00101001",6071 => "00010111",6072 => "10111011",6073 => "00011110",6074 => "11100000",6075 => "11000100",6076 => "00001110",6077 => "00000001",6078 => "10101100",6079 => "10000101",6080 => "00100111",6081 => "10101001",6082 => "11101100",6083 => "01111111",6084 => "00000010",6085 => "11010000",6086 => "01111001",6087 => "11100010",6088 => "10000011",6089 => "01000010",6090 => "00110111",6091 => "10010110",6092 => "11000101",6093 => "10110101",6094 => "10000000",6095 => "11100101",6096 => "10101010",6097 => "01101000",6098 => "01000110",6099 => "10111011",6100 => "10001011",6101 => "01010000",6102 => "11100001",6103 => "10100101",6104 => "00010111",6105 => "11111111",6106 => "11000000",6107 => "11001101",6108 => "11100100",6109 => "11001001",6110 => "10011111",6111 => "01101000",6112 => "00111110",6113 => "01101100",6114 => "01100111",6115 => "10111000",6116 => "11010010",6117 => "00100000",6118 => "10111000",6119 => "00101100",6120 => "11010101",6121 => "11111001",6122 => "01000101",6123 => "10100011",6124 => "00110011",6125 => "01011000",6126 => "01110100",6127 => "00010110",6128 => "00011100",6129 => "11101001",6130 => "10001011",6131 => "10100000",6132 => "01100101",6133 => "01110110",6134 => "10100001",6135 => "00000001",6136 => "11100111",6137 => "01101100",6138 => "00110010",6139 => "11111101",6140 => "10010101",6141 => "10000111",6142 => "00001010",6143 => "11111110",6144 => "01110101",6145 => "11000010",6146 => "11111000",6147 => "00000101",6148 => "10100001",6149 => "10011110",6150 => "10011001",6151 => "00010011",6152 => "01100010",6153 => "10111110",6154 => "01010101",6155 => "10111100",6156 => "11100000",6157 => "10000001",6158 => "00000010",6159 => "00001101",6160 => "00100011",6161 => "11010010",6162 => "11101000",6163 => "11110100",6164 => "00001101",6165 => "10001100",6166 => "10011011",6167 => "00011000",6168 => "01100110",6169 => "00011101",6170 => "00100111",6171 => "00010111",6172 => "10110011",6173 => "11011001",6174 => "00111110",6175 => "10010111",6176 => "11111101",6177 => "11010010",6178 => "00111110",6179 => "01000110",6180 => "11101111",6181 => "01110000",6182 => "11011111",6183 => "11011111",6184 => "11000101",6185 => "10100111",6186 => "01000110",6187 => "11100011",6188 => "00011001",6189 => "01000101",6190 => "11011110",6191 => "10101100",6192 => "11000100",6193 => "11111010",6194 => "10110100",6195 => "10000011",6196 => "11110001",6197 => "11111010",6198 => "00100100",6199 => "11110111",6200 => "10001110",6201 => "01001011",6202 => "00000000",6203 => "10000000",6204 => "11001001",6205 => "11111011",6206 => "01110011",6207 => "00100000",6208 => "00111110",6209 => "10001011",6210 => "10001001",6211 => "00011011",6212 => "10011001",6213 => "00011011",6214 => "01111100",6215 => "11101010",6216 => "01110110",6217 => "10000100",6218 => "10001110",6219 => "00010110",6220 => "11010001",6221 => "00100101",6222 => "00111101",6223 => "11110111",6224 => "00011011",6225 => "00101001",6226 => "11001100",6227 => "11001011",6228 => "01001110",6229 => "00111110",6230 => "00111010",6231 => "10101011",6232 => "10010111",6233 => "00100100",6234 => "11110101",6235 => "11100110",6236 => "11001100",6237 => "10001001",6238 => "11110110",6239 => "10111100",6240 => "11001001",6241 => "01101011",6242 => "11100101",6243 => "01111000",6244 => "00101101",6245 => "10110101",6246 => "00100010",6247 => "10010101",6248 => "11001111",6249 => "00010011",6250 => "11000111",6251 => "10111010",6252 => "01000000",6253 => "11011101",6254 => "10010100",6255 => "11001011",6256 => "11110000",6257 => "00111000",6258 => "10101010",6259 => "11010101",6260 => "01101010",6261 => "00011010",6262 => "00100000",6263 => "10111000",6264 => "11001101",6265 => "00101000",6266 => "11100101",6267 => "01011101",6268 => "10101111",6269 => "01110111",6270 => "01110000",6271 => "00110001",6272 => "00111000",6273 => "00011111",6274 => "01000010",6275 => "00111100",6276 => "00000100",6277 => "10101000",6278 => "01000010",6279 => "10101110",6280 => "01010011",6281 => "00011100",6282 => "10101000",6283 => "00000000",6284 => "00011101",6285 => "11001011",6286 => "11010100",6287 => "01001011",6288 => "01010111",6289 => "01101011",6290 => "00100011",6291 => "01101011",6292 => "11100011",6293 => "10110011",6294 => "10100111",6295 => "11000011",6296 => "00011110",6297 => "01100101",6298 => "11000000",6299 => "00011000",6300 => "10100001",6301 => "00110100",6302 => "00101011",6303 => "11110111",6304 => "01111011",6305 => "11111010",6306 => "10110110",6307 => "01110111",6308 => "00110111",6309 => "01000111",6310 => "10111101",6311 => "00000011",6312 => "00011110",6313 => "10010101",6314 => "10111011",6315 => "00101011",6316 => "00100100",6317 => "00110101",6318 => "00110100",6319 => "00101011",6320 => "10111111",6321 => "11001101",6322 => "01001111",6323 => "01010110",6324 => "10110010",6325 => "00001010",6326 => "11010100",6327 => "10001011",6328 => "01110011",6329 => "10000101",6330 => "10110000",6331 => "10011001",6332 => "11000011",6333 => "00100011",6334 => "10010010",6335 => "10011010",6336 => "01101001",6337 => "00011001",6338 => "11111101",6339 => "10000000",6340 => "00110111",6341 => "00010110",6342 => "01010111",6343 => "10111010",6344 => "11000001",6345 => "00000100",6346 => "01111000",6347 => "11010110",6348 => "01110110",6349 => "11101000",6350 => "00000100",6351 => "01101111",6352 => "11010010",6353 => "00111101",6354 => "00011110",6355 => "11000011",6356 => "01101010",6357 => "11101101",6358 => "10001100",6359 => "01100001",6360 => "01110000",6361 => "10001011",6362 => "00011010",6363 => "10110110",6364 => "01110001",6365 => "01011001",6366 => "11100111",6367 => "00101110",6368 => "00011101",6369 => "11000110",6370 => "11111010",6371 => "10011000",6372 => "01000011",6373 => "11000011",6374 => "10011011",6375 => "00010001",6376 => "10011000",6377 => "01110101",6378 => "11110111",6379 => "00100110",6380 => "10100101",6381 => "00101110",6382 => "11001000",6383 => "10010101",6384 => "10011001",6385 => "10111110",6386 => "01000110",6387 => "10000110",6388 => "11101100",6389 => "11010001",6390 => "01000100",6391 => "00110010",6392 => "11011101",6393 => "11101000",6394 => "01001101",6395 => "00111101",6396 => "01010101",6397 => "01110101",6398 => "00110110",6399 => "11100111",6400 => "10000101",6401 => "11011111",6402 => "00111101",6403 => "11101011",6404 => "10010101",6405 => "11100100",6406 => "01011010",6407 => "00110100",6408 => "11110101",6409 => "00000001",6410 => "00001111",6411 => "01100111",6412 => "10101000",6413 => "00110110",6414 => "01111101",6415 => "11001101",6416 => "10000110",6417 => "00110111",6418 => "01010011",6419 => "11111101",6420 => "01010100",6421 => "11010011",6422 => "10001110",6423 => "01011001",6424 => "01011000",6425 => "00111001",6426 => "11001000",6427 => "01001000",6428 => "11000110",6429 => "00110101",6430 => "01010000",6431 => "10011100",6432 => "10010101",6433 => "00011110",6434 => "01001110",6435 => "11110110",6436 => "10100010",6437 => "11011110",6438 => "01001111",6439 => "11100100",6440 => "00010001",6441 => "00111001",6442 => "01000011",6443 => "00100111",6444 => "00010100",6445 => "11110100",6446 => "00111111",6447 => "00011011",6448 => "01010100",6449 => "01110110",6450 => "11001011",6451 => "01100100",6452 => "11101001",6453 => "10000111",6454 => "01110110",6455 => "01111110",6456 => "01010001",6457 => "00000001",6458 => "10111100",6459 => "01110011",6460 => "10110011",6461 => "00100010",6462 => "01110110",6463 => "11111010",6464 => "01101111",6465 => "01000100",6466 => "10110101",6467 => "10000110",6468 => "10110001",6469 => "11000000",6470 => "01001111",6471 => "01100100",6472 => "01101100",6473 => "11101110",6474 => "10010101",6475 => "01110101",6476 => "10101001",6477 => "00000010",6478 => "00100111",6479 => "10111000",6480 => "11110000",6481 => "11111001",6482 => "11000011",6483 => "00100001",6484 => "10110110",6485 => "11111011",6486 => "10111111",6487 => "10010101",6488 => "00001100",6489 => "00001010",6490 => "01111011",6491 => "01111111",6492 => "00011001",6493 => "00110100",6494 => "00111100",6495 => "00011000",6496 => "10110011",6497 => "01101000",6498 => "01011001",6499 => "00001001",6500 => "00001100",6501 => "11010101",6502 => "11100010",6503 => "00110010",6504 => "01000010",6505 => "01111010",6506 => "10001100",6507 => "10111000",6508 => "00111011",6509 => "00010010",6510 => "11000000",6511 => "00101000",6512 => "00001001",6513 => "11001001",6514 => "00111011",6515 => "00100000",6516 => "00101001",6517 => "00001011",6518 => "10101010",6519 => "00000000",6520 => "00011101",6521 => "00110101",6522 => "00101011",6523 => "10101011",6524 => "11110001",6525 => "10100001",6526 => "11010111",6527 => "00000010",6528 => "00010010",6529 => "01010101",6530 => "11011110",6531 => "01101110",6532 => "10000110",6533 => "10010010",6534 => "01111100",6535 => "01001101",6536 => "00000001",6537 => "00101101",6538 => "01111101",6539 => "01111111",6540 => "00000101",6541 => "00010000",6542 => "01101000",6543 => "10100110",6544 => "01001001",6545 => "01111000",6546 => "01011100",6547 => "00111010",6548 => "11101000",6549 => "10110101",6550 => "11110001",6551 => "00000101",6552 => "01101110",6553 => "11110110",6554 => "01110001",6555 => "01101011",6556 => "10011111",6557 => "01101111",6558 => "10000101",6559 => "00100011",6560 => "11001110",6561 => "01001011",6562 => "01101110",6563 => "01111000",6564 => "11010101",6565 => "00101000",6566 => "11000101",6567 => "00110010",6568 => "01010101",6569 => "11100000",6570 => "10001010",6571 => "10110001",6572 => "10010101",6573 => "00011010",6574 => "01111001",6575 => "11100110",6576 => "11011000",6577 => "11110101",6578 => "10001100",6579 => "01010010",6580 => "00110101",6581 => "01111111",6582 => "01100010",6583 => "11110001",6584 => "00110010",6585 => "00001101",6586 => "10011011",6587 => "10110010",6588 => "00000111",6589 => "10010101",6590 => "01001101",6591 => "10000010",6592 => "01000000",6593 => "01100100",6594 => "11101110",6595 => "10010010",6596 => "11001000",6597 => "01101111",6598 => "10011000",6599 => "01111000",6600 => "01110110",6601 => "11010011",6602 => "10011010",6603 => "11010001",6604 => "00010011",6605 => "00110011",6606 => "00001001",6607 => "11100011",6608 => "01100111",6609 => "11110110",6610 => "10001011",6611 => "10011010",6612 => "01000011",6613 => "10111111",6614 => "01000110",6615 => "11111110",6616 => "11111100",6617 => "11011100",6618 => "11111000",6619 => "10111100",6620 => "01110000",6621 => "11000001",6622 => "01110100",6623 => "00010000",6624 => "00110100",6625 => "01000110",6626 => "00101001",6627 => "11000111",6628 => "11101011",6629 => "01010100",6630 => "01000000",6631 => "01111111",6632 => "10111000",6633 => "10001110",6634 => "00100111",6635 => "10010110",6636 => "00100111",6637 => "00000100",6638 => "01001101",6639 => "10110100",6640 => "10010101",6641 => "10101001",6642 => "00011001",6643 => "01111001",6644 => "00010011",6645 => "00001000",6646 => "11011101",6647 => "10111111",6648 => "11101010",6649 => "10110000",6650 => "00111000",6651 => "00111101",6652 => "11110110",6653 => "00100101",6654 => "11111011",6655 => "00101100",6656 => "00111010",6657 => "00111101",6658 => "00011111",6659 => "11110010",6660 => "11010001",6661 => "11010110",6662 => "11101100",6663 => "11010100",6664 => "10110101",6665 => "01011011",6666 => "00100111",6667 => "01100001",6668 => "00110111",6669 => "01001111",6670 => "11111000",6671 => "01100001",6672 => "01100011",6673 => "10110100",6674 => "00011010",6675 => "01110111",6676 => "11111101",6677 => "11100010",6678 => "01101010",6679 => "10100101",6680 => "11100010",6681 => "10110101",6682 => "10101010",6683 => "11000110",6684 => "00011011",6685 => "10011110",6686 => "10110101",6687 => "11000001",6688 => "11000101",6689 => "01011110",6690 => "10100111",6691 => "11010110",6692 => "11000101",6693 => "00010100",6694 => "01010100",6695 => "00010110",6696 => "01111000",6697 => "00101111",6698 => "10011100",6699 => "11010011",6700 => "10101010",6701 => "00111001",6702 => "01001101",6703 => "01101110",6704 => "11000101",6705 => "10011010",6706 => "00111110",6707 => "01010110",6708 => "10110001",6709 => "00101100",6710 => "11111101",6711 => "00110100",6712 => "10001001",6713 => "01011111",6714 => "11110101",6715 => "01101111",6716 => "00010011",6717 => "00000000",6718 => "10000101",6719 => "01100001",6720 => "00111000",6721 => "00110010",6722 => "00111111",6723 => "11001100",6724 => "11011101",6725 => "00001000",6726 => "11110000",6727 => "01000100",6728 => "11101010",6729 => "10010011",6730 => "10010100",6731 => "01101001",6732 => "01000000",6733 => "01111010",6734 => "10101001",6735 => "01001110",6736 => "00111001",6737 => "10110100",6738 => "11010011",6739 => "11100100",6740 => "11101100",6741 => "10110111",6742 => "00001101",6743 => "11111000",6744 => "00100111",6745 => "11110011",6746 => "10001110",6747 => "00001010",6748 => "11110101",6749 => "11111010",6750 => "10110111",6751 => "11100100",6752 => "11101000",6753 => "01001001",6754 => "10101010",6755 => "11000001",6756 => "00110111",6757 => "01001101",6758 => "11000010",6759 => "10000100",6760 => "01000101",6761 => "01111010",6762 => "10100001",6763 => "10111110",6764 => "00111001",6765 => "00111001",6766 => "01100111",6767 => "11111000",6768 => "10110101",6769 => "11011011",6770 => "00010000",6771 => "11001101",6772 => "11110101",6773 => "00111101",6774 => "11001101",6775 => "01101011",6776 => "10100110",6777 => "01000101",6778 => "11011010",6779 => "11111010",6780 => "01111101",6781 => "10000110",6782 => "11100101",6783 => "10100110",6784 => "00100101",6785 => "11000010",6786 => "11011001",6787 => "00000101",6788 => "01110101",6789 => "11000111",6790 => "01111101",6791 => "10100110",6792 => "10011100",6793 => "01110011",6794 => "11101101",6795 => "10000111",6796 => "10110000",6797 => "00001101",6798 => "00010010",6799 => "11000111",6800 => "00011101",6801 => "01111000",6802 => "10010001",6803 => "00101101",6804 => "11001001",6805 => "11000001",6806 => "01100101",6807 => "00101111",6808 => "00100100",6809 => "00010101",6810 => "10001101",6811 => "10010010",6812 => "01110010",6813 => "10111100",6814 => "01000001",6815 => "10001001",6816 => "01000011",6817 => "11101111",6818 => "01100001",6819 => "01111000",6820 => "11000000",6821 => "11111001",6822 => "10001111",6823 => "10011000",6824 => "01011101",6825 => "01011000",6826 => "11110111",6827 => "10101000",6828 => "11111100",6829 => "01001110",6830 => "00101110",6831 => "00010101",6832 => "10000111",6833 => "11101011",6834 => "11111101",6835 => "00001110",6836 => "10011111",6837 => "10000111",6838 => "00000111",6839 => "01001100",6840 => "01101000",6841 => "00110000",6842 => "11111001",6843 => "10001111",6844 => "10100100",6845 => "10010011",6846 => "00010001",6847 => "01010111",6848 => "00100000",6849 => "00111110",6850 => "11010111",6851 => "11010011",6852 => "10101000",6853 => "01101011",6854 => "11011111",6855 => "10010001",6856 => "10011110",6857 => "00100111",6858 => "11010100",6859 => "01100100",6860 => "00000011",6861 => "10110100",6862 => "10010000",6863 => "01011111",6864 => "10100011",6865 => "10001001",6866 => "10110011",6867 => "10011010",6868 => "11100010",6869 => "10110100",6870 => "00001010",6871 => "11010111",6872 => "00010101",6873 => "10011110",6874 => "11011100",6875 => "00010000",6876 => "11110010",6877 => "00101001",6878 => "10000101",6879 => "00000101",6880 => "00111001",6881 => "11001010",6882 => "00011001",6883 => "11101110",6884 => "01001100",6885 => "01111000",6886 => "11100100",6887 => "01001100",6888 => "10000100",6889 => "10110111",6890 => "00011010",6891 => "11110100",6892 => "10010001",6893 => "01011111",6894 => "01000111",6895 => "00010011",6896 => "11111010",6897 => "00101100",6898 => "01100010",6899 => "10010000",6900 => "01000110",6901 => "11001011",6902 => "00111000",6903 => "00000110",6904 => "11100101",6905 => "00001010",6906 => "11110110",6907 => "01000011",6908 => "01101000",6909 => "10111001",6910 => "11010000",6911 => "01011000",6912 => "00010101",6913 => "10001100",6914 => "01101011",6915 => "00110111",6916 => "01100101",6917 => "11000010",6918 => "10010011",6919 => "01111011",6920 => "10001000",6921 => "11101101",6922 => "10101011",6923 => "10100101",6924 => "11010001",6925 => "00001001",6926 => "11001011",6927 => "01111111",6928 => "11010010",6929 => "00110101",6930 => "00010010",6931 => "10101110",6932 => "11001110",6933 => "10111010",6934 => "00110001",6935 => "11010101",6936 => "11000010",6937 => "01100101",6938 => "01111111",6939 => "00001001",6940 => "01110010",6941 => "00101111",6942 => "00110000",6943 => "11001001",6944 => "10001110",6945 => "00010000",6946 => "10111100",6947 => "00100000",6948 => "10110101",6949 => "10100011",6950 => "00111011",6951 => "01101110",6952 => "01001000",6953 => "01100110",6954 => "10011010",6955 => "10010010",6956 => "11001111",6957 => "10110001",6958 => "11001100",6959 => "01100101",6960 => "01010010",6961 => "10111101",6962 => "10100010",6963 => "01110010",6964 => "10110110",6965 => "00111001",6966 => "01010011",6967 => "00001111",6968 => "10000001",6969 => "10010010",6970 => "01111101",6971 => "10010101",6972 => "10111101",6973 => "00111111",6974 => "00001000",6975 => "01001110",6976 => "00011100",6977 => "00101100",6978 => "01100001",6979 => "10100111",6980 => "00111110",6981 => "01001000",6982 => "01110000",6983 => "11101000",6984 => "10011001",6985 => "00111011",6986 => "01110110",6987 => "01100001",6988 => "01001011",6989 => "00011001",6990 => "01101101",6991 => "11111111",6992 => "01001111",6993 => "10001001",6994 => "11100011",6995 => "00001100",6996 => "11101000",6997 => "00100011",6998 => "00101100",6999 => "11100011",7000 => "01111101",7001 => "10011100",7002 => "10001000",7003 => "01011100",7004 => "11010110",7005 => "11001111",7006 => "10001011",7007 => "01001010",7008 => "01001001",7009 => "00101000",7010 => "11111000",7011 => "11110110",7012 => "11000010",7013 => "11100000",7014 => "01100001",7015 => "00111001",7016 => "00010000",7017 => "01000011",7018 => "10000000",7019 => "00000010",7020 => "01111110",7021 => "10001000",7022 => "01101001",7023 => "11101110",7024 => "11111111",7025 => "00100011",7026 => "01001110",7027 => "01101011",7028 => "00000111",7029 => "10001000",7030 => "10101110",7031 => "10010101",7032 => "11110111",7033 => "00001111",7034 => "00100001",7035 => "00110110",7036 => "00000011",7037 => "00000101",7038 => "10010011",7039 => "10001010",7040 => "00100001",7041 => "11110111",7042 => "11001000",7043 => "01001101",7044 => "01000000",7045 => "10011010",7046 => "00100111",7047 => "00101011",7048 => "01001010",7049 => "01101100",7050 => "01001111",7051 => "01000101",7052 => "00111101",7053 => "01100010",7054 => "01010100",7055 => "00110001",7056 => "10111000",7057 => "00011000",7058 => "01111010",7059 => "00000001",7060 => "10001011",7061 => "01110110",7062 => "01001000",7063 => "11100010",7064 => "11000101",7065 => "01000110",7066 => "10010010",7067 => "10001001",7068 => "01011110",7069 => "01101010",7070 => "10010110",7071 => "00101101",7072 => "00101000",7073 => "10001011",7074 => "10101100",7075 => "01110011",7076 => "10101111",7077 => "00001111",7078 => "01000111",7079 => "00011000",7080 => "11100111",7081 => "01110011",7082 => "00011001",7083 => "00010010",7084 => "10001001",7085 => "10111101",7086 => "11101101",7087 => "11001111",7088 => "00001111",7089 => "10010101",7090 => "00011000",7091 => "00010010",7092 => "01010011",7093 => "10010011",7094 => "11010010",7095 => "11100110",7096 => "10011100",7097 => "11010011",7098 => "01001011",7099 => "00110010",7100 => "10110101",7101 => "01110010",7102 => "01100001",7103 => "00110001",7104 => "11101111",7105 => "11000101",7106 => "10011111",7107 => "00000011",7108 => "01110000",7109 => "11000110",7110 => "01100110",7111 => "11100001",7112 => "10010100",7113 => "00101011",7114 => "01101000",7115 => "11111111",7116 => "00000100",7117 => "11000110",7118 => "11011000",7119 => "00010101",7120 => "10111010",7121 => "00100111",7122 => "01011000",7123 => "01110110",7124 => "01110100",7125 => "01111111",7126 => "01100000",7127 => "10111001",7128 => "11100101",7129 => "10001011",7130 => "00101111",7131 => "00110010",7132 => "00101011",7133 => "10101011",7134 => "10110001",7135 => "01011001",7136 => "00010110",7137 => "01110011",7138 => "10111001",7139 => "10001101",7140 => "10100000",7141 => "10010001",7142 => "10010001",7143 => "11010011",7144 => "10111010",7145 => "01011011",7146 => "10101101",7147 => "11101001",7148 => "10101110",7149 => "00101100",7150 => "00000000",7151 => "11010101",7152 => "10110011",7153 => "01111110",7154 => "11010101",7155 => "10100011",7156 => "10001001",7157 => "00100100",7158 => "10111000",7159 => "00000010",7160 => "10010010",7161 => "00001001",7162 => "10011011",7163 => "10010010",7164 => "10100001",7165 => "10010101",7166 => "10010011",7167 => "11111001",7168 => "00110000",7169 => "00010011",7170 => "10101101",7171 => "11000110",7172 => "10101000",7173 => "10110000",7174 => "00110010",7175 => "10101000",7176 => "01010010",7177 => "10110000",7178 => "01011101",7179 => "00001001",7180 => "00100011",7181 => "11101111",7182 => "11001000",7183 => "01011111",7184 => "11011100",7185 => "10010000",7186 => "00001101",7187 => "00000100",7188 => "11011001",7189 => "01001000",7190 => "10101111",7191 => "10101110",7192 => "11011111",7193 => "10010101",7194 => "10000110",7195 => "00011111",7196 => "11110000",7197 => "10100100",7198 => "00000111",7199 => "01100100",7200 => "10101001",7201 => "10010001",7202 => "10101011",7203 => "00110110",7204 => "11110111",7205 => "00011110",7206 => "10000011",7207 => "01000111",7208 => "10001110",7209 => "11000000",7210 => "10111010",7211 => "11111101",7212 => "01010000",7213 => "01011101",7214 => "11100011",7215 => "11111010",7216 => "00011111",7217 => "01010000",7218 => "10110010",7219 => "11000101",7220 => "11011101",7221 => "01110010",7222 => "00001001",7223 => "10100101",7224 => "11011010",7225 => "00100101",7226 => "11001101",7227 => "10011001",7228 => "01100001",7229 => "10000100",7230 => "01001110",7231 => "00110010",7232 => "10111100",7233 => "10011101",7234 => "00101101",7235 => "00000000",7236 => "00001001",7237 => "10001101",7238 => "10001100",7239 => "01011101",7240 => "11111110",7241 => "10010111",7242 => "01110011",7243 => "10011001",7244 => "10101010",7245 => "10100110",7246 => "01010111",7247 => "10000011",7248 => "10011111",7249 => "01100011",7250 => "01010010",7251 => "01010110",7252 => "01001111",7253 => "10001111",7254 => "11111100",7255 => "11110100",7256 => "00111101",7257 => "10000011",7258 => "11000101",7259 => "00110111",7260 => "01100101",7261 => "10000111",7262 => "11010110",7263 => "01001011",7264 => "11000001",7265 => "01000001",7266 => "10110010",7267 => "10110101",7268 => "00101101",7269 => "00001101",7270 => "11100001",7271 => "10110111",7272 => "00011010",7273 => "10101110",7274 => "10011100",7275 => "01001011",7276 => "00000001",7277 => "00010110",7278 => "01011111",7279 => "00110000",7280 => "01110111",7281 => "10100001",7282 => "01111000",7283 => "01100001",7284 => "10111101",7285 => "00100111",7286 => "10101010",7287 => "01001101",7288 => "11100110",7289 => "00101111",7290 => "10000011",7291 => "10010111",7292 => "11111111",7293 => "11101011",7294 => "10110111",7295 => "11100101",7296 => "11111011",7297 => "01011001",7298 => "01110101",7299 => "00000000",7300 => "10111011",7301 => "00011000",7302 => "10100001",7303 => "11101111",7304 => "10110011",7305 => "00111111",7306 => "11111101",7307 => "10010110",7308 => "11111101",7309 => "10101100",7310 => "01010011",7311 => "01111110",7312 => "01111000",7313 => "10110101",7314 => "11000110",7315 => "10100111",7316 => "11011011",7317 => "11010100",7318 => "00001110",7319 => "01010001",7320 => "10010011",7321 => "01000001",7322 => "00001101",7323 => "01011101",7324 => "00010101",7325 => "00100011",7326 => "10110111",7327 => "10110010",7328 => "00101110",7329 => "00110111",7330 => "01110010",7331 => "10101011",7332 => "10000101",7333 => "11101001",7334 => "01000000",7335 => "00001101",7336 => "01011100",7337 => "00001110",7338 => "10011010",7339 => "00011010",7340 => "00111101",7341 => "10010001",7342 => "00110100",7343 => "01001000",7344 => "11001011",7345 => "10010101",7346 => "00011011",7347 => "00100001",7348 => "00100100",7349 => "01001001",7350 => "01110111",7351 => "11010000",7352 => "01011111",7353 => "11101001",7354 => "00001100",7355 => "01001100",7356 => "11011100",7357 => "01001100",7358 => "11000010",7359 => "00000000",7360 => "11011101",7361 => "01011011",7362 => "01000010",7363 => "01011001",7364 => "01111100",7365 => "01010010",7366 => "11111101",7367 => "01001110",7368 => "01110101",7369 => "01111100",7370 => "11100101",7371 => "10111011",7372 => "00100101",7373 => "11001010",7374 => "00010111",7375 => "11001110",7376 => "11101111",7377 => "11110001",7378 => "11000001",7379 => "10000011",7380 => "00110100",7381 => "10111110",7382 => "10101010",7383 => "00010111",7384 => "01011111",7385 => "01110110",7386 => "11100101",7387 => "00111100",7388 => "11010111",7389 => "01110000",7390 => "01001010",7391 => "10001100",7392 => "00000011",7393 => "10100111",7394 => "01001100",7395 => "10111000",7396 => "10101010",7397 => "10101101",7398 => "11110111",7399 => "10000100",7400 => "01000000",7401 => "01101101",7402 => "11011100",7403 => "10100111",7404 => "11001011",7405 => "11010010",7406 => "11000100",7407 => "11000100",7408 => "01000010",7409 => "00010111",7410 => "01111110",7411 => "10010011",7412 => "10110111",7413 => "01111000",7414 => "10111001",7415 => "10000011",7416 => "10101001",7417 => "10010101",7418 => "01000100",7419 => "11100010",7420 => "01110010",7421 => "00011010",7422 => "00110100",7423 => "01010001",7424 => "00101101",7425 => "01101111",7426 => "00001110",7427 => "01011001",7428 => "00110111",7429 => "01000110",7430 => "01010110",7431 => "10100100",7432 => "00000110",7433 => "10000011",7434 => "10011011",7435 => "01111000",7436 => "01101101",7437 => "00011011",7438 => "11001001",7439 => "10001110",7440 => "11101000",7441 => "00000110",7442 => "10010001",7443 => "10111000",7444 => "10111010",7445 => "01011111",7446 => "01001011",7447 => "00001111",7448 => "01001111",7449 => "00000010",7450 => "11011111",7451 => "01101010",7452 => "11010010",7453 => "10100110",7454 => "00101011",7455 => "00100001",7456 => "01101100",7457 => "01100010",7458 => "00101111",7459 => "01000001",7460 => "10000001",7461 => "00011111",7462 => "10110001",7463 => "11010001",7464 => "00000111",7465 => "00011110",7466 => "00101011",7467 => "11110110",7468 => "10101101",7469 => "10001000",7470 => "00101110",7471 => "01110110",7472 => "00010110",7473 => "11100111",7474 => "11010001",7475 => "11011100",7476 => "11001110",7477 => "11110110",7478 => "11101110",7479 => "10011000",7480 => "10001100",7481 => "01110110",7482 => "01001100",7483 => "00101111",7484 => "00101101",7485 => "11110011",7486 => "10001011",7487 => "01110010",7488 => "00011101",7489 => "10000011",7490 => "01111100",7491 => "10110000",7492 => "00100010",7493 => "00100010",7494 => "00011000",7495 => "10111001",7496 => "00110010",7497 => "11111101",7498 => "11101101",7499 => "01100000",7500 => "01011011",7501 => "01110110",7502 => "10110111",7503 => "10000011",7504 => "11101000",7505 => "11110101",7506 => "00011010",7507 => "01001111",7508 => "01101110",7509 => "10010111",7510 => "10000110",7511 => "01101000",7512 => "10001010",7513 => "10110110",7514 => "10100110",7515 => "01100001",7516 => "11100101",7517 => "00011000",7518 => "00110011",7519 => "11001010",7520 => "01010010",7521 => "00011100",7522 => "00101110",7523 => "11001011",7524 => "10101010",7525 => "01010100",7526 => "10100101",7527 => "10100110",7528 => "00001100",7529 => "01011000",7530 => "00010101",7531 => "10100111",7532 => "00110011",7533 => "11101011",7534 => "10111101",7535 => "00101001",7536 => "11011001",7537 => "11011010",7538 => "01100000",7539 => "10100101",7540 => "00011011",7541 => "11110110",7542 => "01010000",7543 => "10000111",7544 => "01011101",7545 => "11011001",7546 => "01001011",7547 => "01110111",7548 => "01010010",7549 => "11010001",7550 => "10101101",7551 => "10011010",7552 => "11000111",7553 => "10100010",7554 => "01111101",7555 => "11100111",7556 => "00001010",7557 => "01011011",7558 => "00110101",7559 => "11011011",7560 => "01110101",7561 => "10111111",7562 => "01111010",7563 => "01000010",7564 => "01101011",7565 => "10100001",7566 => "01011001",7567 => "00101011",7568 => "01110001",7569 => "10100100",7570 => "11000111",7571 => "00110101",7572 => "10110111",7573 => "10011000",7574 => "01011010",7575 => "00011001",7576 => "01011100",7577 => "11010011",7578 => "11010001",7579 => "10100100",7580 => "01101010",7581 => "10010001",7582 => "10001111",7583 => "11111010",7584 => "01010111",7585 => "01001101",7586 => "11110010",7587 => "11011101",7588 => "11111010",7589 => "10001100",7590 => "10100010",7591 => "01111111",7592 => "11100110",7593 => "01010000",7594 => "10110000",7595 => "00101000",7596 => "01001000",7597 => "01001010",7598 => "10001101",7599 => "11100101",7600 => "01010100",7601 => "10001001",7602 => "11001100",7603 => "10110101",7604 => "01010001",7605 => "01001111",7606 => "00100101",7607 => "01100111",7608 => "11100000",7609 => "01111111",7610 => "00110111",7611 => "10101111",7612 => "01111111",7613 => "00011001",7614 => "11100011",7615 => "10001000",7616 => "11111001",7617 => "10110010",7618 => "11010011",7619 => "11001000",7620 => "10111111",7621 => "11001101",7622 => "10001001",7623 => "10101000",7624 => "00110010",7625 => "01011110",7626 => "00010010",7627 => "11001000",7628 => "01101011",7629 => "00100110",7630 => "10011010",7631 => "01110011",7632 => "00001010",7633 => "01010111",7634 => "10001100",7635 => "11100110",7636 => "10100110",7637 => "10110110",7638 => "10111011",7639 => "00001110",7640 => "11101011",7641 => "11011010",7642 => "11010011",7643 => "11011000",7644 => "00111010",7645 => "00000100",7646 => "11001110",7647 => "00001000",7648 => "11111101",7649 => "00110001",7650 => "11000011",7651 => "11001000",7652 => "01111101",7653 => "10001101",7654 => "10101001",7655 => "10100110",7656 => "11000100",7657 => "01110000",7658 => "01111110",7659 => "10100100",7660 => "01011110",7661 => "01100001",7662 => "10011011",7663 => "00100000",7664 => "01100111",7665 => "10010011",7666 => "11101010",7667 => "01110001",7668 => "01010010",7669 => "01111110",7670 => "11111110",7671 => "00101011",7672 => "01110111",7673 => "11001111",7674 => "01000110",7675 => "00111101",7676 => "00000011",7677 => "00101001",7678 => "10011100",7679 => "01001110",7680 => "11010001",7681 => "10100100",7682 => "10000000",7683 => "11000010",7684 => "11101111",7685 => "01111011",7686 => "11111100",7687 => "10000011",7688 => "11110001",7689 => "11010010",7690 => "11111000",7691 => "10000010",7692 => "01101010",7693 => "11111010",7694 => "01000001",7695 => "00110110",7696 => "11000100",7697 => "01110111",7698 => "01100010",7699 => "01000010",7700 => "10000000",7701 => "01111101",7702 => "11111100",7703 => "01011011",7704 => "11001110",7705 => "10011010",7706 => "00011100",7707 => "11011111",7708 => "10000010",7709 => "00101100",7710 => "11110001",7711 => "00100111",7712 => "11100010",7713 => "00100111",7714 => "10000110",7715 => "01100110",7716 => "11111000",7717 => "11011100",7718 => "10010001",7719 => "01010100",7720 => "10100101",7721 => "00011100",7722 => "00100001",7723 => "00111010",7724 => "11001111",7725 => "01000001",7726 => "11101111",7727 => "00011000",7728 => "01101010",7729 => "11101011",7730 => "10001111",7731 => "10011001",7732 => "10010001",7733 => "01101001",7734 => "11100101",7735 => "00011101",7736 => "10010110",7737 => "11111101",7738 => "01100100",7739 => "00000101",7740 => "11001100",7741 => "00111101",7742 => "11001001",7743 => "00000111",7744 => "01001001",7745 => "01110001",7746 => "01111000",7747 => "10110011",7748 => "00010000",7749 => "00000110",7750 => "11010100",7751 => "11010011",7752 => "11111010",7753 => "10011011",7754 => "10111010",7755 => "10110010",7756 => "01000011",7757 => "01010110",7758 => "11100010",7759 => "11100100",7760 => "10000001",7761 => "01111001",7762 => "01101010",7763 => "01001010",7764 => "01010100",7765 => "10111110",7766 => "00101110",7767 => "10000001",7768 => "01101100",7769 => "01110100",7770 => "11100101",7771 => "10111100",7772 => "10010010",7773 => "01000101",7774 => "01101100",7775 => "01100101",7776 => "00111001",7777 => "11001011",7778 => "00110011",7779 => "00110110",7780 => "10100101",7781 => "10001010",7782 => "10110101",7783 => "00010100",7784 => "10000100",7785 => "11100111",7786 => "00100111",7787 => "01010101",7788 => "01000100",7789 => "00100101",7790 => "00011100",7791 => "11111100",7792 => "10111100",7793 => "10001010",7794 => "00111111",7795 => "11111010",7796 => "00001111",7797 => "10110000",7798 => "11110011",7799 => "10110011",7800 => "10111000",7801 => "11000110",7802 => "01101100",7803 => "00001000",7804 => "11011000",7805 => "10010011",7806 => "01001111",7807 => "11011001",7808 => "11011100",7809 => "00010000",7810 => "00001010",7811 => "00100100",7812 => "11111011",7813 => "10011011",7814 => "00111000",7815 => "00011111",7816 => "01110000",7817 => "10010010",7818 => "11000101",7819 => "00011011",7820 => "10110001",7821 => "10011010",7822 => "10000010",7823 => "00110110",7824 => "11101111",7825 => "10000111",7826 => "01010011",7827 => "11010000",7828 => "00000011",7829 => "10000111",7830 => "11111101",7831 => "10001110",7832 => "10000111",7833 => "01000011",7834 => "10101101",7835 => "10011101",7836 => "10111001",7837 => "11000001",7838 => "10110011",7839 => "00001011",7840 => "10001101",7841 => "01110001",7842 => "11001111",7843 => "10101111",7844 => "01111110",7845 => "00101000",7846 => "00010111",7847 => "01000000",7848 => "00010011",7849 => "11111010",7850 => "01010111",7851 => "11011001",7852 => "11010011",7853 => "11000001",7854 => "10101100",7855 => "01000101",7856 => "00100110",7857 => "00011010",7858 => "11100101",7859 => "00101110",7860 => "01011100",7861 => "11001111",7862 => "00100101",7863 => "10100100",7864 => "00111011",7865 => "00000110",7866 => "10101100",7867 => "01000100",7868 => "10011010",7869 => "00010010",7870 => "00110111",7871 => "01010101",7872 => "01000110",7873 => "11000010",7874 => "11001011",7875 => "01100110",7876 => "01010000",7877 => "10001000",7878 => "11001101",7879 => "11111100",7880 => "11101101",7881 => "10011101",7882 => "01010000",7883 => "10001111",7884 => "10100011",7885 => "11000101",7886 => "00110000",7887 => "01000001",7888 => "01000001",7889 => "10000101",7890 => "11110101",7891 => "00010000",7892 => "01010010",7893 => "10010011",7894 => "00000110",7895 => "01010100",7896 => "01001101",7897 => "01101011",7898 => "11001100",7899 => "11111000",7900 => "01001101",7901 => "00111100",7902 => "11001010",7903 => "00111101",7904 => "11111111",7905 => "10010010",7906 => "11000011",7907 => "01111110",7908 => "11000110",7909 => "10011000",7910 => "01000011",7911 => "01011101",7912 => "11100101",7913 => "10011011",7914 => "01100111",7915 => "10001100",7916 => "00101000",7917 => "01110110",7918 => "00101000",7919 => "11100000",7920 => "00011010",7921 => "01100110",7922 => "11000000",7923 => "10010110",7924 => "01111111",7925 => "10011101",7926 => "01100011",7927 => "00100010",7928 => "10101010",7929 => "11110001",7930 => "00010111",7931 => "10111100",7932 => "01101101",7933 => "10000100",7934 => "00000011",7935 => "10100111",7936 => "01111000",7937 => "10110110",7938 => "00110010",7939 => "10101011",7940 => "01100011",7941 => "10011111",7942 => "11001100",7943 => "11100011",7944 => "01110011",7945 => "10101011",7946 => "01000111",7947 => "00010100",7948 => "00110111",7949 => "00100011",7950 => "11111000",7951 => "11111010",7952 => "01100011",7953 => "11010111",7954 => "00000010",7955 => "10000001",7956 => "10001000",7957 => "00001100",7958 => "11101010",7959 => "11011000",7960 => "00001101",7961 => "00010111",7962 => "01111100",7963 => "11010100",7964 => "10101100",7965 => "01011101",7966 => "00001111",7967 => "11011011",7968 => "00001011",7969 => "00001110",7970 => "11010101",7971 => "01010101",7972 => "10010010",7973 => "11100010",7974 => "11100010",7975 => "00100011",7976 => "10000000",7977 => "10000100",7978 => "10010110",7979 => "10011110",7980 => "00011111",7981 => "00110001",7982 => "11001010",7983 => "00101101",7984 => "00000101",7985 => "11001110",7986 => "10101011",7987 => "00110101",7988 => "10001001",7989 => "01100011",7990 => "10000011",7991 => "10001001",7992 => "00000101",7993 => "11010010",7994 => "10110001",7995 => "11100010",7996 => "01100010",7997 => "00011101",7998 => "00001101",7999 => "10010010",8000 => "10110000",8001 => "01111111",8002 => "11011110",8003 => "00100100",8004 => "10111101",8005 => "00101110",8006 => "00100010",8007 => "11010001",8008 => "00100000",8009 => "01001000",8010 => "01110010",8011 => "10010110",8012 => "11101011",8013 => "01100110",8014 => "00110011",8015 => "10110101",8016 => "01110110",8017 => "00111011",8018 => "00101010",8019 => "00000000",8020 => "01100100",8021 => "01011110",8022 => "11000111",8023 => "00000011",8024 => "11001001",8025 => "00111101",8026 => "00011001",8027 => "00011001",8028 => "10110010",8029 => "11100111",8030 => "10111100",8031 => "10001110",8032 => "01111001",8033 => "00010000",8034 => "01101101",8035 => "00111111",8036 => "01011001",8037 => "10010001",8038 => "00100011",8039 => "10100111",8040 => "00101001",8041 => "01011011",8042 => "00010001",8043 => "10011001",8044 => "10000101",8045 => "00111101",8046 => "11111000",8047 => "10001101",8048 => "00001000",8049 => "00110011",8050 => "11111100",8051 => "00011011",8052 => "00111101",8053 => "01100100",8054 => "11011001",8055 => "11001000",8056 => "01100111",8057 => "10111110",8058 => "10011100",8059 => "11101001",8060 => "01011100",8061 => "11111101",8062 => "11001011",8063 => "10000001",8064 => "10001001",8065 => "01110001",8066 => "01111111",8067 => "01000010",8068 => "11101000",8069 => "00000000",8070 => "11110100",8071 => "10110100",8072 => "00011000",8073 => "10101101",8074 => "01011010",8075 => "01101001",8076 => "11110011",8077 => "00011101",8078 => "01001000",8079 => "00100001",8080 => "00010010",8081 => "01000110",8082 => "10011011",8083 => "01011000",8084 => "00100001",8085 => "10011100",8086 => "10110001",8087 => "00111101",8088 => "00010010",8089 => "00111010",8090 => "00000100",8091 => "10001110",8092 => "10000000",8093 => "00011101",8094 => "00000010",8095 => "00000110",8096 => "00111111",8097 => "01010000",8098 => "11011000",8099 => "01011111",8100 => "00101110",8101 => "11000010",8102 => "00111110",8103 => "11110101",8104 => "10100010",8105 => "11110100",8106 => "10001100",8107 => "11000100",8108 => "01110101",8109 => "10111010",8110 => "10111101",8111 => "01011001",8112 => "01001111",8113 => "10000100",8114 => "11010100",8115 => "01010010",8116 => "10101101",8117 => "10110101",8118 => "11111000",8119 => "00010010",8120 => "11110001",8121 => "01100000",8122 => "01100000",8123 => "01011100",8124 => "00000101",8125 => "01110010",8126 => "01001000",8127 => "01101101",8128 => "01001110",8129 => "10011111",8130 => "11011001",8131 => "00100101",8132 => "10110101",8133 => "00111111",8134 => "01110101",8135 => "01001101",8136 => "01001001",8137 => "01000000",8138 => "11111010",8139 => "11000101",8140 => "11001000",8141 => "11011110",8142 => "11111111",8143 => "01110010",8144 => "10001100",8145 => "01011001",8146 => "11101000",8147 => "00110001",8148 => "10011110",8149 => "00010111",8150 => "11111000",8151 => "11101001",8152 => "01110011",8153 => "01011000",8154 => "00111000",8155 => "01100010",8156 => "01111101",8157 => "11110001",8158 => "10000000",8159 => "01100011",8160 => "00110011",8161 => "11100011",8162 => "11000101",8163 => "00111110",8164 => "01001010",8165 => "11000000",8166 => "10000100",8167 => "10110001",8168 => "11111101",8169 => "01010100",8170 => "01100111",8171 => "10111101",8172 => "00001001",8173 => "11110001",8174 => "10110110",8175 => "10100001",8176 => "01010100",8177 => "00100100",8178 => "00111000",8179 => "01000010",8180 => "01101101",8181 => "10100101",8182 => "11110011",8183 => "01011000",8184 => "10111101",8185 => "11111101",8186 => "00010110",8187 => "10011000",8188 => "10101010",8189 => "01000110",8190 => "11001011",8191 => "10110101",8192 => "01111010",8193 => "00100000",8194 => "10101100",8195 => "10010001",8196 => "10100011",8197 => "10011101",8198 => "01101001",8199 => "10010000",8200 => "10101110",8201 => "11101110",8202 => "11000000",8203 => "10011111",8204 => "10111111",8205 => "00101110",8206 => "11100101",8207 => "10011010",8208 => "10011100",8209 => "11000000",8210 => "10110000",8211 => "00000001",8212 => "00100110",8213 => "00111000",8214 => "10101001",8215 => "11111010",8216 => "10000010",8217 => "11001101",8218 => "10000101",8219 => "11110010",8220 => "10101010",8221 => "00010010",8222 => "01010011",8223 => "00110110",8224 => "11111010",8225 => "00111111",8226 => "11100000",8227 => "00011000",8228 => "00110101",8229 => "00100111",8230 => "11111000",8231 => "01100000",8232 => "10100010",8233 => "10000110",8234 => "00010011",8235 => "11101010",8236 => "01001001",8237 => "10010000",8238 => "01010111",8239 => "01011100",8240 => "00010110",8241 => "00001001",8242 => "11001010",8243 => "00100100",8244 => "01000011",8245 => "00111010",8246 => "10000010",8247 => "01111101",8248 => "01100001",8249 => "00101100",8250 => "11000011",8251 => "10010011",8252 => "10100011",8253 => "10110001",8254 => "11000100",8255 => "01110000",8256 => "11111011",8257 => "00110001",8258 => "11110010",8259 => "10001111",8260 => "10110100",8261 => "00001000",8262 => "00100101",8263 => "00001101",8264 => "10000110",8265 => "01001011",8266 => "01100100",8267 => "00011010",8268 => "10101100",8269 => "00011000",8270 => "11011011",8271 => "01001000",8272 => "10011011",8273 => "00011100",8274 => "11000001",8275 => "10000001",8276 => "01000011",8277 => "00111001",8278 => "01110000",8279 => "00000110",8280 => "11111111",8281 => "10000101",8282 => "10101010",8283 => "01110110",8284 => "11000011",8285 => "01011110",8286 => "00110101",8287 => "01101110",8288 => "00000001",8289 => "11010010",8290 => "01001010",8291 => "11000111",8292 => "00100000",8293 => "01100111",8294 => "00110101",8295 => "00100101",8296 => "11001001",8297 => "00001101",8298 => "01101101",8299 => "10110010",8300 => "01010010",8301 => "01101001",8302 => "11010100",8303 => "00010110",8304 => "11010100",8305 => "11100100",8306 => "11100110",8307 => "00100111",8308 => "00011100",8309 => "11110000",8310 => "10011001",8311 => "11110011",8312 => "01110111",8313 => "00101011",8314 => "01100111",8315 => "01100010",8316 => "00010110",8317 => "01001111",8318 => "10110000",8319 => "01101011",8320 => "10000001",8321 => "00111100",8322 => "01010000",8323 => "01110000",8324 => "00100111",8325 => "00101000",8326 => "11100010",8327 => "00000010",8328 => "11101000",8329 => "00011010",8330 => "10000011",8331 => "11000011",8332 => "11001111",8333 => "10010000",8334 => "10000111",8335 => "10010010",8336 => "01101111",8337 => "10100010",8338 => "01111000",8339 => "00001110",8340 => "10111001",8341 => "11010001",8342 => "01011010",8343 => "01101011",8344 => "01011010",8345 => "10110001",8346 => "11001000",8347 => "01010100",8348 => "01000001",8349 => "01010111",8350 => "11000001",8351 => "01101000",8352 => "00100010",8353 => "01101011",8354 => "01101011",8355 => "10001111",8356 => "01000010",8357 => "11110110",8358 => "01100101",8359 => "11001010",8360 => "11000011",8361 => "01101101",8362 => "01010001",8363 => "00100101",8364 => "11011011",8365 => "00001011",8366 => "10001011",8367 => "00101001",8368 => "00001110",8369 => "00000111",8370 => "10111001",8371 => "11111110",8372 => "00010100",8373 => "11010001",8374 => "00110111",8375 => "10011111",8376 => "01100001",8377 => "00101110",8378 => "01001101",8379 => "11100010",8380 => "11011000",8381 => "10111001",8382 => "00010101",8383 => "10000010",8384 => "01101010",8385 => "10000010",8386 => "10011001",8387 => "00011111",8388 => "00010001",8389 => "11010101",8390 => "00101100",8391 => "10001111",8392 => "01100000",8393 => "00001100",8394 => "10101001",8395 => "11100010",8396 => "11001010",8397 => "00110100",8398 => "01110000",8399 => "10001001",8400 => "11001011",8401 => "00010011",8402 => "10110010",8403 => "11111110",8404 => "00001111",8405 => "11101110",8406 => "11110111",8407 => "10001011",8408 => "11011000",8409 => "11000001",8410 => "00011000",8411 => "01001001",8412 => "01000000",8413 => "00001010",8414 => "01110101",8415 => "10100101",8416 => "11100111",8417 => "01001000",8418 => "01100110",8419 => "10110000",8420 => "00111010",8421 => "00000111",8422 => "00110100",8423 => "10101001",8424 => "10001110",8425 => "00101111",8426 => "10100100",8427 => "01100000",8428 => "00111110",8429 => "10111110",8430 => "11000111",8431 => "01001111",8432 => "11001111",8433 => "00101111",8434 => "11010110",8435 => "01000011",8436 => "01001010",8437 => "11011111",8438 => "01011000",8439 => "10000110",8440 => "10110101",8441 => "10011101",8442 => "00010101",8443 => "10111111",8444 => "00011000",8445 => "11010110",8446 => "00011011",8447 => "11000000",8448 => "01001001",8449 => "00000000",8450 => "00100100",8451 => "10100100",8452 => "01010001",8453 => "10010111",8454 => "00100111",8455 => "10101111",8456 => "01000010",8457 => "00111100",8458 => "11110100",8459 => "10011011",8460 => "10101100",8461 => "10111001",8462 => "11111110",8463 => "11111011",8464 => "10101000",8465 => "11101111",8466 => "01011001",8467 => "00111001",8468 => "01101010",8469 => "11101110",8470 => "01100011",8471 => "01000110",8472 => "11000011",8473 => "10011000",8474 => "11010101",8475 => "10100110",8476 => "01101011",8477 => "10011111",8478 => "01011001",8479 => "11000100",8480 => "01110001",8481 => "00001101",8482 => "00101100",8483 => "11001011",8484 => "00110001",8485 => "01010100",8486 => "01011010",8487 => "01101100",8488 => "00110111",8489 => "11010010",8490 => "01001110",8491 => "11000011",8492 => "01001110",8493 => "00101111",8494 => "01101001",8495 => "11110010",8496 => "00001010",8497 => "01100000",8498 => "01001001",8499 => "10110111",8500 => "10010000",8501 => "10010011",8502 => "11011000",8503 => "11101101",8504 => "01100100",8505 => "10111101",8506 => "10111111",8507 => "00001001",8508 => "01100101",8509 => "01010101",8510 => "11100001",8511 => "10011010",8512 => "01000101",8513 => "00010011",8514 => "11111100",8515 => "11100001",8516 => "11000011",8517 => "00001011",8518 => "00110010",8519 => "11100010",8520 => "11001001",8521 => "11001011",8522 => "00110011",8523 => "11001111",8524 => "01000111",8525 => "10100011",8526 => "01011011",8527 => "00110011",8528 => "01001110",8529 => "01010111",8530 => "10111101",8531 => "00101010",8532 => "11101110",8533 => "11101111",8534 => "00000001",8535 => "00110010",8536 => "10101010",8537 => "01100101",8538 => "10101100",8539 => "01100000",8540 => "00111010",8541 => "11001000",8542 => "10000101",8543 => "10100101",8544 => "01000101",8545 => "00000000",8546 => "00011100",8547 => "00011001",8548 => "00100110",8549 => "01110100",8550 => "11011110",8551 => "10111101",8552 => "11111101",8553 => "01101101",8554 => "00101011",8555 => "00100101",8556 => "00001010",8557 => "10110110",8558 => "11010010",8559 => "00100110",8560 => "01111011",8561 => "10000110",8562 => "00110000",8563 => "11010110",8564 => "00000111",8565 => "00000111",8566 => "01111001",8567 => "11001100",8568 => "10111110",8569 => "11111110",8570 => "11010111",8571 => "01101010",8572 => "11111110",8573 => "10010001",8574 => "00011001",8575 => "11010001",8576 => "10001100",8577 => "10101100",8578 => "11110111",8579 => "10011011",8580 => "10101111",8581 => "00101010",8582 => "10010010",8583 => "10010111",8584 => "11011010",8585 => "00010101",8586 => "10111001",8587 => "11011100",8588 => "01011010",8589 => "11000100",8590 => "11001101",8591 => "11010111",8592 => "11011110",8593 => "11000111",8594 => "11101110",8595 => "01001100",8596 => "11010000",8597 => "10011100",8598 => "01000100",8599 => "00001011",8600 => "11101100",8601 => "10011011",8602 => "01011001",8603 => "11110010",8604 => "11101001",8605 => "00111110",8606 => "10110110",8607 => "00100101",8608 => "10011011",8609 => "11000001",8610 => "00011110",8611 => "10101101",8612 => "01100000",8613 => "10110110",8614 => "10011001",8615 => "01111000",8616 => "10010101",8617 => "11100101",8618 => "01100100",8619 => "00100011",8620 => "00101001",8621 => "00010111",8622 => "01000110",8623 => "00100110",8624 => "00101001",8625 => "10100010",8626 => "01001111",8627 => "10011011",8628 => "01110100",8629 => "01110010",8630 => "11101011",8631 => "01101101",8632 => "10010101",8633 => "10100110",8634 => "00001100",8635 => "11111111",8636 => "11110101",8637 => "01110101",8638 => "00111010",8639 => "00111001",8640 => "11111111",8641 => "01001101",8642 => "00010111",8643 => "11110110",8644 => "11111000",8645 => "10100001",8646 => "00110010",8647 => "01011010",8648 => "11000001",8649 => "11100001",8650 => "01011101",8651 => "10111110",8652 => "01101011",8653 => "00011001",8654 => "01110010",8655 => "00000010",8656 => "01110000",8657 => "01010100",8658 => "11010001",8659 => "00010001",8660 => "10001000",8661 => "11110000",8662 => "11000101",8663 => "11000101",8664 => "01001111",8665 => "01100001",8666 => "11011001",8667 => "00010000",8668 => "01111011",8669 => "11001011",8670 => "11000110",8671 => "10111011",8672 => "01001010",8673 => "01011111",8674 => "10111100",8675 => "00010001",8676 => "00011101",8677 => "01001010",8678 => "01101011",8679 => "11001001",8680 => "00010000",8681 => "00101100",8682 => "00110011",8683 => "01010011",8684 => "01000101",8685 => "00111000",8686 => "01011010",8687 => "01000110",8688 => "01001100",8689 => "10100000",8690 => "10011011",8691 => "11110110",8692 => "01010101",8693 => "10000110",8694 => "01101000",8695 => "00110111",8696 => "10111100",8697 => "10010011",8698 => "10001000",8699 => "10110101",8700 => "10000101",8701 => "01111000",8702 => "10011001",8703 => "11010100",8704 => "00100100",8705 => "10101111",8706 => "10010110",8707 => "00001101",8708 => "00010000",8709 => "00100000",8710 => "10011001",8711 => "01011010",8712 => "00001000",8713 => "10010011",8714 => "00000101",8715 => "00011101",8716 => "10000111",8717 => "10101100",8718 => "10001011",8719 => "11110110",8720 => "01101000",8721 => "10011111",8722 => "11101110",8723 => "01110100",8724 => "00001011",8725 => "10011101",8726 => "10111010",8727 => "01010000",8728 => "11111111",8729 => "00111110",8730 => "11111010",8731 => "01111100",8732 => "00111010",8733 => "01011110",8734 => "11001000",8735 => "10001101",8736 => "11111111",8737 => "00101101",8738 => "11110111",8739 => "00110111",8740 => "00000111",8741 => "11100110",8742 => "10110100",8743 => "11110100",8744 => "10011010",8745 => "11001000",8746 => "11000110",8747 => "10101101",8748 => "11110001",8749 => "11110010",8750 => "10010101",8751 => "01111111",8752 => "10100100",8753 => "01101111",8754 => "01110111",8755 => "10110111",8756 => "11110101",8757 => "10110010",8758 => "00111001",8759 => "10111100",8760 => "00110001",8761 => "00000100",8762 => "01000111",8763 => "01000100",8764 => "10100001",8765 => "10110011",8766 => "11100101",8767 => "10011011",8768 => "10101111",8769 => "01100010",8770 => "00100101",8771 => "01001001",8772 => "01110000",8773 => "10111110",8774 => "00000010",8775 => "11100101",8776 => "10101011",8777 => "10100001",8778 => "01001100",8779 => "01111101",8780 => "10100011",8781 => "10011101",8782 => "01111110",8783 => "01110101",8784 => "11001110",8785 => "00000011",8786 => "01001010",8787 => "11000010",8788 => "00010110",8789 => "01010100",8790 => "01001001",8791 => "11110111",8792 => "01111110",8793 => "00001001",8794 => "01110011",8795 => "11111001",8796 => "00100111",8797 => "01011011",8798 => "01101011",8799 => "10110010",8800 => "00011010",8801 => "00110010",8802 => "01100100",8803 => "00000111",8804 => "10110100",8805 => "11001011",8806 => "00100100",8807 => "01111100",8808 => "01101000",8809 => "11100100",8810 => "01010011",8811 => "10110111",8812 => "01101100",8813 => "00101111",8814 => "00010100",8815 => "00011011",8816 => "11010100",8817 => "00000101",8818 => "00010001",8819 => "10000011",8820 => "01100010",8821 => "11000000",8822 => "00010111",8823 => "11101101",8824 => "11000111",8825 => "10101101",8826 => "01011001",8827 => "10001000",8828 => "10111111",8829 => "11110110",8830 => "01111000",8831 => "11110000",8832 => "00101101",8833 => "10111001",8834 => "10110010",8835 => "00010110",8836 => "11001110",8837 => "01101001",8838 => "10011110",8839 => "10110101",8840 => "11111111",8841 => "01011010",8842 => "10001001",8843 => "11101110",8844 => "00100100",8845 => "10000100",8846 => "10010110",8847 => "00010110",8848 => "01111101",8849 => "11011110",8850 => "00111111",8851 => "01100111",8852 => "11000011",8853 => "00100101",8854 => "01110000",8855 => "00111000",8856 => "11010011",8857 => "11111110",8858 => "10111001",8859 => "00111110",8860 => "11100111",8861 => "01111101",8862 => "11101000",8863 => "00010110",8864 => "01100011",8865 => "11001000",8866 => "00111111",8867 => "11000000",8868 => "00010101",8869 => "11001100",8870 => "00111001",8871 => "10101001",8872 => "10000001",8873 => "00010111",8874 => "00110011",8875 => "11010001",8876 => "10111001",8877 => "00001110",8878 => "01000000",8879 => "11110010",8880 => "01011101",8881 => "00011011",8882 => "10111111",8883 => "10100100",8884 => "11110000",8885 => "00110010",8886 => "00011001",8887 => "10001111",8888 => "01100101",8889 => "11110100",8890 => "01000000",8891 => "00110001",8892 => "00110110",8893 => "10001100",8894 => "01000011",8895 => "01101110",8896 => "10011000",8897 => "00001110",8898 => "10010011",8899 => "11010001",8900 => "11110110",8901 => "01111011",8902 => "11110101",8903 => "00001010",8904 => "11010100",8905 => "11011011",8906 => "11010110",8907 => "10110000",8908 => "01011011",8909 => "11001100",8910 => "00110101",8911 => "01010000",8912 => "11100010",8913 => "00101111",8914 => "10011000",8915 => "01111101",8916 => "11010100",8917 => "00101110",8918 => "10111101",8919 => "01100011",8920 => "00110010",8921 => "00110100",8922 => "00110010",8923 => "10110010",8924 => "10011101",8925 => "10100101",8926 => "01000010",8927 => "11001100",8928 => "11000101",8929 => "00000000",8930 => "00110000",8931 => "10010110",8932 => "10111001",8933 => "11100001",8934 => "00001101",8935 => "01010110",8936 => "11101000",8937 => "00001110",8938 => "00101101",8939 => "11101001",8940 => "11100000",8941 => "11011011",8942 => "10011101",8943 => "01001000",8944 => "10111101",8945 => "11100101",8946 => "10111110",8947 => "01101010",8948 => "00100001",8949 => "11011011",8950 => "01011111",8951 => "10111001",8952 => "01100111",8953 => "01001111",8954 => "01110101",8955 => "11011110",8956 => "01010001",8957 => "01101101",8958 => "10111110",8959 => "00101011",8960 => "00000110",8961 => "11110110",8962 => "01011000",8963 => "10100111",8964 => "10001011",8965 => "11000000",8966 => "00000010",8967 => "10111101",8968 => "11011001",8969 => "00000010",8970 => "00000111",8971 => "11010100",8972 => "00011110",8973 => "11111100",8974 => "01011110",8975 => "11010100",8976 => "01100111",8977 => "11000111",8978 => "10100011",8979 => "00110101",8980 => "11110001",8981 => "10111001",8982 => "11011000",8983 => "10111111",8984 => "00000101",8985 => "10100011",8986 => "10100110",8987 => "00001111",8988 => "01010001",8989 => "10100011",8990 => "10000010",8991 => "01001100",8992 => "10110010",8993 => "11000001",8994 => "01001111",8995 => "00101111",8996 => "11000100",8997 => "10011110",8998 => "01000010",8999 => "10010001",9000 => "10001000",9001 => "01101101",9002 => "10001100",9003 => "01101110",9004 => "00001100",9005 => "11001011",9006 => "10000111",9007 => "11101100",9008 => "10000111",9009 => "00000010",9010 => "01000010",9011 => "10110010",9012 => "11110101",9013 => "10011011",9014 => "01000001",9015 => "10110011",9016 => "10000011",9017 => "11101101",9018 => "00110100",9019 => "11010010",9020 => "00111000",9021 => "01100111",9022 => "10110100",9023 => "11010011",9024 => "01101001",9025 => "11111010",9026 => "11110000",9027 => "00101010",9028 => "01000101",9029 => "11001100",9030 => "01011000",9031 => "10101001",9032 => "01000000",9033 => "11100100",9034 => "00011001",9035 => "00101101",9036 => "11000111",9037 => "10101110",9038 => "00010110",9039 => "11110010",9040 => "01010111",9041 => "11111101",9042 => "00101110",9043 => "00001101",9044 => "01011101",9045 => "11111101",9046 => "00001110",9047 => "00100100",9048 => "00110001",9049 => "11100110",9050 => "11010011",9051 => "01010100",9052 => "11100010",9053 => "11010101",9054 => "00110011",9055 => "11000010",9056 => "01101101",9057 => "10100101",9058 => "11000110",9059 => "11000011",9060 => "01010011",9061 => "01000010",9062 => "00001001",9063 => "10101101",9064 => "10001001",9065 => "01011010",9066 => "01010100",9067 => "10001000",9068 => "01001111",9069 => "00101100",9070 => "10100010",9071 => "00111110",9072 => "11110101",9073 => "00011100",9074 => "11010010",9075 => "10101100",9076 => "11011110",9077 => "11010011",9078 => "10011010",9079 => "00000100",9080 => "01011101",9081 => "01100001",9082 => "10100000",9083 => "00111100",9084 => "10110111",9085 => "10110111",9086 => "01110000",9087 => "10001101",9088 => "00010111",9089 => "10111011",9090 => "00011000",9091 => "00010011",9092 => "00001100",9093 => "00010110",9094 => "01001010",9095 => "01001101",9096 => "10010110",9097 => "00001111",9098 => "01111011",9099 => "01010110",9100 => "01001111",9101 => "01000000",9102 => "01100011",9103 => "01100110",9104 => "00100000",9105 => "01001001",9106 => "00100010",9107 => "11010001",9108 => "11110101",9109 => "10000011",9110 => "00000110",9111 => "10101010",9112 => "10111000",9113 => "10110110",9114 => "00101101",9115 => "01111000",9116 => "00011010",9117 => "00111111",9118 => "01001000",9119 => "00111010",9120 => "01111011",9121 => "11001100",9122 => "10010101",9123 => "01101110",9124 => "01100110",9125 => "00000000",9126 => "01110100",9127 => "11111100",9128 => "11110100",9129 => "10100001",9130 => "00110001",9131 => "00110011",9132 => "00111001",9133 => "00010101",9134 => "01010001",9135 => "00010110",9136 => "10000011",9137 => "00001010",9138 => "11100100",9139 => "11100000",9140 => "00000001",9141 => "11010110",9142 => "00001100",9143 => "01101100",9144 => "11001100",9145 => "01111100",9146 => "10111001",9147 => "01101110",9148 => "01111111",9149 => "11011000",9150 => "01111000",9151 => "00110011",9152 => "01110100",9153 => "01010111",9154 => "01111101",9155 => "11101111",9156 => "11110011",9157 => "11110010",9158 => "11101011",9159 => "00101000",9160 => "11110000",9161 => "11010011",9162 => "11100100",9163 => "01000010",9164 => "00100100",9165 => "11100100",9166 => "11110100",9167 => "10111010",9168 => "10010000",9169 => "00100000",9170 => "00110100",9171 => "10100101",9172 => "01101101",9173 => "01101010",9174 => "10010011",9175 => "01100100",9176 => "01010011",9177 => "11001100",9178 => "01100110",9179 => "01001011",9180 => "01100110",9181 => "10001001",9182 => "10010010",9183 => "11110110",9184 => "01011100",9185 => "11110010",9186 => "00011110",9187 => "01100110",9188 => "10001000",9189 => "10001001",9190 => "11001001",9191 => "10110110",9192 => "01101001",9193 => "01111000",9194 => "00011111",9195 => "10100100",9196 => "10100001",9197 => "01010000",9198 => "00110110",9199 => "00001101",9200 => "11111011",9201 => "01111110",9202 => "00001011",9203 => "00010101",9204 => "11001101",9205 => "00001011",9206 => "01110000",9207 => "11111101",9208 => "01101100",9209 => "11100010",9210 => "11010100",9211 => "11101111",9212 => "00111111",9213 => "10001100",9214 => "01101000",9215 => "01111101",9216 => "01100010",9217 => "01011110",9218 => "10010011",9219 => "01100101",9220 => "01100101",9221 => "01110000",9222 => "10001100",9223 => "00000010",9224 => "00011111",9225 => "11111111",9226 => "00101000",9227 => "10111111",9228 => "10101000",9229 => "11001010",9230 => "11110111",9231 => "11100001",9232 => "00110011",9233 => "10100111",9234 => "00001111",9235 => "00110110",9236 => "00001010",9237 => "10011100",9238 => "11110111",9239 => "00110111",9240 => "11110011",9241 => "11101010",9242 => "00011100",9243 => "11001111",9244 => "01010111",9245 => "11010000",9246 => "10100010",9247 => "10000001",9248 => "00001100",9249 => "00010010",9250 => "00000000",9251 => "00110010",9252 => "11001011",9253 => "00010111",9254 => "01011100",9255 => "11101010",9256 => "11100010",9257 => "01001000",9258 => "11100101",9259 => "11110100",9260 => "11101110",9261 => "01000010",9262 => "10011110",9263 => "10001010",9264 => "11101010",9265 => "01101011",9266 => "11111101",9267 => "11100001",9268 => "11011001",9269 => "00101100",9270 => "00101100",9271 => "10101110",9272 => "10100001",9273 => "10110110",9274 => "11100110",9275 => "11110010",9276 => "00010010",9277 => "10110111",9278 => "01111001",9279 => "01100100",9280 => "00000000",9281 => "10001100",9282 => "11011010",9283 => "11001100",9284 => "11000100",9285 => "01000010",9286 => "11011111",9287 => "10100001",9288 => "10010010",9289 => "10010101",9290 => "01010111",9291 => "10100111",9292 => "01000101",9293 => "01100100",9294 => "00000101",9295 => "10001000",9296 => "11100010",9297 => "00001001",9298 => "10000101",9299 => "11011010",9300 => "01111001",9301 => "00111001",9302 => "10101110",9303 => "01001110",9304 => "01010011",9305 => "10011010",9306 => "10100011",9307 => "10000010",9308 => "11000000",9309 => "11010001",9310 => "10010010",9311 => "10110100",9312 => "00110001",9313 => "11100111",9314 => "00011011",9315 => "10111001",9316 => "01010100",9317 => "00011011",9318 => "01100101",9319 => "10010100",9320 => "11010111",9321 => "01100110",9322 => "11110101",9323 => "00010011",9324 => "11011100",9325 => "01101111",9326 => "10001001",9327 => "01001110",9328 => "00110000",9329 => "11000111",9330 => "10000111",9331 => "10111100",9332 => "11010100",9333 => "01110111",9334 => "10000000",9335 => "01001111",9336 => "00101111",9337 => "00111010",9338 => "10001111",9339 => "10101010",9340 => "10101000",9341 => "00010101",9342 => "10011111",9343 => "00011010",9344 => "10101110",9345 => "10110000",9346 => "11010110",9347 => "01101001",9348 => "00100101",9349 => "11100011",9350 => "00001111",9351 => "01110101",9352 => "11101001",9353 => "01011000",9354 => "01110111",9355 => "11100101",9356 => "01001100",9357 => "01010111",9358 => "01110000",9359 => "10001101",9360 => "00110110",9361 => "00101011",9362 => "01000010",9363 => "10011110",9364 => "10011011",9365 => "11001100",9366 => "11010010",9367 => "00001011",9368 => "01111010",9369 => "10001110",9370 => "10111101",9371 => "00111100",9372 => "11011110",9373 => "10010011",9374 => "01000010",9375 => "00100010",9376 => "10011000",9377 => "11010000",9378 => "11010100",9379 => "01011010",9380 => "11111111",9381 => "11101111",9382 => "10000011",9383 => "01110111",9384 => "00111110",9385 => "01011111",9386 => "00100000",9387 => "00101111",9388 => "01000000",9389 => "10100001",9390 => "00101101",9391 => "01001001",9392 => "00101011",9393 => "11010110",9394 => "10101110",9395 => "01111000",9396 => "11001010",9397 => "00100010",9398 => "00010101",9399 => "00011101",9400 => "00000000",9401 => "00010100",9402 => "11110010",9403 => "00111100",9404 => "00011111",9405 => "10011111",9406 => "00011000",9407 => "00111111",9408 => "01111101",9409 => "11010100",9410 => "10011011",9411 => "01101010",9412 => "11000110",9413 => "01100111",9414 => "00011111",9415 => "01000001",9416 => "10001110",9417 => "11000011",9418 => "11010000",9419 => "01111001",9420 => "00000100",9421 => "10111111",9422 => "00111101",9423 => "00011101",9424 => "00001100",9425 => "00011010",9426 => "11101011",9427 => "11110010",9428 => "00110000",9429 => "00101001",9430 => "01010110",9431 => "01101001",9432 => "11101001",9433 => "00100111",9434 => "10000110",9435 => "10000011",9436 => "10111001",9437 => "10111010",9438 => "00111110",9439 => "00010010",9440 => "11100010",9441 => "10101110",9442 => "10010110",9443 => "00011010",9444 => "00000110",9445 => "00001011",9446 => "00110011",9447 => "10011010",9448 => "00011111",9449 => "01001001",9450 => "10111010",9451 => "01110110",9452 => "00000110",9453 => "00011000",9454 => "10011100",9455 => "11100011",9456 => "00101000",9457 => "10110001",9458 => "01110000",9459 => "01001001",9460 => "10000011",9461 => "01110110",9462 => "00111101",9463 => "00000000",9464 => "00001011",9465 => "10101111",9466 => "00100001",9467 => "10000011",9468 => "00110000",9469 => "01111000",9470 => "00101011",9471 => "01101100",9472 => "11011111",9473 => "00000111",9474 => "01110111",9475 => "00001101",9476 => "11000001",9477 => "01111001",9478 => "01010100",9479 => "00111110",9480 => "00001101",9481 => "10000100",9482 => "00011000",9483 => "10100100",9484 => "11101011",9485 => "11010100",9486 => "00011001",9487 => "11110111",9488 => "00011001",9489 => "00110010",9490 => "00000001",9491 => "10001000",9492 => "11011100",9493 => "00010011",9494 => "10110101",9495 => "00001101",9496 => "00100011",9497 => "10001110",9498 => "10011111",9499 => "00111100",9500 => "01010000",9501 => "10100111",9502 => "01101101",9503 => "11110001",9504 => "10011011",9505 => "11110100",9506 => "00011011",9507 => "01010010",9508 => "11100011",9509 => "11101001",9510 => "10010100",9511 => "10000010",9512 => "10111111",9513 => "00111001",9514 => "11001010",9515 => "11011000",9516 => "01111011",9517 => "11100000",9518 => "10111010",9519 => "01001101",9520 => "10010110",9521 => "10000110",9522 => "01011010",9523 => "00111001",9524 => "01101010",9525 => "01110101",9526 => "00100101",9527 => "11011100",9528 => "11111110",9529 => "01101110",9530 => "10110100",9531 => "10111100",9532 => "00111110",9533 => "00111111",9534 => "11100011",9535 => "00100000",9536 => "11011010",9537 => "10111011",9538 => "01011001",9539 => "00101100",9540 => "11101010",9541 => "00100101",9542 => "11001101",9543 => "10111000",9544 => "11000111",9545 => "10011100",9546 => "00011100",9547 => "11010110",9548 => "01001011",9549 => "00101110",9550 => "10111011",9551 => "01000110",9552 => "10100110",9553 => "10110111",9554 => "10100110",9555 => "00001101",9556 => "11011111",9557 => "01100000",9558 => "00101011",9559 => "11000110",9560 => "01000000",9561 => "01110000",9562 => "00101101",9563 => "00100010",9564 => "01101100",9565 => "10101011",9566 => "11000011",9567 => "00010001",9568 => "10100000",9569 => "11010111",9570 => "11010011",9571 => "11100010",9572 => "11001110",9573 => "01010101",9574 => "10110100",9575 => "00011101",9576 => "00001010",9577 => "00111010",9578 => "11001001",9579 => "00101100",9580 => "00110001",9581 => "11101011",9582 => "11101000",9583 => "01111000",9584 => "10010100",9585 => "01001100",9586 => "11111001",9587 => "11100101",9588 => "10110011",9589 => "00101110",9590 => "00101101",9591 => "10001100",9592 => "11011110",9593 => "11001100",9594 => "00101111",9595 => "01011111",9596 => "00100001",9597 => "00011100",9598 => "00010001",9599 => "00111011",9600 => "10010110",9601 => "01001110",9602 => "01010111",9603 => "11100011",9604 => "11111010",9605 => "10111110",9606 => "00001010",9607 => "00001011",9608 => "01000111",9609 => "01100101",9610 => "10011110",9611 => "11011010",9612 => "01100010",9613 => "00011100",9614 => "00011000",9615 => "10001100",9616 => "01000111",9617 => "10000110",9618 => "00001111",9619 => "10110111",9620 => "11111100",9621 => "00111110",9622 => "01110101",9623 => "10101000",9624 => "10011111",9625 => "10011101",9626 => "10000110",9627 => "00100000",9628 => "10001001",9629 => "01010110",9630 => "11011011",9631 => "01010001",9632 => "01110111",9633 => "01000011",9634 => "10010010",9635 => "01001101",9636 => "00111010",9637 => "00001100",9638 => "00001110",9639 => "10110100",9640 => "10001101",9641 => "10011101",9642 => "00000110",9643 => "01000000",9644 => "10001011",9645 => "10001100",9646 => "10011101",9647 => "01111101",9648 => "11011011",9649 => "00010001",9650 => "01000011",9651 => "01111001",9652 => "01101010",9653 => "10011100",9654 => "11011011",9655 => "10101000",9656 => "00111011",9657 => "00111111",9658 => "11110011",9659 => "10011011",9660 => "11100001",9661 => "00101000",9662 => "10010010",9663 => "01011001",9664 => "01010110",9665 => "11100001",9666 => "11101001",9667 => "11101011",9668 => "00001011",9669 => "01100011",9670 => "10111011",9671 => "00101100",9672 => "01001101",9673 => "11101011",9674 => "10110010",9675 => "00010101",9676 => "10100001",9677 => "10010000",9678 => "01000111",9679 => "01011001",9680 => "10010110",9681 => "01000100",9682 => "00011011",9683 => "01011000",9684 => "11101001",9685 => "10000011",9686 => "00010000",9687 => "01010110",9688 => "01000011",9689 => "11111101",9690 => "11101000",9691 => "01000100",9692 => "01011110",9693 => "00110001",9694 => "00011011",9695 => "11110100",9696 => "00110011",9697 => "10100100",9698 => "00101111",9699 => "00100111",9700 => "11000011",9701 => "01100100",9702 => "10011010",9703 => "01110010",9704 => "00010100",9705 => "11110010",9706 => "10010011",9707 => "10011001",9708 => "00000011",9709 => "01011011",9710 => "11100100",9711 => "00001100",9712 => "01001110",9713 => "00100111",9714 => "01101100",9715 => "11100111",9716 => "11101000",9717 => "11001011",9718 => "10010001",9719 => "00001111",9720 => "11011010",9721 => "00000111",9722 => "10111110",9723 => "00010001",9724 => "01111100",9725 => "00100111",9726 => "00000101",9727 => "11100110",9728 => "11011101",9729 => "11100011",9730 => "00011000",9731 => "00001101",9732 => "01110111",9733 => "00100011",9734 => "01110010",9735 => "11101011",9736 => "11111001",9737 => "10111100",9738 => "01001111",9739 => "10111100",9740 => "00010000",9741 => "00011101",9742 => "10111110",9743 => "11001010",9744 => "11011110",9745 => "01100101",9746 => "11011101",9747 => "10111101",9748 => "01101000",9749 => "10000000",9750 => "01001100",9751 => "01001010",9752 => "11100110",9753 => "01010111",9754 => "01000110",9755 => "10111101",9756 => "00101110",9757 => "01000010",9758 => "10111001",9759 => "01010100",9760 => "01011100",9761 => "01110101",9762 => "00110010",9763 => "10010011",9764 => "11000010",9765 => "01111010",9766 => "00100001",9767 => "10100011",9768 => "10111000",9769 => "10001000",9770 => "10100010",9771 => "11010010",9772 => "00110101",9773 => "10100110",9774 => "10000101",9775 => "00011010",9776 => "11100001",9777 => "11011110",9778 => "00011011",9779 => "01101110",9780 => "10111100",9781 => "01100110",9782 => "10010101",9783 => "01111111",9784 => "01010101",9785 => "01111001",9786 => "00000010",9787 => "00001001",9788 => "01100011",9789 => "00111110",9790 => "00011001",9791 => "11100101",9792 => "11101011",9793 => "11011111",9794 => "10010010",9795 => "01100100",9796 => "11100010",9797 => "11011001",9798 => "11000001",9799 => "00001101",9800 => "11110010",9801 => "10101110",9802 => "10010001",9803 => "00011000",9804 => "11011010",9805 => "11111110",9806 => "10100101",9807 => "01100100",9808 => "00110010",9809 => "11011110",9810 => "10010110",9811 => "00001111",9812 => "11011111",9813 => "11001110",9814 => "11111001",9815 => "11000010",9816 => "11011001",9817 => "00001000",9818 => "00011011",9819 => "01010111",9820 => "00100011",9821 => "01100111",9822 => "01111111",9823 => "11010000",9824 => "11110100",9825 => "11001011",9826 => "10001011",9827 => "01111001",9828 => "01111010",9829 => "00001000",9830 => "00111011",9831 => "11010111",9832 => "00111110",9833 => "10000110",9834 => "00001010",9835 => "10011111",9836 => "11110100",9837 => "00010011",9838 => "10011111",9839 => "10001001",9840 => "00001110",9841 => "00000001",9842 => "00011111",9843 => "01010111",9844 => "00011100",9845 => "11100110",9846 => "01011101",9847 => "11110010",9848 => "11001111",9849 => "11111110",9850 => "10010100",9851 => "01001110",9852 => "00100101",9853 => "10001011",9854 => "01000000",9855 => "10100100",9856 => "01010001",9857 => "01100000",9858 => "10101111",9859 => "01011011",9860 => "00111110",9861 => "01011100",9862 => "11100001",9863 => "00011011",9864 => "00111011",9865 => "10001001",9866 => "11001100",9867 => "10001101",9868 => "10111101",9869 => "11110101",9870 => "10011010",9871 => "11111101",9872 => "10000110",9873 => "01101010",9874 => "00101100",9875 => "00110111",9876 => "11001010",9877 => "10100111",9878 => "11100010",9879 => "01000110",9880 => "01011000",9881 => "00100110",9882 => "01001100",9883 => "00000011",9884 => "01100100",9885 => "00110110",9886 => "00101000",9887 => "01010010",9888 => "01111101",9889 => "00001100",9890 => "01110101",9891 => "11110101",9892 => "01010111",9893 => "01000111",9894 => "10111100",9895 => "10010011",9896 => "00011110",9897 => "11100001",9898 => "00101110",9899 => "01101001",9900 => "01101011",9901 => "00111000",9902 => "00110101",9903 => "00101100",9904 => "10110000",9905 => "11000100",9906 => "00011110",9907 => "10000010",9908 => "10111111",9909 => "00101000",9910 => "10010110",9911 => "11000101",9912 => "11000101",9913 => "00110011",9914 => "10111011",9915 => "00100000",9916 => "00010010",9917 => "01100001",9918 => "00110000",9919 => "11110100",9920 => "01001111",9921 => "01100101",9922 => "00110001",9923 => "10010001",9924 => "10110010",9925 => "10100001",9926 => "01110010",9927 => "11011010",9928 => "10101111",9929 => "11011011",9930 => "10110110",9931 => "01001011",9932 => "00111011",9933 => "10011001",9934 => "00001011",9935 => "01101011",9936 => "00010000",9937 => "00100110",9938 => "10100100",9939 => "11101110",9940 => "00000001",9941 => "00101101",9942 => "11111010",9943 => "01011000",9944 => "11100111",9945 => "11100101",9946 => "00010010",9947 => "11101001",9948 => "00011100",9949 => "01100011",9950 => "10010010",9951 => "00011000",9952 => "11100000",9953 => "11001111",9954 => "00000111",9955 => "01100101",9956 => "10111111",9957 => "01100010",9958 => "01011111",9959 => "01011010",9960 => "10001100",9961 => "01010001",9962 => "01100100",9963 => "00011001",9964 => "01101010",9965 => "10100011",9966 => "11111111",9967 => "10110010",9968 => "10101110",9969 => "01110001",9970 => "01100111",9971 => "10100101",9972 => "11000111",9973 => "00001101",9974 => "00010100",9975 => "01100010",9976 => "10000011",9977 => "01010010",9978 => "01101011",9979 => "10000001",9980 => "11100111",9981 => "01110110",9982 => "00110101",9983 => "10100011",9984 => "00010000",9985 => "11010100",9986 => "10101110",9987 => "10111010",9988 => "10100001",9989 => "10111111",9990 => "00111101",9991 => "10111110",9992 => "00010100",9993 => "11111100",9994 => "01011000",9995 => "01011111",9996 => "11110001",9997 => "11011001",9998 => "01111101",9999 => "01011101",10000 => "10111010",10001 => "01111101",10002 => "11101110",10003 => "01110010",10004 => "10100000",10005 => "11111101",10006 => "01110010",10007 => "10110101",10008 => "01001011",10009 => "01001101",10010 => "00111011",10011 => "01011110",10012 => "10001100",10013 => "11001101",10014 => "01110001",10015 => "00110011",10016 => "11001010",10017 => "00010101",10018 => "11101010",10019 => "01001010",10020 => "10101111",10021 => "00010010",10022 => "11000100",10023 => "10000100",10024 => "11010110",10025 => "01011101",10026 => "10010101",10027 => "01011010",10028 => "00101000",10029 => "11110011",10030 => "10000000",10031 => "10001111",10032 => "11100111",10033 => "00010111",10034 => "11001111",10035 => "10011001",10036 => "10000010",10037 => "10100010",10038 => "10101000",10039 => "10110100",10040 => "10100011",10041 => "10111100",10042 => "00111110",10043 => "10010011",10044 => "01110001",10045 => "00101000",10046 => "01100010",10047 => "00111101",10048 => "01010111",10049 => "01110011",10050 => "11010101",10051 => "11101100",10052 => "11100101",10053 => "01100000",10054 => "10001111",10055 => "01100000",10056 => "00110011",10057 => "00011110",10058 => "01110110",10059 => "01101100",10060 => "11001101",10061 => "01111011",10062 => "01001000",10063 => "11010100",10064 => "10111111",10065 => "11111000",10066 => "01011011",10067 => "11011011",10068 => "10110000",10069 => "00000010",10070 => "01000101",10071 => "11011101",10072 => "01001001",10073 => "11110100",10074 => "01111100",10075 => "01010010",10076 => "10010100",10077 => "00010000",10078 => "11010100",10079 => "11111010",10080 => "01101100",10081 => "10101110",10082 => "01110010",10083 => "10110010",10084 => "11111000",10085 => "11100000",10086 => "11001010",10087 => "01001000",10088 => "11001000",10089 => "01010010",10090 => "10100011",10091 => "11001111",10092 => "10010110",10093 => "01111001",10094 => "01111000",10095 => "11011100",10096 => "11000011",10097 => "11011101",10098 => "11000100",10099 => "11000001",10100 => "00011100",10101 => "11010010",10102 => "10010110",10103 => "00101110",10104 => "10111010",10105 => "01001110",10106 => "11101001",10107 => "01110000",10108 => "11010011",10109 => "11100001",10110 => "11000111",10111 => "10011010",10112 => "10001000",10113 => "11110000",10114 => "00111101",10115 => "01011110",10116 => "01110101",10117 => "01011000",10118 => "11110110",10119 => "11100000",10120 => "01110000",10121 => "01001011",10122 => "10101100",10123 => "10110110",10124 => "10010111",10125 => "10010001",10126 => "11010111",10127 => "01111111",10128 => "00101100",10129 => "01011101",10130 => "01101110",10131 => "01000110",10132 => "00100101",10133 => "00010110",10134 => "11100000",10135 => "01111100",10136 => "11010010",10137 => "00110111",10138 => "11010010",10139 => "10010001",10140 => "01111001",10141 => "11100100",10142 => "00100011",10143 => "00111110",10144 => "00011000",10145 => "00101011",10146 => "01101110",10147 => "01110101",10148 => "11110101",10149 => "10101011",10150 => "00001101",10151 => "11101100",10152 => "01111011",10153 => "10101111",10154 => "10111111",10155 => "00100110",10156 => "01000011",10157 => "00010000",10158 => "10101011",10159 => "11110100",10160 => "01100001",10161 => "01101100",10162 => "11101101",10163 => "01101010",10164 => "11001001",10165 => "11000011",10166 => "10100101",10167 => "01110100",10168 => "00110010",10169 => "11110101",10170 => "10010010",10171 => "10101010",10172 => "01011111",10173 => "11011101",10174 => "01111000",10175 => "00100011",10176 => "00101011",10177 => "11111011",10178 => "10101011",10179 => "00110110",10180 => "10010011",10181 => "00000000",10182 => "10111101",10183 => "00100011",10184 => "10010011",10185 => "00100100",10186 => "11111010",10187 => "00100001",10188 => "00010001",10189 => "01111110",10190 => "11010001",10191 => "00101100",10192 => "00110100",10193 => "00011101",10194 => "10000000",10195 => "00010111",10196 => "11110110",10197 => "00111110",10198 => "00011110",10199 => "00010100",10200 => "11001011",10201 => "01101100",10202 => "10110001",10203 => "10010011",10204 => "11010111",10205 => "10010100",10206 => "01111011",10207 => "00010101",10208 => "00011101",10209 => "01101001",10210 => "00011001",10211 => "11100001",10212 => "01110001",10213 => "10001101",10214 => "10010011",10215 => "01000101",10216 => "10011111",10217 => "00001001",10218 => "00111111",10219 => "11000111",10220 => "01010010",10221 => "00110100",10222 => "10100001",10223 => "01011010",10224 => "00100100",10225 => "01011001",10226 => "00101100",10227 => "10110010",10228 => "10001010",10229 => "10001011",10230 => "10101101",10231 => "10111011",10232 => "00011010",10233 => "01110100",10234 => "01110100",10235 => "00000101",10236 => "00101101",10237 => "10111111",10238 => "00110101",10239 => "10011110",10240 => "00010010",10241 => "01011111",10242 => "11011110",10243 => "10010101",10244 => "00100000",10245 => "11011101",10246 => "01111111",10247 => "11001101",10248 => "11000000",10249 => "11101001",10250 => "00100011",10251 => "10111100",10252 => "01001000",10253 => "01110100",10254 => "10100010",10255 => "10001101",10256 => "11111101",10257 => "11101101",10258 => "00001000",10259 => "11111111",10260 => "10011100",10261 => "10000111",10262 => "00101001",10263 => "10011101",10264 => "11101111",10265 => "10101110",10266 => "10011010",10267 => "01111110",10268 => "01100000",10269 => "00001101",10270 => "10101111",10271 => "00011110",10272 => "00010011",10273 => "11010100",10274 => "00001100",10275 => "11001010",10276 => "00110100",10277 => "01111000",10278 => "00010001",10279 => "11011110",10280 => "11100111",10281 => "00100000",10282 => "10110101",10283 => "10010000",10284 => "10111011",10285 => "01100101",10286 => "11110010",10287 => "00110111",10288 => "10010100",10289 => "10010111",10290 => "00010111",10291 => "10111000",10292 => "00010000",10293 => "11111010",10294 => "11000001",10295 => "10000101",10296 => "01111010",10297 => "00010000",10298 => "01110101",10299 => "00100111",10300 => "11001111",10301 => "11011010",10302 => "11011110",10303 => "00001100",10304 => "10101001",10305 => "11000011",10306 => "10101111",10307 => "10000110",10308 => "10111111",10309 => "00111010",10310 => "10111100",10311 => "00111000",10312 => "00110110",10313 => "11011000",10314 => "00011001",10315 => "10011100",10316 => "10101001",10317 => "01000110",10318 => "10100101",10319 => "10101101",10320 => "00111001",10321 => "11010100",10322 => "10010111",10323 => "00001000",10324 => "00110100",10325 => "00101110",10326 => "10100011",10327 => "01110111",10328 => "00010111",10329 => "01111000",10330 => "11110001",10331 => "11100111",10332 => "00010110",10333 => "10011000",10334 => "00001100",10335 => "11000111",10336 => "11111101",10337 => "00110010",10338 => "01111111",10339 => "11000011",10340 => "11011010",10341 => "00000011",10342 => "01110110",10343 => "11011001",10344 => "00010110",10345 => "01100010",10346 => "10010001",10347 => "10010101",10348 => "11011010",10349 => "01001000",10350 => "10001001",10351 => "01000011",10352 => "11100011",10353 => "10010110",10354 => "00110011",10355 => "10000000",10356 => "10101001",10357 => "11100011",10358 => "11001011",10359 => "00100010",10360 => "01000000",10361 => "10111001",10362 => "00001110",10363 => "01111100",10364 => "00100110",10365 => "00111000",10366 => "00001001",10367 => "01100110",10368 => "10000100",10369 => "11110011",10370 => "00100101",10371 => "11110001",10372 => "00010100",10373 => "01011011",10374 => "10110001",10375 => "00101101",10376 => "11111010",10377 => "01011100",10378 => "01010000",10379 => "00111010",10380 => "11110000",10381 => "00011110",10382 => "01101011",10383 => "01011010",10384 => "11010110",10385 => "10110100",10386 => "01000010",10387 => "10010001",10388 => "00001111",10389 => "10100100",10390 => "00001110",10391 => "00011111",10392 => "01000011",10393 => "01000100",10394 => "00111001",10395 => "00101101",10396 => "11000101",10397 => "01011001",10398 => "10101100",10399 => "00010110",10400 => "00000010",10401 => "11011110",10402 => "10000110",10403 => "00010111",10404 => "11100100",10405 => "10000110",10406 => "10001111",10407 => "11110011",10408 => "00100000",10409 => "10011001",10410 => "01000000",10411 => "01101101",10412 => "01110111",10413 => "10111110",10414 => "11110110",10415 => "01111101",10416 => "01111000",10417 => "00110001",10418 => "11101000",10419 => "10011010",10420 => "01110000",10421 => "01100101",10422 => "01011100",10423 => "00000000",10424 => "11110000",10425 => "01101111",10426 => "11100001",10427 => "11001111",10428 => "00010000",10429 => "10001110",10430 => "11010110",10431 => "11000001",10432 => "10001110",10433 => "11000100",10434 => "10100110",10435 => "01100011",10436 => "10010101",10437 => "00111110",10438 => "00001101",10439 => "11101111",10440 => "01010000",10441 => "00111110",10442 => "10110101",10443 => "01000110",10444 => "11101111",10445 => "10110000",10446 => "01010000",10447 => "10001110",10448 => "10001101",10449 => "10000001",10450 => "11111001",10451 => "01001001",10452 => "01100000",10453 => "00001100",10454 => "11100011",10455 => "00000001",10456 => "10011101",10457 => "00110001",10458 => "00111001",10459 => "10000111",10460 => "01111001",10461 => "11000000",10462 => "00111010",10463 => "00010000",10464 => "10100110",10465 => "10001010",10466 => "11001001",10467 => "10100000",10468 => "10101011",10469 => "11101101",10470 => "01000100",10471 => "01111100",10472 => "10011100",10473 => "11101001",10474 => "00111011",10475 => "01011100",10476 => "01101100",10477 => "00001111",10478 => "01110011",10479 => "11111111",10480 => "10000110",10481 => "00000111",10482 => "00011010",10483 => "00110011",10484 => "00100000",10485 => "00001001",10486 => "00101011",10487 => "10010001",10488 => "10110010",10489 => "10110101",10490 => "10101100",10491 => "11011011",10492 => "10110011",10493 => "11111011",10494 => "01101111",10495 => "01101100",10496 => "10111100",10497 => "10010001",10498 => "10011010",10499 => "11010000",10500 => "10011101",10501 => "11111101",10502 => "11100001",10503 => "10101010",10504 => "11101111",10505 => "01001100",10506 => "00111000",10507 => "00000010",10508 => "10101100",10509 => "10111000",10510 => "01101111",10511 => "11010101",10512 => "10001000",10513 => "10000100",10514 => "01011101",10515 => "10010001",10516 => "10011011",10517 => "01111110",10518 => "01011100",10519 => "01100100",10520 => "00110011",10521 => "01010111",10522 => "11000001",10523 => "00111110",10524 => "10111000",10525 => "00111011",10526 => "01010010",10527 => "00110001",10528 => "11110100",10529 => "01011010",10530 => "00111111",10531 => "10001011",10532 => "00000100",10533 => "01111000",10534 => "01111101",10535 => "11000100",10536 => "10010011",10537 => "01111111",10538 => "10110110",10539 => "10011110",10540 => "00010011",10541 => "00010011",10542 => "10111010",10543 => "00000100",10544 => "11101111",10545 => "01011001",10546 => "11111000",10547 => "10011111",10548 => "10000110",10549 => "00100010",10550 => "01000110",10551 => "10111101",10552 => "11001111",10553 => "10100110",10554 => "01011010",10555 => "01110001",10556 => "01000100",10557 => "00010100",10558 => "10110100",10559 => "01101001",10560 => "01110101",10561 => "00101001",10562 => "10110111",10563 => "01110010",10564 => "11001011",10565 => "10001011",10566 => "10110111",10567 => "00001100",10568 => "11010011",10569 => "01001111",10570 => "00111001",10571 => "01010010",10572 => "11110101",10573 => "00000101",10574 => "00110110",10575 => "01110010",10576 => "10010010",10577 => "01010011",10578 => "00110001",10579 => "10110101",10580 => "00011011",10581 => "11111010",10582 => "00001101",10583 => "11101000",10584 => "01001001",10585 => "10101111",10586 => "01010110",10587 => "11100001",10588 => "11000111",10589 => "10000010",10590 => "10101100",10591 => "00000100",10592 => "01100001",10593 => "00010111",10594 => "01010011",10595 => "01100110",10596 => "10001001",10597 => "01111011",10598 => "11011000",10599 => "10000000",10600 => "01100011",10601 => "11011110",10602 => "00110010",10603 => "10100011",10604 => "00101000",10605 => "11101111",10606 => "01110000",10607 => "11011011",10608 => "00000111",10609 => "00001101",10610 => "00111111",10611 => "00000110",10612 => "00101011",10613 => "00101011",10614 => "11110001",10615 => "11000010",10616 => "01110010",10617 => "11100111",10618 => "10111101",10619 => "00001010",10620 => "10000000",10621 => "01011010",10622 => "10111001",10623 => "01100000",10624 => "10011000",10625 => "11110011",10626 => "10110110",10627 => "00101010",10628 => "00101111",10629 => "10101000",10630 => "01000001",10631 => "10101010",10632 => "01000010",10633 => "11101101",10634 => "10010010",10635 => "11011111",10636 => "01001011",10637 => "01110101",10638 => "00001101",10639 => "00011110",10640 => "01000101",10641 => "01100101",10642 => "11110000",10643 => "00100101",10644 => "00011101",10645 => "01110100",10646 => "10000000",10647 => "00111111",10648 => "10110010",10649 => "00100011",10650 => "01011111",10651 => "01010010",10652 => "11100100",10653 => "10101010",10654 => "01101010",10655 => "10101000",10656 => "01101101",10657 => "01000110",10658 => "01111110",10659 => "11110100",10660 => "00001110",10661 => "00110101",10662 => "01110000",10663 => "11011101",10664 => "01101101",10665 => "00111001",10666 => "00000011",10667 => "01100101",10668 => "11000000",10669 => "10000100",10670 => "11100111",10671 => "11011100",10672 => "00101010",10673 => "01111001",10674 => "00111110",10675 => "11111110",10676 => "01110011",10677 => "01000100",10678 => "01011011",10679 => "10000101",10680 => "01001000",10681 => "10001111",10682 => "11111010",10683 => "10011100",10684 => "10000111",10685 => "11011010",10686 => "11100001",10687 => "11100111",10688 => "10010111",10689 => "01001010",10690 => "11100000",10691 => "10101111",10692 => "01100000",10693 => "01110101",10694 => "11011110",10695 => "10000110",10696 => "01101100",10697 => "01001011",10698 => "11111100",10699 => "10100001",10700 => "10001101",10701 => "00001011",10702 => "01001010",10703 => "01001100",10704 => "01010111",10705 => "00000000",10706 => "00100110",10707 => "11000010",10708 => "00100000",10709 => "00110000",10710 => "10111101",10711 => "01000111",10712 => "11000111",10713 => "01110001",10714 => "01101101",10715 => "10000001",10716 => "00101100",10717 => "01111011",10718 => "10110110",10719 => "10011111",10720 => "00110010",10721 => "00110011",10722 => "01100100",10723 => "00000000",10724 => "00111000",10725 => "01000011",10726 => "11101000",10727 => "00110110",10728 => "10001000",10729 => "01000010",10730 => "00110011",10731 => "10101110",10732 => "10010110",10733 => "10111110",10734 => "00100001",10735 => "11110001",10736 => "01000010",10737 => "11101101",10738 => "01111101",10739 => "00011110",10740 => "00011100",10741 => "01100100",10742 => "00100101",10743 => "00000100",10744 => "10100010",10745 => "01111101",10746 => "00101111",10747 => "01011110",10748 => "00101110",10749 => "10100111",10750 => "10100011",10751 => "00111100",10752 => "10101101",10753 => "10111011",10754 => "00110101",10755 => "00000000",10756 => "11000100",10757 => "01000000",10758 => "10011110",10759 => "01101010",10760 => "11011001",10761 => "11001000",10762 => "10111101",10763 => "11001110",10764 => "11101010",10765 => "01010100",10766 => "11111111",10767 => "11010100",10768 => "00000000",10769 => "00000110",10770 => "01101110",10771 => "11101011",10772 => "11101000",10773 => "10101000",10774 => "00001100",10775 => "01010000",10776 => "01010011",10777 => "10000000",10778 => "01110010",10779 => "00000001",10780 => "10001000",10781 => "01001001",10782 => "10101000",10783 => "01001010",10784 => "00100010",10785 => "10001110",10786 => "10011001",10787 => "10101010",10788 => "00000111",10789 => "01001001",10790 => "00011100",10791 => "11111110",10792 => "11111000",10793 => "00100011",10794 => "00000101",10795 => "00111011",10796 => "00100010",10797 => "11011110",10798 => "10001011",10799 => "01001111",10800 => "01011100",10801 => "10101010",10802 => "10010111",10803 => "10001100",10804 => "01111001",10805 => "10010001",10806 => "11010100",10807 => "10100000",10808 => "00000010",10809 => "01011100",10810 => "10110000",10811 => "10001110",10812 => "00111101",10813 => "10110110",10814 => "00011100",10815 => "10000100",10816 => "10111111",10817 => "00101000",10818 => "01011110",10819 => "00001111",10820 => "00011110",10821 => "01000000",10822 => "01101100",10823 => "01111100",10824 => "11111101",10825 => "01111100",10826 => "01111011",10827 => "10010100",10828 => "01000010",10829 => "00010111",10830 => "10000110",10831 => "11000111",10832 => "00100000",10833 => "10000010",10834 => "01010101",10835 => "11010001",10836 => "10101100",10837 => "01100100",10838 => "01001110",10839 => "10010101",10840 => "01001011",10841 => "00000111",10842 => "01000011",10843 => "01011010",10844 => "00010101",10845 => "11011110",10846 => "11001000",10847 => "01111101",10848 => "00001110",10849 => "10101111",10850 => "00111000",10851 => "10100100",10852 => "01101011",10853 => "01111011",10854 => "00001101",10855 => "01111001",10856 => "10001001",10857 => "00110100",10858 => "00100000",10859 => "10010011",10860 => "11100110",10861 => "01011000",10862 => "01100001",10863 => "11100110",10864 => "01110100",10865 => "10011110",10866 => "01000100",10867 => "10110000",10868 => "01101011",10869 => "10010011",10870 => "00111101",10871 => "01000011",10872 => "00001110",10873 => "01011011",10874 => "11111010",10875 => "01111110",10876 => "01101100",10877 => "01000011",10878 => "10001011",10879 => "01110001",10880 => "10000111",10881 => "01001010",10882 => "11001001",10883 => "01011001",10884 => "10001000",10885 => "00011111",10886 => "10000111",10887 => "11100101",10888 => "01011111",10889 => "01101000",10890 => "10101110",10891 => "10110101",10892 => "00100000",10893 => "10110100",10894 => "11011101",10895 => "11000000",10896 => "01011110",10897 => "00001110",10898 => "10001100",10899 => "00101011",10900 => "11111010",10901 => "01101101",10902 => "10001101",10903 => "00100001",10904 => "10000100",10905 => "11110101",10906 => "10001010",10907 => "01111110",10908 => "01000101",10909 => "01100010",10910 => "01000111",10911 => "10111011",10912 => "01011101",10913 => "11101110",10914 => "00111100",10915 => "11110101",10916 => "01000011",10917 => "10110110",10918 => "00001110",10919 => "11110001",10920 => "11101110",10921 => "00010011",10922 => "10010001",10923 => "01111111",10924 => "01001011",10925 => "00011110",10926 => "11101001",10927 => "10101011",10928 => "00101010",10929 => "00010110",10930 => "01111100",10931 => "01111001",10932 => "10110110",10933 => "00000010",10934 => "10000100",10935 => "01010000",10936 => "00111100",10937 => "11011010",10938 => "01110100",10939 => "01010111",10940 => "10000011",10941 => "01101011",10942 => "11100111",10943 => "00011111",10944 => "01011100",10945 => "00000011",10946 => "11000001",10947 => "10101001",10948 => "01001100",10949 => "01111000",10950 => "11100100",10951 => "01110111",10952 => "11001111",10953 => "10011001",10954 => "10010010",10955 => "10100101",10956 => "01001110",10957 => "00001001",10958 => "11010001",10959 => "10100001",10960 => "11100010",10961 => "11001111",10962 => "11011100",10963 => "00101011",10964 => "01110000",10965 => "10101011",10966 => "00001110",10967 => "01101001",10968 => "01110011",10969 => "11000010",10970 => "00110010",10971 => "01001100",10972 => "01111000",10973 => "01100100",10974 => "10100010",10975 => "00010100",10976 => "01000001",10977 => "01100111",10978 => "01101111",10979 => "00010101",10980 => "01101011",10981 => "00011100",10982 => "00111100",10983 => "01101001",10984 => "01001010",10985 => "00110001",10986 => "00100001",10987 => "11100010",10988 => "10110110",10989 => "10100011",10990 => "11111101",10991 => "00010010",10992 => "01001111",10993 => "11010010",10994 => "11110010",10995 => "10000110",10996 => "00011110",10997 => "00111110",10998 => "00011011",10999 => "01111001",11000 => "10111100",11001 => "01011110",11002 => "00110000",11003 => "11100111",11004 => "00001000",11005 => "01011001",11006 => "00000100",11007 => "11011100",11008 => "11111000",11009 => "11111000",11010 => "10110101",11011 => "10111110",11012 => "00101111",11013 => "10010101",11014 => "01110111",11015 => "00010010",11016 => "10100001",11017 => "00101111",11018 => "00010000",11019 => "01100111",11020 => "10100111",11021 => "00101100",11022 => "10011000",11023 => "00011010",11024 => "01010010",11025 => "11011100",11026 => "11111010",11027 => "11110111",11028 => "11110101",11029 => "11001101",11030 => "10111010",11031 => "11111000",11032 => "10111111",11033 => "10101110",11034 => "01101100",11035 => "01010111",11036 => "10111101",11037 => "11101100",11038 => "10111010",11039 => "10100000",11040 => "00101100",11041 => "11101000",11042 => "10110100",11043 => "01001011",11044 => "10010111",11045 => "00000001",11046 => "00110101",11047 => "01001111",11048 => "11001111",11049 => "10101011",11050 => "00011101",11051 => "01101101",11052 => "11011001",11053 => "00011111",11054 => "00100110",11055 => "01100010",11056 => "01010110",11057 => "01001010",11058 => "01001111",11059 => "01110101",11060 => "01011111",11061 => "10010010",11062 => "11011001",11063 => "01101010",11064 => "10110011",11065 => "10010110",11066 => "01000110",11067 => "11111010",11068 => "11000011",11069 => "01001000",11070 => "10110001",11071 => "11110100",11072 => "11110111",11073 => "11100001",11074 => "00110101",11075 => "00111000",11076 => "00000111",11077 => "00100110",11078 => "11101110",11079 => "11010000",11080 => "01000100",11081 => "01011000",11082 => "10011100",11083 => "01010001",11084 => "11011100",11085 => "01001101",11086 => "10011000",11087 => "00010011",11088 => "00100111",11089 => "10101110",11090 => "11011111",11091 => "00010000",11092 => "10101001",11093 => "10010110",11094 => "01111101",11095 => "01100100",11096 => "00001101",11097 => "11010110",11098 => "00111001",11099 => "10011011",11100 => "10011111",11101 => "00111111",11102 => "00101111",11103 => "01010100",11104 => "11000001",11105 => "01110010",11106 => "10111010",11107 => "10100001",11108 => "10111100",11109 => "10100000",11110 => "10111011",11111 => "10100010",11112 => "10110010",11113 => "11010100",11114 => "01010111",11115 => "01110001",11116 => "10010111",11117 => "01111110",11118 => "10010001",11119 => "01000111",11120 => "01011100",11121 => "00101001",11122 => "11110011",11123 => "11011110",11124 => "00110100",11125 => "11101100",11126 => "10010101",11127 => "01110001",11128 => "11001110",11129 => "11100000",11130 => "01111100",11131 => "00100110",11132 => "11110001",11133 => "11101110",11134 => "11000110",11135 => "00100110",11136 => "01010010",11137 => "01010100",11138 => "10001001",11139 => "00110010",11140 => "10000010",11141 => "01111111",11142 => "11000111",11143 => "00011000",11144 => "01011001",11145 => "01101010",11146 => "00111111",11147 => "10111011",11148 => "11101111",11149 => "00100001",11150 => "01111111",11151 => "10001011",11152 => "10101110",11153 => "00010011",11154 => "11110011",11155 => "00011100",11156 => "11111010",11157 => "01001010",11158 => "00101100",11159 => "10101100",11160 => "00110000",11161 => "01010001",11162 => "01011010",11163 => "10001110",11164 => "00010101",11165 => "10011100",11166 => "10001001",11167 => "11100010",11168 => "11010110",11169 => "00000111",11170 => "01010110",11171 => "10101011",11172 => "11100111",11173 => "11001110",11174 => "10111011",11175 => "11110001",11176 => "10011001",11177 => "10110001",11178 => "10000010",11179 => "11010000",11180 => "00110101",11181 => "00001001",11182 => "10000000",11183 => "00101011",11184 => "01101110",11185 => "01110001",11186 => "01111100",11187 => "01101100",11188 => "01010110",11189 => "00010100",11190 => "10100000",11191 => "01011010",11192 => "10101000",11193 => "00001111",11194 => "00010010",11195 => "00100011",11196 => "11110111",11197 => "00111100",11198 => "01001011",11199 => "00111001",11200 => "10101010",11201 => "10101101",11202 => "10100000",11203 => "01100100",11204 => "10011001",11205 => "10010000",11206 => "01010100",11207 => "11011000",11208 => "00010100",11209 => "11001111",11210 => "11110011",11211 => "11010011",11212 => "00001100",11213 => "11010010",11214 => "10100111",11215 => "11100001",11216 => "00011101",11217 => "00010000",11218 => "00111001",11219 => "01001000",11220 => "11100110",11221 => "01111111",11222 => "01001010",11223 => "11111101",11224 => "01001101",11225 => "00100100",11226 => "00110001",11227 => "01010011",11228 => "01100011",11229 => "01101010",11230 => "10010001",11231 => "11000111",11232 => "01011011",11233 => "00101011",11234 => "10100010",11235 => "10011110",11236 => "01010011",11237 => "00111100",11238 => "00101011",11239 => "01101110",11240 => "01111001",11241 => "10100110",11242 => "00000000",11243 => "11000110",11244 => "10011000",11245 => "01000100",11246 => "01010101",11247 => "11000010",11248 => "10110011",11249 => "00000001",11250 => "10100001",11251 => "00101111",11252 => "11010100",11253 => "10010001",11254 => "10011001",11255 => "01010000",11256 => "10111110",11257 => "10111001",11258 => "01011111",11259 => "11111100",11260 => "11110001",11261 => "10100000",11262 => "11111100",11263 => "11000111",11264 => "01011101",11265 => "00110101",11266 => "11110010",11267 => "10100111",11268 => "11101000",11269 => "11001101",11270 => "11100011",11271 => "10001111",11272 => "01001010",11273 => "10001001",11274 => "10111111",11275 => "01000001",11276 => "00010111",11277 => "01100001",11278 => "00011011",11279 => "00011000",11280 => "01100111",11281 => "10100001",11282 => "11001011",11283 => "01101001",11284 => "10001110",11285 => "11111011",11286 => "01001110",11287 => "10101110",11288 => "11101001",11289 => "10110001",11290 => "11011101",11291 => "10111011",11292 => "10001101",11293 => "00001101",11294 => "11111011",11295 => "10100101",11296 => "10111110",11297 => "00111111",11298 => "10101101",11299 => "10110010",11300 => "00001100",11301 => "01000001",11302 => "11001110",11303 => "10110110",11304 => "10001111",11305 => "11111111",11306 => "11000100",11307 => "00110101",11308 => "10011011",11309 => "11100100",11310 => "11000101",11311 => "00001000",11312 => "00110101",11313 => "10111111",11314 => "01010000",11315 => "11011101",11316 => "11001001",11317 => "11101110",11318 => "11101010",11319 => "01100001",11320 => "10011000",11321 => "11110110",11322 => "11100010",11323 => "00011100",11324 => "10011101",11325 => "01001111",11326 => "00001011",11327 => "00011101",11328 => "10100000",11329 => "11001111",11330 => "10011111",11331 => "01101101",11332 => "10011111",11333 => "01001001",11334 => "11001110",11335 => "00000101",11336 => "01111100",11337 => "00111110",11338 => "01110010",11339 => "01111010",11340 => "10010001",11341 => "01011010",11342 => "01011110",11343 => "01111001",11344 => "11111100",11345 => "11000101",11346 => "11100001",11347 => "10111111",11348 => "00101100",11349 => "11100000",11350 => "01010001",11351 => "01100011",11352 => "00011010",11353 => "11100100",11354 => "10011110",11355 => "10001100",11356 => "00001110",11357 => "10000100",11358 => "01011100",11359 => "00110101",11360 => "00000111",11361 => "01001111",11362 => "11110010",11363 => "11001110",11364 => "10111100",11365 => "10110011",11366 => "01010011",11367 => "01010101",11368 => "10111011",11369 => "01100010",11370 => "01100101",11371 => "01011101",11372 => "01000010",11373 => "00101010",11374 => "10101100",11375 => "01101100",11376 => "10100110",11377 => "11110100",11378 => "11110011",11379 => "00110011",11380 => "11111000",11381 => "11000110",11382 => "11001001",11383 => "00101000",11384 => "11001110",11385 => "11111101",11386 => "00000100",11387 => "00100100",11388 => "11011000",11389 => "10011101",11390 => "10100000",11391 => "11100010",11392 => "01110000",11393 => "00100111",11394 => "01100111",11395 => "11101100",11396 => "10101010",11397 => "10111100",11398 => "00000101",11399 => "11011010",11400 => "00001000",11401 => "01001111",11402 => "10100000",11403 => "01010111",11404 => "01110010",11405 => "10110001",11406 => "01110000",11407 => "10110111",11408 => "01010100",11409 => "01000110",11410 => "00000011",11411 => "11001111",11412 => "01111011",11413 => "01101111",11414 => "00110011",11415 => "01000111",11416 => "11101011",11417 => "11010110",11418 => "00000110",11419 => "01011011",11420 => "11100011",11421 => "01000011",11422 => "11111100",11423 => "01100000",11424 => "00111000",11425 => "11001001",11426 => "11011101",11427 => "00000010",11428 => "01001101",11429 => "00101101",11430 => "10001111",11431 => "10011011",11432 => "11101110",11433 => "01100011",11434 => "01111100",11435 => "11111000",11436 => "11010001",11437 => "11110111",11438 => "10010110",11439 => "10011111",11440 => "01001111",11441 => "00011010",11442 => "11010000",11443 => "10110111",11444 => "01011010",11445 => "01001101",11446 => "11010010",11447 => "00111111",11448 => "01011101",11449 => "11101010",11450 => "01111010",11451 => "01100110",11452 => "00000100",11453 => "10001011",11454 => "01011010",11455 => "11001011",11456 => "11101000",11457 => "11010010",11458 => "00001000",11459 => "10101010",11460 => "10110010",11461 => "11100000",11462 => "00000011",11463 => "11001001",11464 => "00110111",11465 => "10111111",11466 => "00001110",11467 => "11110011",11468 => "01111010",11469 => "00110100",11470 => "00111011",11471 => "10111101",11472 => "00111101",11473 => "10100011",11474 => "11010100",11475 => "00010100",11476 => "01000010",11477 => "00101011",11478 => "11010100",11479 => "11110100",11480 => "11000100",11481 => "00111110",11482 => "10001100",11483 => "10011011",11484 => "10101001",11485 => "01011111",11486 => "11111011",11487 => "01001111",11488 => "00101001",11489 => "10011100",11490 => "00001101",11491 => "10110111",11492 => "11110110",11493 => "11111101",11494 => "10000101",11495 => "11100011",11496 => "00101011",11497 => "00110111",11498 => "11000001",11499 => "00101011",11500 => "11000101",11501 => "11011010",11502 => "01001000",11503 => "01100111",11504 => "11101110",11505 => "00110011",11506 => "00000001",11507 => "00100001",11508 => "10110011",11509 => "11110000",11510 => "10001001",11511 => "01000100",11512 => "00010110",11513 => "01011100",11514 => "11111001",11515 => "10011000",11516 => "10100100",11517 => "10000011",11518 => "01011011",11519 => "00100000",11520 => "11110110",11521 => "10001001",11522 => "01010110",11523 => "01001101",11524 => "00110001",11525 => "11000000",11526 => "11111010",11527 => "10111001",11528 => "01111000",11529 => "11100111",11530 => "11011000",11531 => "00101111",11532 => "10100110",11533 => "01101000",11534 => "10011101",11535 => "00111110",11536 => "01110000",11537 => "11000101",11538 => "11111011",11539 => "01110000",11540 => "01110101",11541 => "10101111",11542 => "10010010",11543 => "00000100",11544 => "00110101",11545 => "10111010",11546 => "10111110",11547 => "11110110",11548 => "11000001",11549 => "01000000",11550 => "10100100",11551 => "01011101",11552 => "11000101",11553 => "10010100",11554 => "00100111",11555 => "00111000",11556 => "11001001",11557 => "00000111",11558 => "11011100",11559 => "00011001",11560 => "01010000",11561 => "10110100",11562 => "00110010",11563 => "10101010",11564 => "01111011",11565 => "10010010",11566 => "01000101",11567 => "01101001",11568 => "01010001",11569 => "11111011",11570 => "11101101",11571 => "00100011",11572 => "00001000",11573 => "00011000",11574 => "01011100",11575 => "01010001",11576 => "10011110",11577 => "11011110",11578 => "01001011",11579 => "00011101",11580 => "01101101",11581 => "10101111",11582 => "11111000",11583 => "10011011",11584 => "11101101",11585 => "01010001",11586 => "00011111",11587 => "00010111",11588 => "10000111",11589 => "11111101",11590 => "01110001",11591 => "11010000",11592 => "11000111",11593 => "10010010",11594 => "10000001",11595 => "11001100",11596 => "10001111",11597 => "11100011",11598 => "01110001",11599 => "10110110",11600 => "00000101",11601 => "11111011",11602 => "01010011",11603 => "11000000",11604 => "10010111",11605 => "01111110",11606 => "11111111",11607 => "00001100",11608 => "00001111",11609 => "10011110",11610 => "10100100",11611 => "10000101",11612 => "00100110",11613 => "10111011",11614 => "00011111",11615 => "00001100",11616 => "01110101",11617 => "11010010",11618 => "10110001",11619 => "01110110",11620 => "11000111",11621 => "00011111",11622 => "00101110",11623 => "10101101",11624 => "00011001",11625 => "01100100",11626 => "11011101",11627 => "11111100",11628 => "00111100",11629 => "00011111",11630 => "01011010",11631 => "00011101",11632 => "01000100",11633 => "11011110",11634 => "11010010",11635 => "00111010",11636 => "00000101",11637 => "11110111",11638 => "11001111",11639 => "00011101",11640 => "00100100",11641 => "10110010",11642 => "11111100",11643 => "01000001",11644 => "11010001",11645 => "00010111",11646 => "10100011",11647 => "10100011",11648 => "11001111",11649 => "00110110",11650 => "01100001",11651 => "01100101",11652 => "01010100",11653 => "10100000",11654 => "11010011",11655 => "01111101",11656 => "11000111",11657 => "01011101",11658 => "11101111",11659 => "11111100",11660 => "11110110",11661 => "00101000",11662 => "10100101",11663 => "00000100",11664 => "00101011",11665 => "01001101",11666 => "01111110",11667 => "10101000",11668 => "10010001",11669 => "11101011",11670 => "01010001",11671 => "01101000",11672 => "11011001",11673 => "01010100",11674 => "00111100",11675 => "01110011",11676 => "00101101",11677 => "10101101",11678 => "10011000",11679 => "11010110",11680 => "11010101",11681 => "01010011",11682 => "11101001",11683 => "00111010",11684 => "00111111",11685 => "01000100",11686 => "10010000",11687 => "01100100",11688 => "00100111",11689 => "11111001",11690 => "01111110",11691 => "00010111",11692 => "01000111",11693 => "01000001",11694 => "11010010",11695 => "00110001",11696 => "11000010",11697 => "00000110",11698 => "11010110",11699 => "10111110",11700 => "11100010",11701 => "10101101",11702 => "11110000",11703 => "11010001",11704 => "00011110",11705 => "10101111",11706 => "00100110",11707 => "00111100",11708 => "11000100",11709 => "01010111",11710 => "01100100",11711 => "01100101",11712 => "11100010",11713 => "00000100",11714 => "01110111",11715 => "11110100",11716 => "11011001",11717 => "01010011",11718 => "10001110",11719 => "00011010",11720 => "10000011",11721 => "11100010",11722 => "00101001",11723 => "11111100",11724 => "11100001",11725 => "11010011",11726 => "10110110",11727 => "00000010",11728 => "01100000",11729 => "11001000",11730 => "01001011",11731 => "10001101",11732 => "01010100",11733 => "01011010",11734 => "01011111",11735 => "00001111",11736 => "00110100",11737 => "10011101",11738 => "00110000",11739 => "00101010",11740 => "01001101",11741 => "11101100",11742 => "00110011",11743 => "01000001",11744 => "11110101",11745 => "00111011",11746 => "01001010",11747 => "11000100",11748 => "01000111",11749 => "10000101",11750 => "01110100",11751 => "01100111",11752 => "00110011",11753 => "10110101",11754 => "01110101",11755 => "11000001",11756 => "00011110",11757 => "00101000",11758 => "00010010",11759 => "11110011",11760 => "00011101",11761 => "01111011",11762 => "10010010",11763 => "11001000",11764 => "11110100",11765 => "11011111",11766 => "10100111",11767 => "10000110",11768 => "01111111",11769 => "11011101",11770 => "00000000",11771 => "01000001",11772 => "11000100",11773 => "11010110",11774 => "11011100",11775 => "00010010",11776 => "01000001",11777 => "11101101",11778 => "00010011",11779 => "11011001",11780 => "00110000",11781 => "10101111",11782 => "10110100",11783 => "11000011",11784 => "00101101",11785 => "00001010",11786 => "00000001",11787 => "01101010",11788 => "11000000",11789 => "00100011",11790 => "10111111",11791 => "11000010",11792 => "11110000",11793 => "01001010",11794 => "10101100",11795 => "11011110",11796 => "10110000",11797 => "11000110",11798 => "00111000",11799 => "10111100",11800 => "00100101",11801 => "11001010",11802 => "11010100",11803 => "01110001",11804 => "10000011",11805 => "10100001",11806 => "00111000",11807 => "00001100",11808 => "10000111",11809 => "01010111",11810 => "10001010",11811 => "10000011",11812 => "11111010",11813 => "01000010",11814 => "11011100",11815 => "01101101",11816 => "01111010",11817 => "10101001",11818 => "11110111",11819 => "00011110",11820 => "00100111",11821 => "11111011",11822 => "01001110",11823 => "01000110",11824 => "10111101",11825 => "10000010",11826 => "10111110",11827 => "10100011",11828 => "00010001",11829 => "11000111",11830 => "01000100",11831 => "00011001",11832 => "00110000",11833 => "11000111",11834 => "10000101",11835 => "11011110",11836 => "01010011",11837 => "11110000",11838 => "00001011",11839 => "01101010",11840 => "01000000",11841 => "01111100",11842 => "11100000",11843 => "00001000",11844 => "11011110",11845 => "01000000",11846 => "10000000",11847 => "01001111",11848 => "11110110",11849 => "10111001",11850 => "11110000",11851 => "00111010",11852 => "10100111",11853 => "00011101",11854 => "10110010",11855 => "00011100",11856 => "11010000",11857 => "10000110",11858 => "00001010",11859 => "01101111",11860 => "10100101",11861 => "11000011",11862 => "10110100",11863 => "11101011",11864 => "10110111",11865 => "01010101",11866 => "10110100",11867 => "10101100",11868 => "00011101",11869 => "11111101",11870 => "00011110",11871 => "11111010",11872 => "01011001",11873 => "01011100",11874 => "01111000",11875 => "00110011",11876 => "00100011",11877 => "00010010",11878 => "01101111",11879 => "10010110",11880 => "00010001",11881 => "01010001",11882 => "01010010",11883 => "11101000",11884 => "01000101",11885 => "10010010",11886 => "00000001",11887 => "00001011",11888 => "01010110",11889 => "10010101",11890 => "10101101",11891 => "11011011",11892 => "10111100",11893 => "10110101",11894 => "01111110",11895 => "01101011",11896 => "10010101",11897 => "00111000",11898 => "00010100",11899 => "10001000",11900 => "00000111",11901 => "11011111",11902 => "01000110",11903 => "11100001",11904 => "11010011",11905 => "00111111",11906 => "10000111",11907 => "00001111",11908 => "11111100",11909 => "11101100",11910 => "11011010",11911 => "00000101",11912 => "11100000",11913 => "11101110",11914 => "10011011",11915 => "00101100",11916 => "01000110",11917 => "10100010",11918 => "10100101",11919 => "00000110",11920 => "01100001",11921 => "00010101",11922 => "00000100",11923 => "00101000",11924 => "11000010",11925 => "00100011",11926 => "11101010",11927 => "11010010",11928 => "11110000",11929 => "10101100",11930 => "10011000",11931 => "11010011",11932 => "11001111",11933 => "11010100",11934 => "01001011",11935 => "10100100",11936 => "00001011",11937 => "01101011",11938 => "11100001",11939 => "00000010",11940 => "11111110",11941 => "01111010",11942 => "10000101",11943 => "00000001",11944 => "00100111",11945 => "10011010",11946 => "11001111",11947 => "11100011",11948 => "10000111",11949 => "01100001",11950 => "11110010",11951 => "00001001",11952 => "11101100",11953 => "10111010",11954 => "00010001",11955 => "01011111",11956 => "11010001",11957 => "01101111",11958 => "11110100",11959 => "10000110",11960 => "00111000",11961 => "10000010",11962 => "10100100",11963 => "11100111",11964 => "00011110",11965 => "11011000",11966 => "01001110",11967 => "00111101",11968 => "00011010",11969 => "11001111",11970 => "11000011",11971 => "10101111",11972 => "00110100",11973 => "11010111",11974 => "10000011",11975 => "00010001",11976 => "11011010",11977 => "11001011",11978 => "00000100",11979 => "00110100",11980 => "01110110",11981 => "00110110",11982 => "11110000",11983 => "10010100",11984 => "01001010",11985 => "11111001",11986 => "11000000",11987 => "10100011",11988 => "10111100",11989 => "01101101",11990 => "11101100",11991 => "11001010",11992 => "01011110",11993 => "10101000",11994 => "10010100",11995 => "11010101",11996 => "01011011",11997 => "11110011",11998 => "10111111",11999 => "10101101",12000 => "01011001",12001 => "00110011",12002 => "10110010",12003 => "11010110",12004 => "01010011",12005 => "00000101",12006 => "10000110",12007 => "01111110",12008 => "11001111",12009 => "01100011",12010 => "00000101",12011 => "10001110",12012 => "00100100",12013 => "00111110",12014 => "10110101",12015 => "01100011",12016 => "11111110",12017 => "11000011",12018 => "01111101",12019 => "00000010",12020 => "11110011",12021 => "11011101",12022 => "00110000",12023 => "10010001",12024 => "11001111",12025 => "00001111",12026 => "01111101",12027 => "11000111",12028 => "10100110",12029 => "11000110",12030 => "00011000",12031 => "01000010",12032 => "01111111",12033 => "10101101",12034 => "01100100",12035 => "10100110",12036 => "00011110",12037 => "00010100",12038 => "11100010",12039 => "11010110",12040 => "10101101",12041 => "10001011",12042 => "00101011",12043 => "01000001",12044 => "01000100",12045 => "10011101",12046 => "01000000",12047 => "01101110",12048 => "10011011",12049 => "10001011",12050 => "11000011",12051 => "11101000",12052 => "10100101",12053 => "00100010",12054 => "00110110",12055 => "01100010",12056 => "00001010",12057 => "10011010",12058 => "10111111",12059 => "11110000",12060 => "00110101",12061 => "11001011",12062 => "10011110",12063 => "10100101",12064 => "01110010",12065 => "00000000",12066 => "00011100",12067 => "00110001",12068 => "11000101",12069 => "01111000",12070 => "11110111",12071 => "01110111",12072 => "10100001",12073 => "10000010",12074 => "11110101",12075 => "01010101",12076 => "10110111",12077 => "01100001",12078 => "11000111",12079 => "01011010",12080 => "10101011",12081 => "10100110",12082 => "00011011",12083 => "01001011",12084 => "01001011",12085 => "01010110",12086 => "01101110",12087 => "11111110",12088 => "00100110",12089 => "01001010",12090 => "00000101",12091 => "11110010",12092 => "11111101",12093 => "00101100",12094 => "10010010",12095 => "01110010",12096 => "11000110",12097 => "10001011",12098 => "00110110",12099 => "11101111",12100 => "01101111",12101 => "11100011",12102 => "10110101",12103 => "11101111",12104 => "01010111",12105 => "11010111",12106 => "10101100",12107 => "00000000",12108 => "10000111",12109 => "11000101",12110 => "10001010",12111 => "10111101",12112 => "00010111",12113 => "01000001",12114 => "11100101",12115 => "10010001",12116 => "10011110",12117 => "00001011",12118 => "10111110",12119 => "10010011",12120 => "01000101",12121 => "00100011",12122 => "11010010",12123 => "11010000",12124 => "00011000",12125 => "00100011",12126 => "10010010",12127 => "00111000",12128 => "11011101",12129 => "10101011",12130 => "01111110",12131 => "10011000",12132 => "00011001",12133 => "11011000",12134 => "11100011",12135 => "11110101",12136 => "11111111",12137 => "00011100",12138 => "10000010",12139 => "00111011",12140 => "00101001",12141 => "00011101",12142 => "10010101",12143 => "10001001",12144 => "00111010",12145 => "00111001",12146 => "11101101",12147 => "01111000",12148 => "01001001",12149 => "11000100",12150 => "01101010",12151 => "00100110",12152 => "11000110",12153 => "10101000",12154 => "11110100",12155 => "10110110",12156 => "01110100",12157 => "01101100",12158 => "11011100",12159 => "01010010",12160 => "00110000",12161 => "11101111",12162 => "11110101",12163 => "11110010",12164 => "10000001",12165 => "00010010",12166 => "00001001",12167 => "01110100",12168 => "10101000",12169 => "01110111",12170 => "11011011",12171 => "00111010",12172 => "01010111",12173 => "01010010",12174 => "10100101",12175 => "10111110",12176 => "01110100",12177 => "10101100",12178 => "01010010",12179 => "11000001",12180 => "00000110",12181 => "00010000",12182 => "11101010",12183 => "00001100",12184 => "11011110",12185 => "10000010",12186 => "10110011",12187 => "00010110",12188 => "11000110",12189 => "01110000",12190 => "11111000",12191 => "01111010",12192 => "11011110",12193 => "10111010",12194 => "10100111",12195 => "01110101",12196 => "01101000",12197 => "00110001",12198 => "00001100",12199 => "01111111",12200 => "01001101",12201 => "11010001",12202 => "00100111",12203 => "00111110",12204 => "01000101",12205 => "11010101",12206 => "11001000",12207 => "11101111",12208 => "11010000",12209 => "11100000",12210 => "10101000",12211 => "10010001",12212 => "11110111",12213 => "00010010",12214 => "10001000",12215 => "10010100",12216 => "10100110",12217 => "01111100",12218 => "01011111",12219 => "11010000",12220 => "01110000",12221 => "11000010",12222 => "01110011",12223 => "01111100",12224 => "11101101",12225 => "00100111",12226 => "11111000",12227 => "10110000",12228 => "10001010",12229 => "10001100",12230 => "01100001",12231 => "01110010",12232 => "01011111",12233 => "10111001",12234 => "01111111",12235 => "10011010",12236 => "01100001",12237 => "11101100",12238 => "00000101",12239 => "10111010",12240 => "11111111",12241 => "10001011",12242 => "00110010",12243 => "00011100",12244 => "10110111",12245 => "11011111",12246 => "01011011",12247 => "01101000",12248 => "01111101",12249 => "10001111",12250 => "10111011",12251 => "11010100",12252 => "10110011",12253 => "00010111",12254 => "01110101",12255 => "10010101",12256 => "11101100",12257 => "11011011",12258 => "01100100",12259 => "10100010",12260 => "01111100",12261 => "10011001",12262 => "11101111",12263 => "00111001",12264 => "00100101",12265 => "00110101",12266 => "10010111",12267 => "11010010",12268 => "10001000",12269 => "10000101",12270 => "01011010",12271 => "10011101",12272 => "11010110",12273 => "00010011",12274 => "10110000",12275 => "10000110",12276 => "01100110",12277 => "00110111",12278 => "11000110",12279 => "10101111",12280 => "11011110",12281 => "00010010",12282 => "01110011",12283 => "11111101",12284 => "10100111",12285 => "00110000",12286 => "11111000",12287 => "11110010",12288 => "00100010",12289 => "01110000",12290 => "01101111",12291 => "01111000",12292 => "00101011",12293 => "10100111",12294 => "00010000",12295 => "00010001",12296 => "11101010",12297 => "11011111",12298 => "10000001",12299 => "01110011",12300 => "01110000",12301 => "11110011",12302 => "11110011",12303 => "10101001",12304 => "01101111",12305 => "10101011",12306 => "00001100",12307 => "01101010",12308 => "10000101",12309 => "11001011",12310 => "11000001",12311 => "11010100",12312 => "11111011",12313 => "01001110",12314 => "01110000",12315 => "01110011",12316 => "01001001",12317 => "00001000",12318 => "11010011",12319 => "10101101",12320 => "01101101",12321 => "01100011",12322 => "01010011",12323 => "11110001",12324 => "01101110",12325 => "11000010",12326 => "11000001",12327 => "11000110",12328 => "01110110",12329 => "11101100",12330 => "10011111",12331 => "00001100",12332 => "11110010",12333 => "10111011",12334 => "10111011",12335 => "01000101",12336 => "10011001",12337 => "11100000",12338 => "00011110",12339 => "10001111",12340 => "11100100",12341 => "00110000",12342 => "00010001",12343 => "11110010",12344 => "00000110",12345 => "10010101",12346 => "01010100",12347 => "01011111",12348 => "01101000",12349 => "11110111",12350 => "11100101",12351 => "01001011",12352 => "11000001",12353 => "11001000",12354 => "10110100",12355 => "10000100",12356 => "00101100",12357 => "01111101",12358 => "11111011",12359 => "10100100",12360 => "00000100",12361 => "01011010",12362 => "11110001",12363 => "00110101",12364 => "10000111",12365 => "10001000",12366 => "01010001",12367 => "10100000",12368 => "11100110",12369 => "00110110",12370 => "01110111",12371 => "00110000",12372 => "10101000",12373 => "11111011",12374 => "01110100",12375 => "11100101",12376 => "00010000",12377 => "11001000",12378 => "01110010",12379 => "01000011",12380 => "01100001",12381 => "01111011",12382 => "11011001",12383 => "01101111",12384 => "11001001",12385 => "11000001",12386 => "11010000",12387 => "00011010",12388 => "00101100",12389 => "00101100",12390 => "01111010",12391 => "11101110",12392 => "00101011",12393 => "11101010",12394 => "11011001",12395 => "10101111",12396 => "01110110",12397 => "00111010",12398 => "10001101",12399 => "00011011",12400 => "10111000",12401 => "00000111",12402 => "11001100",12403 => "11011011",12404 => "11000011",12405 => "10000111",12406 => "00111111",12407 => "00011110",12408 => "01011011",12409 => "00011111",12410 => "11111010",12411 => "11011001",12412 => "10001111",12413 => "01110101",12414 => "10111100",12415 => "00101101",12416 => "11100011",12417 => "11101011",12418 => "10010100",12419 => "00010110",12420 => "10000011",12421 => "11000101",12422 => "01110101",12423 => "11111110",12424 => "11010111",12425 => "11101001",12426 => "11010101",12427 => "10100101",12428 => "00101101",12429 => "10100001",12430 => "11111001",12431 => "11110110",12432 => "01010010",12433 => "01100000",12434 => "01011100",12435 => "00001110",12436 => "10011110",12437 => "00000000",12438 => "01101010",12439 => "01110000",12440 => "00010011",12441 => "00001101",12442 => "00001011",12443 => "10100010",12444 => "01111001",12445 => "10010100",12446 => "01110001",12447 => "01100001",12448 => "10110001",12449 => "00011011",12450 => "01011011",12451 => "01100000",12452 => "10100100",12453 => "10100000",12454 => "11000001",12455 => "11000100",12456 => "11111000",12457 => "10111110",12458 => "11101000",12459 => "00000010",12460 => "01110001",12461 => "00010010",12462 => "10001011",12463 => "01010110",12464 => "01011010",12465 => "00101111",12466 => "11001110",12467 => "00010010",12468 => "01111011",12469 => "10111011",12470 => "00100001",12471 => "01100000",12472 => "00011110",12473 => "11101011",12474 => "01001001",12475 => "11000110",12476 => "11001111",12477 => "01000010",12478 => "10000100",12479 => "00010011",12480 => "01100111",12481 => "01000001",12482 => "01100101",12483 => "01000111",12484 => "11110111",12485 => "00011100",12486 => "11100010",12487 => "11011000",12488 => "00010100",12489 => "11001001",12490 => "11111001",12491 => "00110001",12492 => "00010111",12493 => "11100101",12494 => "01101101",12495 => "00100001",12496 => "01011001",12497 => "10000100",12498 => "11110000",12499 => "10101111",12500 => "01010100",12501 => "01111000",12502 => "10001010",12503 => "00001110",12504 => "10000010",12505 => "01111000",12506 => "00110110",12507 => "10011111",12508 => "01100001",12509 => "01011110",12510 => "11000111",12511 => "00100000",12512 => "10100111",12513 => "10010001",12514 => "00001101",12515 => "11000010",12516 => "00111110",12517 => "01011010",12518 => "01111110",12519 => "11100101",12520 => "10110101",12521 => "00011110",12522 => "10101100",12523 => "01100101",12524 => "00000010",12525 => "11010000",12526 => "10101001",12527 => "10000000",12528 => "01101110",12529 => "10110110",12530 => "00000000",12531 => "11100000",12532 => "00111100",12533 => "00110111",12534 => "10010111",12535 => "01011100",12536 => "10001110",12537 => "00110110",12538 => "10001100",12539 => "00101100",12540 => "01110001",12541 => "10011011",12542 => "11110011",12543 => "10001111",12544 => "11011001",12545 => "00111010",12546 => "11000101",12547 => "00001101",12548 => "00000000",12549 => "10110111",12550 => "11010110",12551 => "10000011",12552 => "00000111",12553 => "11001101",12554 => "10011000",12555 => "11001000",12556 => "01111111",12557 => "01001010",12558 => "00111100",12559 => "00010111",12560 => "01101101",12561 => "10010001",12562 => "00000100",12563 => "11001111",12564 => "10111010",12565 => "11111010",12566 => "00000011",12567 => "01100011",12568 => "00010111",12569 => "00000110",12570 => "01010010",12571 => "11111110",12572 => "10110001",12573 => "01111010",12574 => "10111100",12575 => "01011011",12576 => "11011001",12577 => "10101010",12578 => "10010111",12579 => "00100101",12580 => "11001101",12581 => "01000011",12582 => "00010000",12583 => "11100101",12584 => "11010000",12585 => "10011001",12586 => "10011110",12587 => "11010010",12588 => "00111100",12589 => "10111110",12590 => "10001101",12591 => "00110101",12592 => "00100111",12593 => "11100110",12594 => "01011000",12595 => "01011110",12596 => "01111110",12597 => "00100011",12598 => "00110111",12599 => "01001111",12600 => "10111110",12601 => "11000001",12602 => "10001010",12603 => "11111101",12604 => "11001000",12605 => "11110010",12606 => "11000111",12607 => "01011001",12608 => "01000000",12609 => "10110010",12610 => "11010110",12611 => "01101110",12612 => "01111110",12613 => "00101101",12614 => "00000110",12615 => "01001110",12616 => "11101001",12617 => "01001110",12618 => "11011001",12619 => "10111110",12620 => "11111111",12621 => "00100011",12622 => "00101011",12623 => "10111010",12624 => "10001110",12625 => "10000110",12626 => "00110101",12627 => "00000101",12628 => "10111100",12629 => "10110010",12630 => "00011001",12631 => "00010100",12632 => "10000010",12633 => "01000110",12634 => "11100001",12635 => "00011010",12636 => "10101000",12637 => "01111110",12638 => "00001001",12639 => "11010001",12640 => "10111101",12641 => "00010111",12642 => "01010001",12643 => "10101001",12644 => "11001000",12645 => "00010100",12646 => "00100100",12647 => "10100010",12648 => "10011111",12649 => "10111100",12650 => "10001001",12651 => "10001110",12652 => "01101100",12653 => "11001001",12654 => "00101010",12655 => "01011011",12656 => "11111010",12657 => "10011101",12658 => "00111011",12659 => "10100011",12660 => "10011110",12661 => "00000011",12662 => "01110011",12663 => "00000110",12664 => "00001100",12665 => "01110001",12666 => "00000101",12667 => "11100011",12668 => "01111000",12669 => "10110101",12670 => "10111110",12671 => "10011011",12672 => "00010111",12673 => "10001100",12674 => "11010101",12675 => "01111101",12676 => "00000001",12677 => "10010111",12678 => "00001010",12679 => "10010001",12680 => "01101111",12681 => "10100100",12682 => "11011010",12683 => "11100110",12684 => "11001011",12685 => "00110101",12686 => "10000001",12687 => "10101110",12688 => "01010110",12689 => "01001110",12690 => "10010011",12691 => "00111100",12692 => "11000001",12693 => "11011011",12694 => "01010110",12695 => "01010100",12696 => "00001001",12697 => "00000001",12698 => "01100000",12699 => "10110101",12700 => "01001111",12701 => "01000100",12702 => "11001100",12703 => "01100001",12704 => "01000000",12705 => "11101011",12706 => "10100010",12707 => "01101100",12708 => "01001111",12709 => "11011101",12710 => "00100111",12711 => "00101000",12712 => "10100101",12713 => "10010111",12714 => "01000100",12715 => "01101011",12716 => "11000100",12717 => "10100111",12718 => "11001010",12719 => "10101001",12720 => "10101001",12721 => "10111110",12722 => "00111000",12723 => "00110110",12724 => "11001110",12725 => "10101110",12726 => "10001010",12727 => "11101111",12728 => "01100111",12729 => "01101100",12730 => "10010010",12731 => "11010001",12732 => "00111011",12733 => "01101100",12734 => "01110001",12735 => "11100001",12736 => "10110011",12737 => "10101111",12738 => "01010010",12739 => "11111110",12740 => "11010101",12741 => "11111010",12742 => "11110110",12743 => "11000010",12744 => "10110000",12745 => "10100100",12746 => "00000100",12747 => "10100010",12748 => "00111101",12749 => "10001101",12750 => "01010111",12751 => "01110001",12752 => "10111110",12753 => "10000011",12754 => "00000011",12755 => "01010101",12756 => "01010010",12757 => "00101110",12758 => "00010001",12759 => "01111000",12760 => "10010111",12761 => "10101110",12762 => "10100001",12763 => "00111011",12764 => "01001011",12765 => "01110111",12766 => "11010000",12767 => "11000111",12768 => "00111101",12769 => "01010100",12770 => "01100010",12771 => "00000110",12772 => "11010000",12773 => "01011010",12774 => "00001001",12775 => "11101010",12776 => "10100001",12777 => "00111001",12778 => "11100011",12779 => "00100101",12780 => "11011011",12781 => "11110101",12782 => "10110010",12783 => "00010001",12784 => "01000000",12785 => "00111111",12786 => "11111011",12787 => "01100010",12788 => "01110010",12789 => "11011001",12790 => "10001100",12791 => "01000101",12792 => "00111001",12793 => "01110000",12794 => "01110011",12795 => "11010000",12796 => "01011010",12797 => "01001010",12798 => "01111101",12799 => "01100001",12800 => "01011110",12801 => "11110000",12802 => "01101011",12803 => "11100100",12804 => "00011010",12805 => "11001000",12806 => "01101001",12807 => "11110100",12808 => "10110000",12809 => "00110101",12810 => "10000000",12811 => "01101000",12812 => "10010001",12813 => "10000110",12814 => "01101101",12815 => "00000111",12816 => "10001111",12817 => "00001000",12818 => "11101111",12819 => "11101101",12820 => "01010011",12821 => "11100001",12822 => "00000011",12823 => "00110101",12824 => "00010011",12825 => "01010110",12826 => "10001010",12827 => "00010001",12828 => "11101001",12829 => "01001010",12830 => "10010110",12831 => "10010011",12832 => "00001001",12833 => "00100010",12834 => "00111000",12835 => "00110101",12836 => "10010101",12837 => "10011001",12838 => "00100101",12839 => "00010010",12840 => "10100000",12841 => "11010111",12842 => "10001111",12843 => "10000111",12844 => "11011001",12845 => "01101101",12846 => "00111011",12847 => "11010000",12848 => "01111011",12849 => "00001110",12850 => "10011011",12851 => "10110100",12852 => "10101100",12853 => "10101001",12854 => "11010011",12855 => "10100010",12856 => "00010001",12857 => "11011000",12858 => "11111101",12859 => "01100010",12860 => "00110101",12861 => "11111010",12862 => "11110010",12863 => "11000011",12864 => "10101100",12865 => "11001100",12866 => "00010100",12867 => "01000101",12868 => "01001110",12869 => "01101010",12870 => "11100010",12871 => "00100001",12872 => "00111100",12873 => "01010011",12874 => "10100110",12875 => "00100010",12876 => "11100010",12877 => "10010101",12878 => "11110000",12879 => "00000011",12880 => "01111000",12881 => "01010011",12882 => "10010111",12883 => "00001010",12884 => "10110100",12885 => "10011011",12886 => "00110000",12887 => "11010111",12888 => "01011111",12889 => "11110001",12890 => "01011010",12891 => "01101010",12892 => "11010100",12893 => "01011100",12894 => "01111111",12895 => "00100010",12896 => "11110000",12897 => "01010101",12898 => "11000011",12899 => "01000011",12900 => "10010001",12901 => "10101110",12902 => "01001100",12903 => "10011111",12904 => "00001010",12905 => "00010010",12906 => "00010111",12907 => "10111011",12908 => "00111110",12909 => "11001010",12910 => "11110001",12911 => "11101101",12912 => "10111111",12913 => "11110001",12914 => "01000011",12915 => "11110010",12916 => "10010110",12917 => "00001100",12918 => "01001011",12919 => "00001010",12920 => "11000010",12921 => "11011100",12922 => "00010011",12923 => "01110011",12924 => "11110100",12925 => "01110111",12926 => "10100111",12927 => "10100100",12928 => "01100001",12929 => "00111111",12930 => "01001011",12931 => "10001010",12932 => "10110110",12933 => "00100100",12934 => "10100010",12935 => "10010110",12936 => "11111000",12937 => "10110110",12938 => "11100001",12939 => "00101011",12940 => "00101110",12941 => "11000111",12942 => "10111001",12943 => "01100000",12944 => "00011101",12945 => "01100011",12946 => "00100011",12947 => "00001000",12948 => "11101011",12949 => "10010100",12950 => "11100011",12951 => "11110011",12952 => "01111111",12953 => "01111001",12954 => "01100001",12955 => "01010111",12956 => "10000010",12957 => "00011111",12958 => "01000110",12959 => "01111100",12960 => "01110011",12961 => "10111101",12962 => "00000100",12963 => "11110001",12964 => "11110011",12965 => "01101101",12966 => "00100100",12967 => "01111010",12968 => "10111011",12969 => "10110010",12970 => "00001111",12971 => "00010000",12972 => "01000100",12973 => "10100000",12974 => "10111100",12975 => "00101101",12976 => "11100001",12977 => "01000001",12978 => "11110101",12979 => "11000100",12980 => "01110111",12981 => "11001001",12982 => "00000010",12983 => "00011111",12984 => "10100101",12985 => "00001000",12986 => "01001010",12987 => "11000001",12988 => "01101010",12989 => "11010010",12990 => "01001110",12991 => "10111101",12992 => "01110101",12993 => "00011001",12994 => "11001001",12995 => "00100010",12996 => "00011000",12997 => "11110110",12998 => "11010110",12999 => "00010110",13000 => "01000011",13001 => "01110101",13002 => "11001011",13003 => "00010001",13004 => "10110000",13005 => "00110101",13006 => "11110100",13007 => "10001001",13008 => "10011101",13009 => "00001100",13010 => "00101110",13011 => "11110000",13012 => "00111111",13013 => "11000100",13014 => "11010110",13015 => "00000110",13016 => "10011000",13017 => "11011000",13018 => "11111111",13019 => "00011010",13020 => "01100100",13021 => "10101110",13022 => "10100010",13023 => "10001111",13024 => "11100000",13025 => "00100101",13026 => "00100000",13027 => "01010100",13028 => "00101001",13029 => "00011110",13030 => "00111001",13031 => "11001000",13032 => "10111000",13033 => "00101010",13034 => "01000100",13035 => "00011111",13036 => "00111011",13037 => "01011010",13038 => "11111101",13039 => "00100010",13040 => "11111101",13041 => "01011000",13042 => "01011001",13043 => "01100001",13044 => "01000111",13045 => "00110110",13046 => "01000001",13047 => "10101011",13048 => "10001110",13049 => "10111100",13050 => "10110011",13051 => "11001110",13052 => "10000010",13053 => "01110000",13054 => "11010000",13055 => "00010100",13056 => "10111101",13057 => "00101100",13058 => "01011100",13059 => "11001100",13060 => "11000101",13061 => "00011100",13062 => "10000000",13063 => "10101000",13064 => "11110101",13065 => "01101010",13066 => "00100001",13067 => "11000011",13068 => "01010001",13069 => "00010000",13070 => "01111110",13071 => "11011101",13072 => "00111001",13073 => "00010000",13074 => "11111011",13075 => "10001110",13076 => "10100101",13077 => "01110001",13078 => "11110100",13079 => "01111010",13080 => "10001000",13081 => "11010110",13082 => "10011010",13083 => "10110010",13084 => "01101111",13085 => "00100110",13086 => "01100010",13087 => "10010010",13088 => "00101100",13089 => "10101011",13090 => "10110000",13091 => "10000011",13092 => "00010011",13093 => "11000101",13094 => "01011001",13095 => "00010001",13096 => "10111101",13097 => "11010111",13098 => "01111001",13099 => "10101110",13100 => "10001110",13101 => "00011101",13102 => "11000100",13103 => "11101000",13104 => "10001011",13105 => "00001000",13106 => "01011010",13107 => "10011111",13108 => "00011000",13109 => "01111000",13110 => "00010010",13111 => "11000101",13112 => "10001001",13113 => "10000000",13114 => "10111100",13115 => "00001001",13116 => "11011000",13117 => "11111000",13118 => "10110001",13119 => "10101111",13120 => "11100001",13121 => "01010011",13122 => "01000110",13123 => "01010001",13124 => "11110000",13125 => "00010100",13126 => "10100001",13127 => "01001110",13128 => "00100001",13129 => "00011100",13130 => "10011011",13131 => "01000101",13132 => "11110010",13133 => "11111100",13134 => "01001010",13135 => "01100000",13136 => "00011101",13137 => "00110010",13138 => "10011011",13139 => "00110000",13140 => "01010011",13141 => "00100000",13142 => "01001100",13143 => "01111101",13144 => "00011011",13145 => "11011010",13146 => "00011011",13147 => "00010001",13148 => "11000000",13149 => "11011101",13150 => "01001100",13151 => "11101111",13152 => "10111011",13153 => "11001011",13154 => "01101101",13155 => "10110010",13156 => "00100010",13157 => "11100000",13158 => "11100111",13159 => "01011100",13160 => "01010011",13161 => "11010000",13162 => "10010000",13163 => "00111100",13164 => "01101111",13165 => "11111011",13166 => "01100110",13167 => "10010001",13168 => "00100100",13169 => "10100110",13170 => "00110101",13171 => "01101011",13172 => "11111101",13173 => "11011110",13174 => "01010111",13175 => "01000111",13176 => "00011101",13177 => "00101011",13178 => "11000101",13179 => "00111000",13180 => "00111011",13181 => "10111000",13182 => "11001100",13183 => "10001111",13184 => "10111011",13185 => "01010000",13186 => "10111100",13187 => "11011001",13188 => "00101111",13189 => "01100001",13190 => "11001111",13191 => "01000001",13192 => "11000110",13193 => "00111001",13194 => "10110001",13195 => "01111001",13196 => "10111000",13197 => "11101011",13198 => "00110101",13199 => "00110010",13200 => "11101011",13201 => "11101001",13202 => "01001111",13203 => "01101000",13204 => "01110010",13205 => "00010000",13206 => "01110000",13207 => "00000011",13208 => "11111111",13209 => "11011010",13210 => "10100010",13211 => "11010111",13212 => "10110111",13213 => "00101101",13214 => "00101110",13215 => "11001010",13216 => "11010110",13217 => "11010110",13218 => "10110111",13219 => "11101010",13220 => "10000011",13221 => "01101011",13222 => "11000100",13223 => "11011010",13224 => "01111011",13225 => "10001001",13226 => "10010100",13227 => "11101000",13228 => "00010110",13229 => "10101010",13230 => "11000000",13231 => "01101101",13232 => "11010001",13233 => "00100010",13234 => "11111000",13235 => "00011111",13236 => "11100011",13237 => "10100001",13238 => "00110001",13239 => "10111101",13240 => "10110011",13241 => "00101010",13242 => "01011110",13243 => "10000010",13244 => "10010110",13245 => "01011110",13246 => "01111110",13247 => "10111001",13248 => "00101110",13249 => "10001100",13250 => "01011111",13251 => "11110101",13252 => "01000000",13253 => "01101111",13254 => "01010100",13255 => "01000111",13256 => "01000111",13257 => "11101011",13258 => "00110010",13259 => "00011011",13260 => "00100101",13261 => "01110011",13262 => "00000100",13263 => "00000010",13264 => "01100100",13265 => "01010101",13266 => "10111011",13267 => "10001111",13268 => "11100001",13269 => "00101010",13270 => "01000010",13271 => "01000111",13272 => "11100111",13273 => "11010000",13274 => "01101001",13275 => "01101001",13276 => "01101011",13277 => "01000010",13278 => "10001111",13279 => "10011110",13280 => "10000111",13281 => "10000100",13282 => "11000001",13283 => "00011100",13284 => "01110010",13285 => "01110001",13286 => "11000110",13287 => "00001110",13288 => "01111011",13289 => "10010011",13290 => "11010001",13291 => "10010110",13292 => "11110011",13293 => "01111000",13294 => "11101111",13295 => "01100111",13296 => "11110001",13297 => "11111001",13298 => "10100110",13299 => "10101100",13300 => "00011010",13301 => "10010111",13302 => "00011000",13303 => "00001000",13304 => "11110101",13305 => "10101111",13306 => "11101100",13307 => "01110100",13308 => "10001010",13309 => "01110000",13310 => "10110111",13311 => "10101101",13312 => "00000011",13313 => "01011001",13314 => "01100010",13315 => "00101101",13316 => "10101001",13317 => "00100000",13318 => "00100110",13319 => "11000011",13320 => "10010110",13321 => "11010101",13322 => "10100011",13323 => "10100111",13324 => "00010110",13325 => "10100010",13326 => "00100011",13327 => "00001010",13328 => "10010000",13329 => "11101100",13330 => "11100001",13331 => "10101001",13332 => "00000111",13333 => "01110110",13334 => "00011011",13335 => "00110110",13336 => "10010001",13337 => "10111111",13338 => "01101000",13339 => "10011001",13340 => "11101101",13341 => "10001000",13342 => "11001000",13343 => "11100011",13344 => "00011101",13345 => "01111011",13346 => "10101010",13347 => "00110010",13348 => "10010101",13349 => "01100000",13350 => "00011010",13351 => "01011011",13352 => "01100010",13353 => "11110111",13354 => "00100111",13355 => "10000000",13356 => "00010001",13357 => "10011011",13358 => "01010001",13359 => "00011011",13360 => "10000001",13361 => "00011000",13362 => "11011011",13363 => "00000011",13364 => "10010001",13365 => "01010101",13366 => "00101100",13367 => "01011101",13368 => "11101011",13369 => "01001101",13370 => "00011100",13371 => "11111010",13372 => "11101110",13373 => "11110110",13374 => "00000100",13375 => "00100000",13376 => "00000010",13377 => "11101101",13378 => "01110101",13379 => "10110000",13380 => "10000001",13381 => "00110110",13382 => "01000100",13383 => "00011011",13384 => "10010010",13385 => "01101100",13386 => "11111010",13387 => "11111011",13388 => "01001100",13389 => "01110110",13390 => "00001101",13391 => "01111101",13392 => "00111111",13393 => "01010011",13394 => "00100000",13395 => "00111011",13396 => "00111100",13397 => "10010100",13398 => "01000100",13399 => "10110111",13400 => "10011011",13401 => "01110111",13402 => "01011101",13403 => "01110001",13404 => "11101110",13405 => "10011010",13406 => "00011010",13407 => "11100111",13408 => "01111100",13409 => "00000000",13410 => "01011010",13411 => "00100100",13412 => "01110001",13413 => "11100101",13414 => "11000010",13415 => "00100010",13416 => "10101111",13417 => "01100011",13418 => "10101101",13419 => "10011000",13420 => "11010010",13421 => "00011000",13422 => "00001100",13423 => "01010110",13424 => "10001010",13425 => "00011000",13426 => "01011010",13427 => "11100010",13428 => "11011010",13429 => "10010101",13430 => "11001111",13431 => "01111110",13432 => "10101010",13433 => "10111011",13434 => "00000100",13435 => "01100011",13436 => "01110001",13437 => "00101101",13438 => "11000000",13439 => "11010000",13440 => "10011110",13441 => "01000101",13442 => "01110011",13443 => "11111101",13444 => "11001111",13445 => "00000100",13446 => "01101010",13447 => "01101111",13448 => "10011010",13449 => "11101100",13450 => "11111100",13451 => "00111010",13452 => "00101110",13453 => "11110000",13454 => "10010011",13455 => "00110010",13456 => "00011101",13457 => "11111110",13458 => "01111010",13459 => "10100101",13460 => "01111100",13461 => "00111001",13462 => "10110100",13463 => "00011101",13464 => "10011111",13465 => "00010100",13466 => "00110110",13467 => "11000010",13468 => "01000000",13469 => "01011000",13470 => "11011001",13471 => "10010000",13472 => "10010011",13473 => "11101010",13474 => "00110011",13475 => "10010111",13476 => "00001110",13477 => "00001011",13478 => "00010100",13479 => "11111000",13480 => "11100011",13481 => "00001010",13482 => "10011111",13483 => "11100010",13484 => "00001001",13485 => "11110011",13486 => "11110100",13487 => "10011100",13488 => "10110001",13489 => "10100111",13490 => "10001100",13491 => "00101010",13492 => "01010101",13493 => "01100010",13494 => "01110010",13495 => "10000000",13496 => "10110001",13497 => "10010100",13498 => "01111001",13499 => "10010111",13500 => "00110110",13501 => "01001001",13502 => "11011000",13503 => "11110110",13504 => "01010010",13505 => "10111000",13506 => "01011101",13507 => "01110000",13508 => "01000011",13509 => "10001111",13510 => "11000110",13511 => "01100100",13512 => "00110110",13513 => "01010111",13514 => "01110101",13515 => "00111100",13516 => "01110001",13517 => "10010101",13518 => "01100111",13519 => "01110111",13520 => "00111111",13521 => "11001100",13522 => "11101111",13523 => "11100100",13524 => "11011010",13525 => "01100101",13526 => "10000000",13527 => "00101000",13528 => "00100101",13529 => "01110001",13530 => "11110101",13531 => "00011110",13532 => "01111000",13533 => "00000011",13534 => "01101110",13535 => "10011110",13536 => "10010010",13537 => "10110110",13538 => "10000010",13539 => "11100001",13540 => "00011000",13541 => "00011010",13542 => "01101010",13543 => "11100111",13544 => "10100011",13545 => "00011001",13546 => "01010101",13547 => "01110100",13548 => "01010101",13549 => "01011101",13550 => "01001111",13551 => "10110010",13552 => "10001010",13553 => "00001011",13554 => "00010101",13555 => "11111101",13556 => "00000000",13557 => "10001010",13558 => "00100011",13559 => "11101011",13560 => "01011000",13561 => "00011010",13562 => "10011110",13563 => "00110010",13564 => "11010001",13565 => "11011000",13566 => "11111101",13567 => "10100100",13568 => "10010001",13569 => "01011101",13570 => "11111011",13571 => "00100101",13572 => "01101011",13573 => "10001010",13574 => "11111111",13575 => "01011000",13576 => "00011001",13577 => "00000000",13578 => "10010111",13579 => "01110011",13580 => "00011100",13581 => "10111110",13582 => "00001010",13583 => "11100100",13584 => "10011011",13585 => "10011000",13586 => "00101111",13587 => "10001001",13588 => "10101001",13589 => "01011100",13590 => "00011110",13591 => "10110101",13592 => "01101011",13593 => "10111001",13594 => "11111011",13595 => "11000011",13596 => "11001000",13597 => "01000001",13598 => "11111000",13599 => "11010110",13600 => "00001001",13601 => "01011010",13602 => "10101100",13603 => "00101000",13604 => "10111001",13605 => "10000011",13606 => "10101111",13607 => "00011000",13608 => "11001010",13609 => "11010110",13610 => "01110100",13611 => "01100100",13612 => "11100100",13613 => "00011010",13614 => "00110010",13615 => "01101001",13616 => "01110000",13617 => "11011100",13618 => "11000100",13619 => "11110100",13620 => "11010011",13621 => "11110001",13622 => "11111010",13623 => "01010011",13624 => "00010010",13625 => "00110011",13626 => "01111100",13627 => "00111011",13628 => "11011011",13629 => "11111101",13630 => "11110000",13631 => "00000100",13632 => "00101101",13633 => "10110010",13634 => "01000111",13635 => "00000001",13636 => "11001110",13637 => "01101010",13638 => "01010110",13639 => "10101100",13640 => "00010011",13641 => "10011101",13642 => "00011111",13643 => "11100001",13644 => "01110000",13645 => "00000011",13646 => "00110000",13647 => "01101010",13648 => "11110010",13649 => "00100111",13650 => "10011111",13651 => "11101011",13652 => "00001110",13653 => "10010100",13654 => "11011110",13655 => "11010100",13656 => "10001011",13657 => "10100111",13658 => "00101110",13659 => "11011100",13660 => "11010011",13661 => "01001000",13662 => "01011110",13663 => "11110111",13664 => "10011101",13665 => "10111100",13666 => "00000000",13667 => "10111101",13668 => "10000000",13669 => "10011111",13670 => "11100110",13671 => "11111100",13672 => "10100110",13673 => "01100000",13674 => "11110001",13675 => "11101001",13676 => "00100001",13677 => "11001100",13678 => "10101101",13679 => "00110101",13680 => "01011011",13681 => "10010110",13682 => "00001110",13683 => "10001000",13684 => "01111111",13685 => "10101110",13686 => "00010100",13687 => "11101101",13688 => "00111011",13689 => "00011111",13690 => "10011000",13691 => "11001000",13692 => "00000111",13693 => "11101000",13694 => "00101100",13695 => "01101101",13696 => "11110000",13697 => "10001100",13698 => "00111110",13699 => "01100010",13700 => "00011010",13701 => "01111111",13702 => "01110001",13703 => "11011010",13704 => "11111100",13705 => "11100001",13706 => "01100110",13707 => "01011010",13708 => "10101100",13709 => "10001010",13710 => "01010010",13711 => "11101100",13712 => "11110111",13713 => "00000100",13714 => "10011100",13715 => "11001110",13716 => "11100100",13717 => "00011101",13718 => "00110010",13719 => "11001110",13720 => "00101010",13721 => "00100000",13722 => "01111101",13723 => "10110000",13724 => "10100101",13725 => "00110010",13726 => "10111100",13727 => "11101010",13728 => "10011011",13729 => "11001001",13730 => "11101100",13731 => "10001001",13732 => "11000001",13733 => "00001010",13734 => "01001000",13735 => "11001101",13736 => "00010110",13737 => "00011111",13738 => "01001010",13739 => "10000100",13740 => "01011010",13741 => "10101010",13742 => "00111001",13743 => "01001100",13744 => "11101111",13745 => "11101100",13746 => "11111100",13747 => "10101000",13748 => "01010001",13749 => "10110011",13750 => "01110111",13751 => "00001111",13752 => "01111101",13753 => "01010101",13754 => "00011101",13755 => "11101011",13756 => "01011011",13757 => "00010101",13758 => "01110111",13759 => "01111011",13760 => "11110101",13761 => "10010100",13762 => "10000101",13763 => "00011001",13764 => "00000000",13765 => "00111000",13766 => "00100001",13767 => "01010011",13768 => "11000001",13769 => "10010110",13770 => "00111001",13771 => "10100001",13772 => "11001100",13773 => "00010101",13774 => "00001010",13775 => "11110101",13776 => "10100111",13777 => "10100001",13778 => "10000110",13779 => "11110111",13780 => "11111000",13781 => "01011101",13782 => "01111011",13783 => "10010001",13784 => "01001001",13785 => "00000011",13786 => "10011101",13787 => "11000001",13788 => "11111111",13789 => "00101000",13790 => "00000100",13791 => "01000111",13792 => "01001000",13793 => "00001010",13794 => "10010110",13795 => "01011010",13796 => "11101000",13797 => "10011110",13798 => "10000000",13799 => "01011000",13800 => "11100011",13801 => "11101010",13802 => "11101100",13803 => "11011111",13804 => "01011100",13805 => "00001010",13806 => "00101100",13807 => "11111001",13808 => "01110111",13809 => "00110111",13810 => "11011010",13811 => "01101000",13812 => "01110000",13813 => "11001100",13814 => "10110111",13815 => "11010000",13816 => "10001100",13817 => "11010011",13818 => "11100110",13819 => "10111010",13820 => "00101110",13821 => "01111100",13822 => "00011111",13823 => "01000010",13824 => "01110001",13825 => "00110001",13826 => "01011100",13827 => "11101111",13828 => "00100111",13829 => "00110111",13830 => "00001110",13831 => "01000111",13832 => "11011101",13833 => "01011110",13834 => "10111001",13835 => "00101010",13836 => "11101000",13837 => "11100111",13838 => "01010011",13839 => "10010000",13840 => "10011100",13841 => "10011110",13842 => "01010100",13843 => "00101110",13844 => "10110101",13845 => "00110010",13846 => "00001101",13847 => "10001010",13848 => "00010110",13849 => "01100101",13850 => "01110001",13851 => "01111011",13852 => "10000110",13853 => "01000111",13854 => "00011011",13855 => "10011010",13856 => "11011101",13857 => "11110000",13858 => "10010011",13859 => "00001000",13860 => "11011010",13861 => "11101111",13862 => "10011001",13863 => "01100100",13864 => "01010000",13865 => "11011001",13866 => "10011001",13867 => "00010011",13868 => "00000111",13869 => "10011110",13870 => "00001101",13871 => "10010100",13872 => "11110010",13873 => "10101010",13874 => "10001010",13875 => "00010001",13876 => "01101101",13877 => "01100110",13878 => "10001011",13879 => "10000010",13880 => "11101001",13881 => "00101111",13882 => "01000000",13883 => "01111110",13884 => "10011110",13885 => "10001001",13886 => "10000100",13887 => "11101000",13888 => "10100100",13889 => "00010001",13890 => "11111101",13891 => "10010000",13892 => "00110101",13893 => "01111011",13894 => "11000000",13895 => "01010001",13896 => "10011011",13897 => "00010000",13898 => "00101101",13899 => "00110001",13900 => "01111111",13901 => "01111110",13902 => "11011100",13903 => "10000001",13904 => "00101100",13905 => "00010111",13906 => "10001101",13907 => "11001001",13908 => "11000101",13909 => "11010001",13910 => "10101111",13911 => "10000101",13912 => "01101000",13913 => "00010111",13914 => "01011101",13915 => "10110010",13916 => "10100111",13917 => "11110011",13918 => "00101011",13919 => "10100101",13920 => "11001111",13921 => "11111011",13922 => "11001000",13923 => "01100001",13924 => "00101111",13925 => "10101001",13926 => "11000001",13927 => "10100011",13928 => "01001001",13929 => "01101000",13930 => "00010110",13931 => "00110010",13932 => "11100111",13933 => "01110101",13934 => "01101110",13935 => "11010110",13936 => "00000100",13937 => "01110110",13938 => "10000110",13939 => "10101011",13940 => "01101010",13941 => "11100110",13942 => "01100010",13943 => "00110001",13944 => "10011000",13945 => "01010010",13946 => "01101100",13947 => "00011010",13948 => "10110110",13949 => "01011001",13950 => "11001001",13951 => "00000111",13952 => "00011100",13953 => "10010111",13954 => "01000011",13955 => "10011000",13956 => "00011000",13957 => "11101000",13958 => "11111001",13959 => "00000100",13960 => "11100001",13961 => "11100001",13962 => "10110001",13963 => "11010100",13964 => "10010100",13965 => "11001110",13966 => "00001001",13967 => "01011101",13968 => "10111101",13969 => "00111011",13970 => "10001101",13971 => "01001011",13972 => "01111001",13973 => "11000111",13974 => "01000111",13975 => "00111101",13976 => "01010111",13977 => "10110110",13978 => "00110001",13979 => "11110110",13980 => "01101011",13981 => "01111111",13982 => "11001001",13983 => "11010001",13984 => "11001110",13985 => "11011001",13986 => "11010000",13987 => "01100110",13988 => "01011100",13989 => "11011011",13990 => "11111011",13991 => "11001101",13992 => "11100000",13993 => "01001101",13994 => "10011111",13995 => "10010001",13996 => "00010100",13997 => "11111111",13998 => "01111110",13999 => "10011000",14000 => "01110010",14001 => "01100011",14002 => "00111011",14003 => "11111011",14004 => "01101111",14005 => "11000000",14006 => "11011100",14007 => "10001001",14008 => "00011000",14009 => "11000101",14010 => "01000001",14011 => "00101000",14012 => "10010101",14013 => "10010000",14014 => "11100100",14015 => "11101111",14016 => "01001100",14017 => "01000101",14018 => "01000101",14019 => "11100101",14020 => "00011000",14021 => "10011010",14022 => "00100000",14023 => "10100100",14024 => "01110001",14025 => "10100101",14026 => "11110010",14027 => "10000101",14028 => "11001101",14029 => "11101011",14030 => "01111101",14031 => "10000101",14032 => "00000101",14033 => "01100000",14034 => "01101000",14035 => "10111011",14036 => "01010011",14037 => "10101011",14038 => "01100000",14039 => "00101001",14040 => "00111100",14041 => "01000000",14042 => "00101010",14043 => "11001100",14044 => "11101100",14045 => "11010110",14046 => "11111100",14047 => "01010101",14048 => "10001001",14049 => "10111001",14050 => "01111101",14051 => "11001100",14052 => "11111111",14053 => "10111100",14054 => "00000101",14055 => "00001111",14056 => "11101011",14057 => "11110001",14058 => "01101011",14059 => "11001011",14060 => "00110010",14061 => "11101111",14062 => "10100011",14063 => "00111000",14064 => "11010010",14065 => "10101000",14066 => "00111000",14067 => "11111100",14068 => "00100001",14069 => "10000100",14070 => "00010110",14071 => "01010100",14072 => "00011111",14073 => "01110100",14074 => "00100001",14075 => "11111011",14076 => "01100000",14077 => "00000100",14078 => "10000100",14079 => "10101100",14080 => "10001001",14081 => "10010011",14082 => "01100110",14083 => "11111110",14084 => "10010011",14085 => "00011110",14086 => "10110000",14087 => "11011010",14088 => "01110000",14089 => "00101101",14090 => "10001001",14091 => "11111100",14092 => "01011110",14093 => "00110110",14094 => "11100100",14095 => "10000100",14096 => "10011010",14097 => "10010011",14098 => "00001000",14099 => "00111100",14100 => "11101100",14101 => "10000111",14102 => "01101000",14103 => "00101101",14104 => "11001001",14105 => "01000010",14106 => "01111010",14107 => "10101011",14108 => "00110110",14109 => "01010011",14110 => "11101010",14111 => "10010010",14112 => "10110110",14113 => "10100000",14114 => "00011110",14115 => "00100011",14116 => "11010000",14117 => "11110100",14118 => "00011101",14119 => "00000110",14120 => "10001001",14121 => "10010001",14122 => "00000000",14123 => "10010100",14124 => "11010001",14125 => "11001100",14126 => "11111111",14127 => "11011010",14128 => "00111110",14129 => "11111001",14130 => "00010010",14131 => "10111000",14132 => "10100100",14133 => "10010100",14134 => "01010001",14135 => "01011010",14136 => "00101100",14137 => "11011000",14138 => "00000101",14139 => "00110001",14140 => "01110000",14141 => "11010001",14142 => "01100000",14143 => "00011011",14144 => "11010000",14145 => "11011000",14146 => "11111010",14147 => "10110000",14148 => "11111110",14149 => "10000111",14150 => "01011000",14151 => "01011001",14152 => "01111001",14153 => "10001010",14154 => "01111100",14155 => "11011000",14156 => "00000010",14157 => "01001000",14158 => "01011011",14159 => "10111010",14160 => "00011100",14161 => "11000100",14162 => "10100111",14163 => "11110101",14164 => "01001100",14165 => "00011101",14166 => "11110111",14167 => "10111100",14168 => "01000000",14169 => "11101111",14170 => "11101011",14171 => "00000100",14172 => "11101110",14173 => "00101101",14174 => "10000111",14175 => "11011001",14176 => "10000010",14177 => "00100100",14178 => "10001011",14179 => "00110001",14180 => "10100111",14181 => "00111001",14182 => "11000010",14183 => "10101111",14184 => "01101010",14185 => "10111101",14186 => "00100101",14187 => "11111110",14188 => "10010010",14189 => "00010010",14190 => "01111101",14191 => "11001001",14192 => "00000010",14193 => "01111111",14194 => "00101011",14195 => "10011101",14196 => "00101100",14197 => "10001110",14198 => "11011011",14199 => "00110000",14200 => "01010001",14201 => "11100010",14202 => "10011110",14203 => "00101110",14204 => "00000110",14205 => "11110000",14206 => "00101001",14207 => "11000101",14208 => "10001110",14209 => "11010011",14210 => "01000101",14211 => "10010111",14212 => "11101111",14213 => "10100100",14214 => "00000000",14215 => "01110110",14216 => "01010101",14217 => "01100010",14218 => "11010110",14219 => "00010011",14220 => "01111111",14221 => "11100110",14222 => "11101101",14223 => "10110100",14224 => "10101010",14225 => "11101101",14226 => "11000101",14227 => "00111110",14228 => "01100011",14229 => "10110110",14230 => "00110111",14231 => "01000110",14232 => "11011110",14233 => "01001100",14234 => "10101011",14235 => "10100011",14236 => "11001110",14237 => "00100010",14238 => "10110001",14239 => "01111100",14240 => "11110100",14241 => "01000111",14242 => "10011100",14243 => "11011011",14244 => "01111011",14245 => "01000010",14246 => "11011111",14247 => "01110001",14248 => "10111100",14249 => "10010110",14250 => "11000000",14251 => "00111010",14252 => "01001100",14253 => "11001011",14254 => "00010010",14255 => "00111001",14256 => "01111111",14257 => "11010111",14258 => "01101101",14259 => "10110000",14260 => "01110000",14261 => "11111110",14262 => "11111100",14263 => "01101011",14264 => "11001011",14265 => "00101001",14266 => "10111011",14267 => "00111010",14268 => "01100101",14269 => "10000011",14270 => "10100111",14271 => "10011011",14272 => "11011011",14273 => "11101001",14274 => "10111100",14275 => "01010101",14276 => "10111100",14277 => "01111101",14278 => "11110011",14279 => "00000011",14280 => "11000010",14281 => "00000000",14282 => "10001000",14283 => "10110111",14284 => "01111100",14285 => "00101111",14286 => "10101110",14287 => "00001111",14288 => "00110011",14289 => "11111110",14290 => "11110100",14291 => "00011110",14292 => "11100101",14293 => "00000101",14294 => "00110001",14295 => "10001001",14296 => "11110001",14297 => "00011101",14298 => "10111001",14299 => "00011100",14300 => "11001111",14301 => "00111101",14302 => "11011000",14303 => "11010001",14304 => "10110110",14305 => "11010111",14306 => "01101000",14307 => "01111111",14308 => "11000111",14309 => "00111010",14310 => "01110100",14311 => "10111110",14312 => "00010111",14313 => "00001110",14314 => "10010010",14315 => "10110001",14316 => "00001011",14317 => "10001110",14318 => "01111011",14319 => "11011100",14320 => "10010001",14321 => "01010000",14322 => "11101110",14323 => "00011111",14324 => "10011110",14325 => "11000110",14326 => "00011001",14327 => "01111100",14328 => "11001000",14329 => "01011111",14330 => "11111100",14331 => "11011110",14332 => "10110011",14333 => "01000111",14334 => "11001000",14335 => "11010110",14336 => "10101000",14337 => "00100001",14338 => "11100001",14339 => "01000100",14340 => "01111000",14341 => "00001010",14342 => "00100010",14343 => "00100011",14344 => "00110010",14345 => "10111111",14346 => "10110000",14347 => "00110000",14348 => "10111100",14349 => "01110101",14350 => "11111010",14351 => "10111000",14352 => "10111101",14353 => "01110011",14354 => "11010010",14355 => "01011011",14356 => "01010001",14357 => "11010100",14358 => "10000101",14359 => "01100100",14360 => "10111101",14361 => "01110100",14362 => "11001100",14363 => "00011010",14364 => "10011110",14365 => "01000011",14366 => "01100001",14367 => "11001111",14368 => "01110100",14369 => "00111001",14370 => "10111010",14371 => "10110011",14372 => "01011101",14373 => "11001000",14374 => "10100101",14375 => "11011010",14376 => "00110101",14377 => "10010111",14378 => "01101110",14379 => "00110001",14380 => "01001101",14381 => "00001110",14382 => "11100100",14383 => "11110111",14384 => "00001010",14385 => "01000001",14386 => "01011110",14387 => "00000111",14388 => "10110111",14389 => "10011011",14390 => "11011001",14391 => "01011000",14392 => "10111010",14393 => "01000000",14394 => "10011100",14395 => "01101001",14396 => "00000001",14397 => "00110101",14398 => "11000010",14399 => "11101101",14400 => "00100011",14401 => "00011101",14402 => "11110100",14403 => "00000100",14404 => "11101001",14405 => "11000100",14406 => "11100010",14407 => "10010001",14408 => "00111011",14409 => "00100001",14410 => "00100001",14411 => "11010001",14412 => "11111010",14413 => "01010101",14414 => "10100011",14415 => "00100011",14416 => "01110000",14417 => "00010000",14418 => "00110111",14419 => "00101110",14420 => "10110100",14421 => "10011110",14422 => "00101111",14423 => "10110101",14424 => "10110011",14425 => "01101000",14426 => "00000001",14427 => "01010010",14428 => "11011110",14429 => "01110010",14430 => "00101000",14431 => "11001101",14432 => "11001111",14433 => "01000101",14434 => "01000010",14435 => "10010110",14436 => "00101111",14437 => "11000101",14438 => "11111100",14439 => "01001100",14440 => "11101000",14441 => "10111101",14442 => "11001010",14443 => "01111110",14444 => "11111101",14445 => "00001100",14446 => "00000000",14447 => "01011111",14448 => "10101100",14449 => "10111000",14450 => "11111011",14451 => "00111100",14452 => "01000010",14453 => "11100010",14454 => "10011110",14455 => "10001100",14456 => "10100101",14457 => "10111001",14458 => "01000100",14459 => "10010000",14460 => "11111001",14461 => "01000110",14462 => "11111000",14463 => "11001110",14464 => "11010111",14465 => "01100011",14466 => "10000000",14467 => "10110111",14468 => "11100101",14469 => "10101100",14470 => "01110011",14471 => "00011010",14472 => "11101001",14473 => "10100111",14474 => "11000110",14475 => "10110011",14476 => "01010001",14477 => "01000111",14478 => "11100111",14479 => "11000001",14480 => "01001101",14481 => "11101011",14482 => "10010110",14483 => "10010101",14484 => "00110000",14485 => "01100011",14486 => "11111001",14487 => "10011100",14488 => "11101110",14489 => "11110011",14490 => "01101110",14491 => "10101010",14492 => "11100101",14493 => "10111110",14494 => "00111111",14495 => "11111110",14496 => "11001000",14497 => "11001100",14498 => "10111100",14499 => "11000001",14500 => "10010001",14501 => "10101101",14502 => "00000100",14503 => "00000010",14504 => "10110101",14505 => "10001111",14506 => "01110000",14507 => "10010010",14508 => "01010011",14509 => "11100000",14510 => "01010111",14511 => "10000001",14512 => "10010010",14513 => "00111101",14514 => "11001101",14515 => "11111100",14516 => "10100001",14517 => "11101010",14518 => "00110010",14519 => "00010100",14520 => "11000110",14521 => "10101011",14522 => "10100000",14523 => "01110011",14524 => "01101010",14525 => "01110100",14526 => "11110101",14527 => "01000111",14528 => "11011101",14529 => "00101100",14530 => "01111010",14531 => "11111010",14532 => "01101110",14533 => "10110111",14534 => "00111100",14535 => "00010111",14536 => "00001011",14537 => "00111111",14538 => "00100101",14539 => "10101101",14540 => "01010111",14541 => "00011101",14542 => "00101011",14543 => "10011010",14544 => "01111000",14545 => "10101010",14546 => "01110010",14547 => "00101110",14548 => "00010011",14549 => "10011100",14550 => "11100100",14551 => "10000000",14552 => "00111000",14553 => "11001000",14554 => "11001011",14555 => "10111110",14556 => "11111000",14557 => "01110101",14558 => "01101010",14559 => "01010100",14560 => "10101000",14561 => "00111101",14562 => "10111010",14563 => "01110111",14564 => "11011000",14565 => "01100110",14566 => "01011010",14567 => "01001100",14568 => "00001011",14569 => "10100110",14570 => "11010000",14571 => "11001101",14572 => "10111011",14573 => "00111101",14574 => "10011111",14575 => "11100110",14576 => "10001110",14577 => "01000110",14578 => "11000011",14579 => "00110011",14580 => "01110111",14581 => "10101101",14582 => "00010001",14583 => "11100000",14584 => "00110110",14585 => "00100010",14586 => "00110011",14587 => "11110000",14588 => "01010001",14589 => "00000001",14590 => "01010000",14591 => "00110011",14592 => "10110101",14593 => "10110011",14594 => "11111111",14595 => "11010100",14596 => "10100011",14597 => "00001011",14598 => "01101101",14599 => "01001101",14600 => "10010010",14601 => "00000000",14602 => "01100101",14603 => "00001111",14604 => "01101000",14605 => "10010010",14606 => "11000000",14607 => "10100000",14608 => "10001111",14609 => "01000101",14610 => "10111111",14611 => "11011110",14612 => "00100100",14613 => "11100011",14614 => "11101010",14615 => "00011111",14616 => "01001110",14617 => "00101010",14618 => "11001110",14619 => "01101001",14620 => "00001010",14621 => "01011101",14622 => "00110000",14623 => "00110111",14624 => "11111111",14625 => "01010111",14626 => "00110111",14627 => "00010110",14628 => "11011100",14629 => "01010101",14630 => "01101110",14631 => "00101001",14632 => "00001001",14633 => "00011101",14634 => "11011011",14635 => "00010101",14636 => "11011101",14637 => "11101001",14638 => "00101011",14639 => "00101100",14640 => "10000001",14641 => "00010010",14642 => "01010111",14643 => "00010000",14644 => "00010001",14645 => "11110010",14646 => "11011010",14647 => "11010001",14648 => "10111111",14649 => "10100000",14650 => "10010100",14651 => "00001000",14652 => "01101111",14653 => "11101110",14654 => "01011111",14655 => "00101011",14656 => "10111101",14657 => "10111100",14658 => "01100010",14659 => "10110100",14660 => "11100010",14661 => "00100001",14662 => "11111001",14663 => "10110010",14664 => "10100010",14665 => "10001100",14666 => "00110010",14667 => "10010100",14668 => "00101111",14669 => "10011100",14670 => "11101001",14671 => "10111100",14672 => "01100010",14673 => "10010000",14674 => "01001110",14675 => "00111101",14676 => "01001101",14677 => "00101010",14678 => "00101110",14679 => "10011110",14680 => "01011100",14681 => "10100001",14682 => "11101111",14683 => "10000101",14684 => "01001010",14685 => "11000011",14686 => "01001010",14687 => "00101100",14688 => "01010110",14689 => "11000101",14690 => "11100100",14691 => "00001110",14692 => "11111001",14693 => "00100100",14694 => "11011010",14695 => "10100000",14696 => "00101000",14697 => "11010100",14698 => "01110010",14699 => "11101111",14700 => "10110100",14701 => "00101110",14702 => "01100110",14703 => "00101011",14704 => "11110011",14705 => "00111111",14706 => "11001011",14707 => "00110010",14708 => "01110011",14709 => "10001111",14710 => "11000000",14711 => "10011001",14712 => "10110101",14713 => "10011110",14714 => "00101100",14715 => "01100001",14716 => "11011000",14717 => "00010110",14718 => "01000000",14719 => "00101100",14720 => "00001100",14721 => "00011111",14722 => "00100110",14723 => "01101111",14724 => "10000011",14725 => "10001101",14726 => "10101011",14727 => "00010001",14728 => "01111111",14729 => "10110000",14730 => "00111101",14731 => "10110010",14732 => "11100111",14733 => "01110000",14734 => "11100100",14735 => "01000101",14736 => "00110011",14737 => "00010101",14738 => "01101011",14739 => "00111000",14740 => "11011110",14741 => "01111100",14742 => "11001111",14743 => "00111011",14744 => "11100111",14745 => "11110110",14746 => "01100111",14747 => "10111011",14748 => "01100100",14749 => "10100001",14750 => "00110011",14751 => "11010100",14752 => "01110000",14753 => "10110101",14754 => "10110001",14755 => "10010101",14756 => "10101101",14757 => "10010110",14758 => "01000000",14759 => "01000001",14760 => "00010000",14761 => "00100000",14762 => "00010110",14763 => "10100100",14764 => "00010111",14765 => "10111100",14766 => "11111101",14767 => "10110010",14768 => "11001000",14769 => "01110101",14770 => "10010100",14771 => "01111100",14772 => "00111101",14773 => "00000011",14774 => "00001100",14775 => "00101110",14776 => "11111001",14777 => "01110001",14778 => "10010000",14779 => "11000111",14780 => "10110100",14781 => "11110101",14782 => "00100110",14783 => "11101100",14784 => "01100111",14785 => "00100011",14786 => "00100110",14787 => "10001011",14788 => "01010011",14789 => "00010100",14790 => "01010110",14791 => "11111011",14792 => "10100101",14793 => "00001011",14794 => "11000100",14795 => "11100011",14796 => "00100101",14797 => "11111011",14798 => "11001110",14799 => "10000111",14800 => "00111101",14801 => "10100010",14802 => "11111100",14803 => "00011000",14804 => "10101001",14805 => "00010101",14806 => "00110001",14807 => "01010111",14808 => "00011000",14809 => "10011101",14810 => "10000011",14811 => "01110010",14812 => "11111011",14813 => "10110110",14814 => "11100000",14815 => "01011111",14816 => "00110111",14817 => "11100001",14818 => "11000111",14819 => "11110000",14820 => "10011010",14821 => "10111110",14822 => "00000001",14823 => "11001010",14824 => "10000011",14825 => "00101000",14826 => "00011011",14827 => "01011001",14828 => "00010101",14829 => "00010001",14830 => "10111010",14831 => "10010010",14832 => "10000000",14833 => "11110001",14834 => "10011010",14835 => "01000000",14836 => "11101001",14837 => "11101011",14838 => "10011010",14839 => "01100000",14840 => "00001101",14841 => "01111100",14842 => "01101101",14843 => "00011111",14844 => "00110000",14845 => "11110100",14846 => "00010001",14847 => "01011101",14848 => "00101001",14849 => "11101000",14850 => "11001010",14851 => "01010001",14852 => "01001101",14853 => "10011011",14854 => "11010011",14855 => "01101110",14856 => "00011100",14857 => "10000010",14858 => "10000010",14859 => "00001000",14860 => "10110110",14861 => "01001001",14862 => "01110011",14863 => "01001001",14864 => "10110011",14865 => "10110011",14866 => "01000101",14867 => "01001110",14868 => "11101000",14869 => "11111101",14870 => "01001000",14871 => "10101001",14872 => "10001010",14873 => "00011101",14874 => "11000111",14875 => "11100001",14876 => "11111101",14877 => "11010100",14878 => "01101110",14879 => "01001101",14880 => "10000010",14881 => "00011101",14882 => "11101001",14883 => "11111011",14884 => "11011010",14885 => "00001100",14886 => "10001010",14887 => "01100010",14888 => "11101000",14889 => "00000101",14890 => "00111000",14891 => "01001001",14892 => "00110100",14893 => "10110100",14894 => "01111001",14895 => "01000101",14896 => "11000010",14897 => "11101001",14898 => "00111010",14899 => "10110100",14900 => "01010100",14901 => "11011000",14902 => "01001111",14903 => "00101100",14904 => "00010000",14905 => "00111100",14906 => "01010100",14907 => "01010011",14908 => "11010100",14909 => "10101011",14910 => "11000111",14911 => "01101010",14912 => "11010011",14913 => "00100000",14914 => "01011010",14915 => "10101111",14916 => "01011110",14917 => "01011110",14918 => "10011000",14919 => "11000111",14920 => "00100011",14921 => "01111101",14922 => "11111010",14923 => "11000111",14924 => "10111100",14925 => "00010010",14926 => "11111000",14927 => "00101110",14928 => "10011110",14929 => "11000000",14930 => "00010101",14931 => "01011100",14932 => "10100011",14933 => "01110000",14934 => "10111000",14935 => "00101010",14936 => "10000000",14937 => "01100000",14938 => "01010101",14939 => "11000110",14940 => "01100100",14941 => "00101000",14942 => "11111011",14943 => "00100001",14944 => "01001100",14945 => "11110001",14946 => "11000101",14947 => "10011111",14948 => "01001101",14949 => "01111101",14950 => "10101111",14951 => "11111000",14952 => "00101001",14953 => "10110111",14954 => "11001001",14955 => "10111110",14956 => "00000000",14957 => "01100000",14958 => "00100011",14959 => "10010100",14960 => "11101010",14961 => "11110111",14962 => "11100111",14963 => "00100110",14964 => "01000100",14965 => "10001011",14966 => "00011101",14967 => "00110000",14968 => "10110101",14969 => "00001010",14970 => "00111011",14971 => "10000000",14972 => "10000000",14973 => "00110110",14974 => "11010000",14975 => "11010110",14976 => "10110111",14977 => "11011000",14978 => "00010100",14979 => "11010011",14980 => "00101100",14981 => "00110110",14982 => "01111110",14983 => "00111101",14984 => "10101100",14985 => "01011011",14986 => "01100111",14987 => "00101110",14988 => "10111111",14989 => "00000100",14990 => "00011111",14991 => "01010000",14992 => "00100111",14993 => "11101111",14994 => "11000011",14995 => "01110110",14996 => "01111101",14997 => "10110101",14998 => "01100011",14999 => "11001111",15000 => "10001001",15001 => "11001001",15002 => "00010000",15003 => "10100100",15004 => "00110000",15005 => "00000011",15006 => "11010101",15007 => "01001100",15008 => "00101101",15009 => "10010110",15010 => "10001000",15011 => "00000010",15012 => "01010100",15013 => "01000111",15014 => "01011111",15015 => "00010001",15016 => "01010101",15017 => "01001100",15018 => "11111000",15019 => "11110011",15020 => "00011111",15021 => "00001001",15022 => "00100001",15023 => "00000110",15024 => "00000100",15025 => "00101001",15026 => "00110100",15027 => "00000010",15028 => "10101100",15029 => "01011001",15030 => "11000101",15031 => "00110111",15032 => "01110011",15033 => "01101100",15034 => "10110101",15035 => "11000011",15036 => "11111110",15037 => "01101001",15038 => "00101010",15039 => "10011001",15040 => "10101011",15041 => "11001111",15042 => "00101011",15043 => "01000111",15044 => "11100101",15045 => "00010111",15046 => "00101110",15047 => "10010010",15048 => "10110111",15049 => "00011111",15050 => "10001010",15051 => "10110111",15052 => "11001111",15053 => "11001100",15054 => "00001000",15055 => "00110111",15056 => "01011000",15057 => "00011001",15058 => "00011000",15059 => "00101001",15060 => "01101010",15061 => "10110110",15062 => "11011111",15063 => "01101100",15064 => "10010110",15065 => "11000010",15066 => "01010010",15067 => "01101100",15068 => "11011010",15069 => "00000110",15070 => "01100000",15071 => "11011000",15072 => "10001110",15073 => "10110101",15074 => "11010100",15075 => "10100110",15076 => "00001001",15077 => "01101100",15078 => "01110111",15079 => "10010100",15080 => "00101000",15081 => "11011101",15082 => "01001110",15083 => "11001110",15084 => "10011000",15085 => "00001011",15086 => "11011110",15087 => "10001011",15088 => "10110010",15089 => "11011001",15090 => "11010010",15091 => "00001001",15092 => "10100000",15093 => "10111000",15094 => "01000100",15095 => "10110000",15096 => "00110000",15097 => "00101000",15098 => "00001011",15099 => "11000111",15100 => "11010001",15101 => "11100100",15102 => "01001001",15103 => "01000001",15104 => "11000001",15105 => "00010100",15106 => "00010101",15107 => "11111100",15108 => "01110100",15109 => "10010111",15110 => "00000100",15111 => "01100010",15112 => "00110001",15113 => "11010010",15114 => "01011000",15115 => "10100010",15116 => "00101010",15117 => "01011000",15118 => "01110011",15119 => "01000000",15120 => "01011011",15121 => "10010111",15122 => "10110010",15123 => "11111011",15124 => "00111001",15125 => "00100110",15126 => "01001010",15127 => "10111010",15128 => "01101000",15129 => "11110110",15130 => "01101100",15131 => "10110111",15132 => "01111100",15133 => "11101001",15134 => "01100000",15135 => "11111101",15136 => "01010110",15137 => "01010111",15138 => "11100101",15139 => "01110100",15140 => "01101100",15141 => "10011001",15142 => "11110100",15143 => "00110100",15144 => "00111010",15145 => "00110000",15146 => "00101101",15147 => "00111100",15148 => "01010001",15149 => "10100100",15150 => "11010111",15151 => "11000001",15152 => "10111001",15153 => "01000101",15154 => "11101111",15155 => "00001111",15156 => "10011010",15157 => "01110000",15158 => "11100000",15159 => "01111011",15160 => "01000011",15161 => "11111000",15162 => "10000111",15163 => "00110101",15164 => "11001011",15165 => "10010010",15166 => "00100101",15167 => "11110100",15168 => "01011001",15169 => "11001110",15170 => "01100111",15171 => "00101011",15172 => "00110111",15173 => "10100010",15174 => "11001111",15175 => "10111000",15176 => "10011111",15177 => "00001000",15178 => "00000101",15179 => "00101101",15180 => "01010100",15181 => "11111100",15182 => "01111010",15183 => "00110100",15184 => "11000100",15185 => "11101000",15186 => "01110001",15187 => "10011011",15188 => "01101100",15189 => "11110000",15190 => "00011001",15191 => "00111000",15192 => "00001100",15193 => "11011001",15194 => "10001110",15195 => "00101000",15196 => "11000111",15197 => "01111001",15198 => "00110010",15199 => "00110100",15200 => "10010101",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00111011" report "FAIL high bits" severity failure;
assert RAM(0) = "01100000" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
