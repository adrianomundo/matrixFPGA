 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01101010",3 => "10001010",4 => "10000011",5 => "00100010",6 => "00010010",7 => "00111001",8 => "10101111",9 => "00010101",10 => "01000001",11 => "11100100",12 => "11101011",13 => "11100110",14 => "01110011",15 => "10011011",16 => "00111011",17 => "11100111",18 => "11100011",19 => "01111101",20 => "11111000",21 => "10001111",22 => "10001101",23 => "01100100",24 => "10101001",25 => "00011010",26 => "01000110",27 => "00111011",28 => "11110001",29 => "00111110",30 => "01111010",31 => "10011100",32 => "01011110",33 => "11100101",34 => "11101110",35 => "10101001",36 => "00001111",37 => "11011001",38 => "01111111",39 => "00100101",40 => "00110101",41 => "01101101",42 => "10010011",43 => "11011111",44 => "11011100",45 => "01110011",46 => "00011001",47 => "11011011",48 => "11111000",49 => "11110111",50 => "01011010",51 => "10100001",52 => "10110000",53 => "00010110",54 => "00110101",55 => "11110011",56 => "10000001",57 => "00010110",58 => "10010101",59 => "00001001",60 => "11111101",61 => "10101010",62 => "01010011",63 => "11011100",64 => "01000011",65 => "11000010",66 => "11101000",67 => "00010000",68 => "00000000",69 => "00010001",70 => "11110010",71 => "11110011",72 => "01111001",73 => "10110001",74 => "10110001",75 => "11000110",76 => "01101101",77 => "00001000",78 => "01010011",79 => "01011010",80 => "11101111",81 => "00101100",82 => "11101111",83 => "11110000",84 => "01010000",85 => "01000110",86 => "01100101",87 => "10011110",88 => "10011010",89 => "00110110",90 => "11010000",91 => "10000111",92 => "11000100",93 => "00001001",94 => "10010011",95 => "10001100",96 => "01101100",97 => "11000111",98 => "00001100",99 => "00100111",100 => "01100011",101 => "10100001",102 => "01110101",103 => "10001111",104 => "11001000",105 => "11010110",106 => "10010100",107 => "10110011",108 => "01001011",109 => "01001110",110 => "00000010",111 => "01101010",112 => "11110111",113 => "10010110",114 => "11001110",115 => "01110110",116 => "10110111",117 => "11010001",118 => "01110010",119 => "11101100",120 => "00100111",121 => "10010000",122 => "10100100",123 => "01010110",124 => "01001000",125 => "01011010",126 => "00100111",127 => "11100000",128 => "11100011",129 => "11000100",130 => "01000110",131 => "00010011",132 => "01101110",133 => "00100000",134 => "11100001",135 => "00011011",136 => "00000110",137 => "11001101",138 => "00100011",139 => "01000100",140 => "00000010",141 => "00111000",142 => "10010111",143 => "00010000",144 => "01100001",145 => "01100101",146 => "00110000",147 => "10101011",148 => "11110001",149 => "10010100",150 => "00100110",151 => "01011010",152 => "01101010",153 => "01111000",154 => "00011100",155 => "01101111",156 => "11111110",157 => "01110100",158 => "01110111",159 => "00100000",160 => "10011110",161 => "10011100",162 => "11100111",163 => "01100110",164 => "11111110",165 => "11000010",166 => "00010101",167 => "01011100",168 => "01110010",169 => "10111000",170 => "01111101",171 => "00000001",172 => "01010110",173 => "00101101",174 => "11000110",175 => "01010010",176 => "11100110",177 => "01010101",178 => "01000100",179 => "10000011",180 => "10111111",181 => "00110001",182 => "00101101",183 => "10000001",184 => "11001111",185 => "01011011",186 => "00110101",187 => "11101000",188 => "11101000",189 => "00100001",190 => "10001001",191 => "11111110",192 => "00011011",193 => "00000101",194 => "01000101",195 => "00000000",196 => "10010101",197 => "11010000",198 => "10111111",199 => "00001110",200 => "10101100",201 => "00000000",202 => "10100000",203 => "10100101",204 => "00110111",205 => "01001010",206 => "01101100",207 => "00110100",208 => "01011010",209 => "11010011",210 => "11001110",211 => "11010100",212 => "00000101",213 => "00100000",214 => "01111101",215 => "11000111",216 => "01110001",217 => "01000011",218 => "01110001",219 => "11111010",220 => "01111111",221 => "11001000",222 => "11010111",223 => "11110001",224 => "10111000",225 => "00001111",226 => "01111110",227 => "10100111",228 => "11110101",229 => "01111111",230 => "10010001",231 => "01000100",232 => "10110101",233 => "10110011",234 => "00111001",235 => "11010100",236 => "11000001",237 => "01100010",238 => "10100100",239 => "11111011",240 => "11110010",241 => "01010110",242 => "00010010",243 => "10001110",244 => "11110011",245 => "11001101",246 => "00010100",247 => "01001011",248 => "11010001",249 => "11101011",250 => "01110110",251 => "01101011",252 => "11001011",253 => "11000110",254 => "10110010",255 => "11100011",256 => "10100001",257 => "11101010",258 => "11100000",259 => "10000101",260 => "10111111",261 => "10110000",262 => "01110010",263 => "00100010",264 => "11111101",265 => "11111001",266 => "00000001",267 => "11101000",268 => "10011111",269 => "10001011",270 => "00000000",271 => "01000101",272 => "11110101",273 => "01001000",274 => "10000101",275 => "11100000",276 => "01111110",277 => "11011010",278 => "00101000",279 => "10010100",280 => "00101110",281 => "10111100",282 => "11101110",283 => "11111010",284 => "01010010",285 => "00101100",286 => "01111110",287 => "10110110",288 => "00011100",289 => "00000000",290 => "11100011",291 => "11001111",292 => "10001000",293 => "01001010",294 => "00011101",295 => "10011111",296 => "10111111",297 => "01101101",298 => "00000110",299 => "01010001",300 => "00010001",301 => "00110000",302 => "00001011",303 => "00101010",304 => "10110001",305 => "10001110",306 => "11111000",307 => "00100000",308 => "10111011",309 => "11101110",310 => "01010011",311 => "11110001",312 => "10000110",313 => "11111011",314 => "00111001",315 => "10001011",316 => "10100001",317 => "00011110",318 => "01110110",319 => "00011111",320 => "01000010",321 => "01010001",322 => "11100101",323 => "10011100",324 => "10011110",325 => "10000101",326 => "00011110",327 => "11110111",328 => "01111100",329 => "01111010",330 => "01111010",331 => "11010110",332 => "01110101",333 => "00101010",334 => "11101011",335 => "00011000",336 => "00111011",337 => "11010001",338 => "01011011",339 => "00001110",340 => "11011010",341 => "00111110",342 => "10001111",343 => "01011011",344 => "01101001",345 => "00110111",346 => "00100110",347 => "10000100",348 => "10001001",349 => "10111110",350 => "11100110",351 => "01100001",352 => "01100011",353 => "01010101",354 => "01101101",355 => "01100101",356 => "01000101",357 => "11001000",358 => "10110110",359 => "00001100",360 => "00100110",361 => "00101010",362 => "00100001",363 => "11101101",364 => "10010100",365 => "00100001",366 => "01110010",367 => "01000101",368 => "00000011",369 => "00010011",370 => "01010000",371 => "01110111",372 => "01110100",373 => "00101001",374 => "11100100",375 => "00010001",376 => "01001001",377 => "10110111",378 => "10110111",379 => "11100010",380 => "10011101",381 => "11100101",382 => "11001100",383 => "01110011",384 => "01110110",385 => "11001100",386 => "11000011",387 => "01001100",388 => "00110000",389 => "00110010",390 => "01111001",391 => "10011110",392 => "10001000",393 => "11011110",394 => "11010000",395 => "00000101",396 => "00010110",397 => "01001000",398 => "11100110",399 => "00110100",400 => "10101100",401 => "11010111",402 => "01111011",403 => "00100000",404 => "10100101",405 => "01010110",406 => "00001010",407 => "11110000",408 => "00001011",409 => "01010101",410 => "00110101",411 => "00100111",412 => "10001001",413 => "11011110",414 => "01110001",415 => "10100111",416 => "11000011",417 => "01001010",418 => "10110001",419 => "00101000",420 => "11111111",421 => "10100110",422 => "10101010",423 => "01110000",424 => "11011000",425 => "00111010",426 => "11110101",427 => "00111111",428 => "01110111",429 => "10100100",430 => "01001011",431 => "11110110",432 => "11100001",433 => "00000011",434 => "00100100",435 => "00101001",436 => "00000011",437 => "11001101",438 => "01000111",439 => "00100000",440 => "11010110",441 => "10100101",442 => "01111110",443 => "11100000",444 => "01010000",445 => "10101101",446 => "00010110",447 => "01101000",448 => "11100100",449 => "10110000",450 => "01110010",451 => "00100100",452 => "00101010",453 => "10010001",454 => "01111001",455 => "11111101",456 => "00111011",457 => "10110010",458 => "11000011",459 => "11011100",460 => "11000111",461 => "01011111",462 => "01111011",463 => "11010011",464 => "01110000",465 => "10110001",466 => "11111000",467 => "00010010",468 => "00011010",469 => "01100010",470 => "10001010",471 => "01101101",472 => "01000111",473 => "00111110",474 => "10110100",475 => "11111110",476 => "00011001",477 => "11101010",478 => "00111000",479 => "11001011",480 => "00111101",481 => "01101001",482 => "11110001",483 => "00100100",484 => "00011111",485 => "00001110",486 => "11011010",487 => "10111100",488 => "10000110",489 => "11101010",490 => "11100011",491 => "10001011",492 => "01000111",493 => "00101110",494 => "00011100",495 => "00011100",496 => "11101110",497 => "11100111",498 => "11000101",499 => "00101000",500 => "10000001",501 => "10011001",502 => "11001010",503 => "01101101",504 => "11010100",505 => "01000110",506 => "01100001",507 => "00000111",508 => "10111110",509 => "01100100",510 => "01000001",511 => "10000111",512 => "01011110",513 => "00000100",514 => "00100001",515 => "01010011",516 => "10101101",517 => "01001111",518 => "11100100",519 => "01110010",520 => "01100001",521 => "10110011",522 => "00110101",523 => "01010110",524 => "01010110",525 => "01111011",526 => "01001001",527 => "01111111",528 => "10000111",529 => "10110110",530 => "10000110",531 => "01000101",532 => "00100010",533 => "10010000",534 => "00001011",535 => "10010110",536 => "10011110",537 => "00001000",538 => "00111011",539 => "11001110",540 => "10101000",541 => "01000001",542 => "10010100",543 => "10001101",544 => "11011111",545 => "01100100",546 => "00100000",547 => "10010100",548 => "10111111",549 => "00101110",550 => "01110110",551 => "01000001",552 => "01111100",553 => "11001100",554 => "11110000",555 => "01100010",556 => "01100010",557 => "10101111",558 => "11011111",559 => "10101110",560 => "10000110",561 => "10111001",562 => "01110100",563 => "11001011",564 => "00010001",565 => "00111000",566 => "11101011",567 => "00111101",568 => "01011111",569 => "10000101",570 => "01110111",571 => "11011000",572 => "00011001",573 => "11001010",574 => "01101101",575 => "10100110",576 => "10101000",577 => "11100111",578 => "00100011",579 => "11101010",580 => "11101110",581 => "00000000",582 => "00110010",583 => "01001101",584 => "00100000",585 => "00011010",586 => "10000001",587 => "11010011",588 => "11001110",589 => "11011010",590 => "11110100",591 => "00011110",592 => "01011011",593 => "11010001",594 => "01100000",595 => "00111010",596 => "11100101",597 => "11000011",598 => "01110000",599 => "10000110",600 => "11000001",601 => "00100001",602 => "01111100",603 => "00010000",604 => "11100011",605 => "00101111",606 => "00001101",607 => "00101010",608 => "00101110",609 => "10100001",610 => "11001000",611 => "11100100",612 => "00101101",613 => "01111111",614 => "10111110",615 => "10011000",616 => "11000110",617 => "00010100",618 => "10011100",619 => "01000011",620 => "00111101",621 => "11101000",622 => "00110000",623 => "01110100",624 => "00000001",625 => "10110101",626 => "10010000",627 => "00100001",628 => "00101011",629 => "01011101",630 => "11101001",631 => "00100011",632 => "10011000",633 => "11100110",634 => "11000100",635 => "01011100",636 => "00101001",637 => "00100000",638 => "10000000",639 => "10001000",640 => "11010011",641 => "01111011",642 => "01100010",643 => "11010101",644 => "11101011",645 => "00000110",646 => "00110111",647 => "11011100",648 => "10111111",649 => "11110000",650 => "00100011",651 => "01111101",652 => "00111000",653 => "10011110",654 => "10001101",655 => "11111111",656 => "10101111",657 => "00100001",658 => "00110000",659 => "01111101",660 => "01111110",661 => "01000001",662 => "10000001",663 => "10010101",664 => "10111100",665 => "01111000",666 => "10000000",667 => "10011000",668 => "01010101",669 => "00011001",670 => "10000010",671 => "00011010",672 => "01101011",673 => "10001001",674 => "01001101",675 => "10100001",676 => "11110110",677 => "10000000",678 => "10100101",679 => "10010101",680 => "10100010",681 => "00111110",682 => "10100110",683 => "11001111",684 => "11001100",685 => "00110001",686 => "10100110",687 => "11000101",688 => "01110011",689 => "01111101",690 => "01111010",691 => "11011110",692 => "10011000",693 => "00110101",694 => "11010111",695 => "10000001",696 => "10001011",697 => "01000011",698 => "01011011",699 => "01000010",700 => "10000101",701 => "11010111",702 => "01110101",703 => "00100101",704 => "00111111",705 => "10010011",706 => "11010101",707 => "00100001",708 => "01111101",709 => "11101010",710 => "01100101",711 => "11101011",712 => "01101001",713 => "10011100",714 => "11101101",715 => "00010110",716 => "10111011",717 => "01000011",718 => "11001001",719 => "01111011",720 => "11100110",721 => "10000100",722 => "00101001",723 => "10000011",724 => "11011110",725 => "00100101",726 => "01101010",727 => "10101111",728 => "10110011",729 => "10101001",730 => "11001111",731 => "10001011",732 => "10011101",733 => "10010010",734 => "01110110",735 => "00010100",736 => "00100001",737 => "00110010",738 => "01110010",739 => "01100111",740 => "01010101",741 => "00101101",742 => "00001110",743 => "10010010",744 => "01111110",745 => "01101111",746 => "10100100",747 => "10001000",748 => "11001000",749 => "01101001",750 => "11110100",751 => "00101010",752 => "00101011",753 => "11100001",754 => "10001001",755 => "10001011",756 => "10000101",757 => "01110110",758 => "10101011",759 => "11110111",760 => "10100110",761 => "01111001",762 => "10010010",763 => "00010011",764 => "00110111",765 => "11000110",766 => "01110101",767 => "00010101",768 => "00110010",769 => "10001101",770 => "01000011",771 => "01001000",772 => "11101000",773 => "01011011",774 => "10111100",775 => "01101101",776 => "11010101",777 => "10101010",778 => "11011110",779 => "01110001",780 => "11110010",781 => "01111101",782 => "10110010",783 => "10001111",784 => "01010001",785 => "11010011",786 => "01010110",787 => "01100011",788 => "10100001",789 => "11011100",790 => "11111101",791 => "10011111",792 => "11111010",793 => "11110011",794 => "00010011",795 => "11100100",796 => "11100101",797 => "00101111",798 => "01011011",799 => "00001011",800 => "00100101",801 => "00010100",802 => "00000111",803 => "10101100",804 => "00110001",805 => "11110010",806 => "10100100",807 => "11100001",808 => "11110110",809 => "11011101",810 => "00111111",811 => "10110010",812 => "00011011",813 => "11011111",814 => "10011000",815 => "10111111",816 => "01010110",817 => "01110011",818 => "11110100",819 => "01101100",820 => "01010110",821 => "11111110",822 => "11000010",823 => "11110101",824 => "10111000",825 => "11010111",826 => "01111110",827 => "11111101",828 => "00111111",829 => "01011111",830 => "11100000",831 => "01111001",832 => "10010100",833 => "11110000",834 => "11111001",835 => "11101110",836 => "01011111",837 => "01100000",838 => "00100011",839 => "01110100",840 => "11111010",841 => "11000111",842 => "01011010",843 => "00001001",844 => "10111011",845 => "10000101",846 => "01010111",847 => "10011110",848 => "00111110",849 => "11001101",850 => "11110101",851 => "00011111",852 => "01001101",853 => "10111001",854 => "11101000",855 => "10011100",856 => "00111010",857 => "00101111",858 => "11001110",859 => "11000110",860 => "11111110",861 => "01011001",862 => "10101011",863 => "11010010",864 => "01001100",865 => "01110100",866 => "10010111",867 => "10110001",868 => "10001100",869 => "01101011",870 => "01111110",871 => "10100000",872 => "00010110",873 => "01001011",874 => "00011011",875 => "00010101",876 => "11001011",877 => "00011001",878 => "10101001",879 => "01110100",880 => "11111110",881 => "01001110",882 => "00011010",883 => "10100011",884 => "00010100",885 => "10110100",886 => "00010010",887 => "10001101",888 => "01001011",889 => "10010110",890 => "11011010",891 => "01001001",892 => "10100000",893 => "11111110",894 => "01001010",895 => "11110100",896 => "00111101",897 => "10001010",898 => "00111000",899 => "11100011",900 => "01000111",901 => "11101101",902 => "01000100",903 => "01110110",904 => "11111111",905 => "10110111",906 => "11010111",907 => "10111001",908 => "11100010",909 => "11110000",910 => "00000111",911 => "00111110",912 => "11101101",913 => "00001010",914 => "11111101",915 => "01011101",916 => "00100000",917 => "00101101",918 => "01110100",919 => "10100100",920 => "11110001",921 => "01101001",922 => "11110001",923 => "11000001",924 => "00010101",925 => "01000100",926 => "01000001",927 => "11100101",928 => "00111011",929 => "00101110",930 => "00101011",931 => "01011010",932 => "11010110",933 => "10000111",934 => "00110011",935 => "01110100",936 => "01110101",937 => "10111000",938 => "00000011",939 => "11011110",940 => "01101010",941 => "10100010",942 => "11100010",943 => "10001001",944 => "01110000",945 => "10110011",946 => "01110101",947 => "01010100",948 => "00110011",949 => "10000000",950 => "01011101",951 => "00110101",952 => "11110010",953 => "10101100",954 => "11000000",955 => "00111001",956 => "00001111",957 => "11111101",958 => "01000101",959 => "10010001",960 => "11010011",961 => "01001001",962 => "10111111",963 => "00000110",964 => "10111010",965 => "10010101",966 => "00100101",967 => "11001011",968 => "00111110",969 => "01000101",970 => "10101110",971 => "11000011",972 => "10001101",973 => "11011100",974 => "11111000",975 => "00110100",976 => "01111001",977 => "10010010",978 => "00011111",979 => "10001101",980 => "10100110",981 => "11001010",982 => "01010111",983 => "01101110",984 => "11001100",985 => "11000100",986 => "01000011",987 => "11111011",988 => "10111111",989 => "01011101",990 => "10001011",991 => "11011101",992 => "01011000",993 => "10100010",994 => "10111010",995 => "11111011",996 => "01010100",997 => "00000000",998 => "11100110",999 => "11101111",1000 => "01110011",1001 => "00110010",1002 => "00010001",1003 => "11100100",1004 => "11011000",1005 => "01100110",1006 => "00100001",1007 => "10111011",1008 => "11010100",1009 => "01101100",1010 => "01001010",1011 => "10000010",1012 => "01000100",1013 => "10101001",1014 => "01100001",1015 => "11110111",1016 => "00101100",1017 => "11011011",1018 => "00010111",1019 => "00001010",1020 => "00000111",1021 => "00100001",1022 => "11100101",1023 => "11110111",1024 => "01001001",1025 => "01011110",1026 => "10000000",1027 => "01001010",1028 => "11110010",1029 => "11111011",1030 => "01100100",1031 => "10011001",1032 => "10111111",1033 => "00100001",1034 => "00011110",1035 => "10100010",1036 => "10110011",1037 => "10111110",1038 => "10100110",1039 => "00011111",1040 => "01011111",1041 => "01010101",1042 => "11111111",1043 => "01111110",1044 => "00001110",1045 => "00011011",1046 => "11110111",1047 => "11011010",1048 => "11101110",1049 => "11011010",1050 => "11001000",1051 => "00101010",1052 => "01011101",1053 => "00000101",1054 => "01011101",1055 => "10011111",1056 => "10100001",1057 => "01001011",1058 => "01111110",1059 => "00000000",1060 => "11000110",1061 => "01111111",1062 => "01001111",1063 => "11100011",1064 => "10101110",1065 => "11101000",1066 => "00001001",1067 => "00110001",1068 => "11101001",1069 => "00110100",1070 => "11111111",1071 => "00001010",1072 => "10011111",1073 => "11000110",1074 => "10100011",1075 => "00111000",1076 => "00101011",1077 => "00101100",1078 => "11001010",1079 => "10010001",1080 => "01000110",1081 => "10100111",1082 => "10001011",1083 => "01010011",1084 => "10111100",1085 => "00101000",1086 => "01010110",1087 => "11011010",1088 => "10001111",1089 => "01011110",1090 => "10000001",1091 => "10001110",1092 => "01111010",1093 => "01001000",1094 => "01101001",1095 => "11001111",1096 => "10001110",1097 => "00010011",1098 => "01011100",1099 => "01111101",1100 => "01000011",1101 => "11001101",1102 => "11100011",1103 => "11101011",1104 => "11001000",1105 => "10111110",1106 => "11111110",1107 => "01101011",1108 => "11000010",1109 => "10000111",1110 => "11100001",1111 => "01011100",1112 => "10110101",1113 => "01010101",1114 => "01001100",1115 => "10101111",1116 => "10101110",1117 => "00101010",1118 => "10001011",1119 => "11110100",1120 => "11110111",1121 => "01110000",1122 => "11101011",1123 => "11110100",1124 => "10000100",1125 => "11100000",1126 => "11000110",1127 => "10111100",1128 => "01010111",1129 => "11000110",1130 => "10010001",1131 => "01101111",1132 => "11100111",1133 => "11011000",1134 => "00011010",1135 => "10101100",1136 => "11111011",1137 => "11011010",1138 => "10011100",1139 => "10001110",1140 => "00000000",1141 => "00010000",1142 => "11000111",1143 => "01110101",1144 => "11000110",1145 => "01000111",1146 => "00110111",1147 => "01011110",1148 => "11100110",1149 => "10111010",1150 => "10101110",1151 => "11010101",1152 => "10101011",1153 => "10100010",1154 => "10001010",1155 => "01011111",1156 => "00101011",1157 => "11011011",1158 => "00001100",1159 => "11100001",1160 => "01001111",1161 => "11000110",1162 => "10010011",1163 => "00110001",1164 => "11000001",1165 => "00001100",1166 => "00000101",1167 => "01001111",1168 => "10010100",1169 => "00011111",1170 => "10000001",1171 => "10001000",1172 => "00100101",1173 => "00000100",1174 => "11100010",1175 => "01011100",1176 => "01111101",1177 => "11010001",1178 => "10101010",1179 => "11001110",1180 => "10011101",1181 => "11100100",1182 => "01111100",1183 => "00111010",1184 => "00001010",1185 => "11100010",1186 => "11100100",1187 => "10011100",1188 => "10010000",1189 => "00100011",1190 => "00100010",1191 => "10101100",1192 => "11010111",1193 => "10001110",1194 => "00101011",1195 => "11100100",1196 => "01100000",1197 => "01100010",1198 => "11001101",1199 => "01111101",1200 => "01110100",1201 => "01010111",1202 => "01101000",1203 => "11101011",1204 => "10101011",1205 => "11011010",1206 => "01011000",1207 => "00011100",1208 => "11100110",1209 => "11010011",1210 => "01001101",1211 => "01100011",1212 => "01111010",1213 => "10001100",1214 => "01000110",1215 => "01010110",1216 => "11111001",1217 => "11101011",1218 => "00011101",1219 => "01000110",1220 => "01001011",1221 => "01100011",1222 => "10111101",1223 => "01111101",1224 => "01101000",1225 => "01110101",1226 => "00111111",1227 => "11011010",1228 => "10010101",1229 => "11010000",1230 => "00001000",1231 => "01010110",1232 => "00110100",1233 => "11101100",1234 => "01110000",1235 => "00101010",1236 => "01101000",1237 => "10010001",1238 => "01100110",1239 => "10110001",1240 => "01110101",1241 => "10100110",1242 => "11100101",1243 => "10111110",1244 => "01011001",1245 => "01010111",1246 => "01101011",1247 => "10110111",1248 => "01010111",1249 => "10111111",1250 => "10111110",1251 => "10100011",1252 => "11010101",1253 => "10100000",1254 => "11000110",1255 => "11010100",1256 => "11110000",1257 => "00100111",1258 => "00111010",1259 => "00111111",1260 => "11111011",1261 => "11100101",1262 => "00100000",1263 => "01000101",1264 => "10101000",1265 => "00011110",1266 => "00111011",1267 => "00101001",1268 => "00101111",1269 => "11111010",1270 => "01111001",1271 => "01100000",1272 => "10010010",1273 => "11010011",1274 => "00010000",1275 => "01101111",1276 => "10011110",1277 => "10110001",1278 => "01110110",1279 => "01110001",1280 => "01110111",1281 => "11011111",1282 => "01011110",1283 => "11111111",1284 => "00011000",1285 => "11100001",1286 => "01111110",1287 => "00100100",1288 => "10001000",1289 => "11010000",1290 => "10110010",1291 => "00010110",1292 => "00011001",1293 => "00111011",1294 => "00110100",1295 => "10011001",1296 => "00001101",1297 => "11110000",1298 => "10110101",1299 => "11000111",1300 => "01100100",1301 => "01010111",1302 => "00010110",1303 => "01000010",1304 => "00010001",1305 => "11111011",1306 => "00011101",1307 => "00010001",1308 => "10100110",1309 => "11001001",1310 => "11100011",1311 => "00001110",1312 => "11001001",1313 => "10111101",1314 => "01111001",1315 => "10011011",1316 => "11011100",1317 => "10000000",1318 => "11001000",1319 => "00011010",1320 => "00000000",1321 => "11010011",1322 => "00001010",1323 => "10011000",1324 => "01011101",1325 => "00100111",1326 => "01000110",1327 => "00111100",1328 => "00110011",1329 => "10111100",1330 => "00100101",1331 => "10110110",1332 => "11000011",1333 => "01010101",1334 => "10101111",1335 => "11010011",1336 => "11010110",1337 => "00111110",1338 => "10011001",1339 => "11010000",1340 => "11000100",1341 => "00110100",1342 => "00000001",1343 => "00001111",1344 => "00010001",1345 => "01010011",1346 => "01011001",1347 => "11100000",1348 => "00110111",1349 => "00011101",1350 => "11110100",1351 => "00000001",1352 => "01001100",1353 => "10001111",1354 => "00101000",1355 => "00011101",1356 => "10000011",1357 => "11010010",1358 => "10000101",1359 => "10100101",1360 => "10001000",1361 => "10101111",1362 => "00011010",1363 => "11110110",1364 => "11010100",1365 => "01100111",1366 => "01010111",1367 => "01110110",1368 => "11110111",1369 => "11110011",1370 => "01001100",1371 => "01111111",1372 => "11011100",1373 => "11011111",1374 => "10010111",1375 => "01010111",1376 => "10110110",1377 => "00100110",1378 => "11010011",1379 => "00101000",1380 => "00110110",1381 => "01000110",1382 => "01000111",1383 => "01010001",1384 => "00011111",1385 => "11000001",1386 => "01011110",1387 => "01101101",1388 => "00110110",1389 => "00001101",1390 => "01011000",1391 => "01010011",1392 => "11001011",1393 => "11010000",1394 => "11001100",1395 => "00100010",1396 => "01111101",1397 => "11001011",1398 => "00000101",1399 => "01101100",1400 => "10111111",1401 => "00101010",1402 => "10010010",1403 => "10011010",1404 => "01011101",1405 => "00111111",1406 => "10010000",1407 => "11100101",1408 => "00100010",1409 => "11000100",1410 => "11010011",1411 => "00100101",1412 => "01011000",1413 => "11011110",1414 => "01100000",1415 => "01000011",1416 => "10111010",1417 => "00111000",1418 => "10000110",1419 => "01011000",1420 => "00000111",1421 => "01100101",1422 => "10000010",1423 => "00010100",1424 => "01100101",1425 => "00101000",1426 => "01101101",1427 => "10010000",1428 => "10111101",1429 => "00001011",1430 => "10011100",1431 => "00010101",1432 => "00100110",1433 => "10001110",1434 => "10010101",1435 => "00000000",1436 => "11101010",1437 => "11000010",1438 => "11110101",1439 => "10001011",1440 => "10101111",1441 => "11111101",1442 => "01001110",1443 => "01110010",1444 => "10001101",1445 => "11001010",1446 => "10011100",1447 => "10001000",1448 => "11010011",1449 => "01001001",1450 => "00111001",1451 => "11010011",1452 => "01010001",1453 => "00010100",1454 => "00111110",1455 => "01001111",1456 => "00100101",1457 => "00001001",1458 => "01001011",1459 => "00010100",1460 => "01110000",1461 => "01111010",1462 => "10101011",1463 => "01111111",1464 => "10010000",1465 => "00101100",1466 => "10100101",1467 => "00000101",1468 => "00111001",1469 => "10000101",1470 => "11000111",1471 => "11000111",1472 => "00110011",1473 => "00001001",1474 => "01100110",1475 => "01110001",1476 => "01111001",1477 => "10111111",1478 => "01010100",1479 => "01010000",1480 => "10010111",1481 => "00101011",1482 => "10001010",1483 => "01101101",1484 => "01100000",1485 => "11010000",1486 => "01010111",1487 => "00100001",1488 => "01110000",1489 => "01010010",1490 => "00110001",1491 => "01100110",1492 => "10010101",1493 => "10100001",1494 => "10000101",1495 => "00001001",1496 => "00100111",1497 => "10010011",1498 => "10011010",1499 => "11011111",1500 => "00110111",1501 => "00101100",1502 => "01000010",1503 => "11101000",1504 => "11000100",1505 => "10000000",1506 => "10010000",1507 => "00101010",1508 => "11110110",1509 => "00100010",1510 => "01110010",1511 => "10001100",1512 => "10010011",1513 => "10010011",1514 => "11001110",1515 => "11010011",1516 => "00110110",1517 => "10001100",1518 => "10100001",1519 => "10001100",1520 => "11000011",1521 => "01001100",1522 => "00011001",1523 => "00010100",1524 => "10101000",1525 => "01000010",1526 => "11001011",1527 => "01100110",1528 => "10110110",1529 => "01000111",1530 => "10010110",1531 => "01000011",1532 => "11111010",1533 => "11010101",1534 => "01110100",1535 => "01100110",1536 => "11111010",1537 => "10101100",1538 => "10000010",1539 => "01011000",1540 => "00110101",1541 => "01100101",1542 => "11111010",1543 => "10111101",1544 => "01111111",1545 => "10101111",1546 => "11101010",1547 => "10110010",1548 => "00001011",1549 => "11110000",1550 => "01010100",1551 => "01011110",1552 => "00010111",1553 => "10011001",1554 => "01111101",1555 => "00100111",1556 => "00010011",1557 => "00000011",1558 => "11101001",1559 => "00000110",1560 => "01010110",1561 => "00010011",1562 => "01000001",1563 => "11111010",1564 => "00100011",1565 => "11000010",1566 => "10011110",1567 => "10000111",1568 => "00010101",1569 => "01101000",1570 => "10001001",1571 => "01011110",1572 => "01001110",1573 => "00000110",1574 => "11001101",1575 => "10111000",1576 => "00101111",1577 => "11100101",1578 => "00101011",1579 => "00001110",1580 => "10100011",1581 => "10010111",1582 => "00100101",1583 => "01001001",1584 => "00101100",1585 => "01010010",1586 => "00010110",1587 => "01001111",1588 => "11000100",1589 => "10011101",1590 => "00010011",1591 => "01111101",1592 => "00111101",1593 => "00111001",1594 => "10110010",1595 => "00100101",1596 => "10100011",1597 => "01100001",1598 => "00010111",1599 => "01001111",1600 => "10011010",1601 => "11010101",1602 => "01111110",1603 => "11010000",1604 => "10100000",1605 => "11001100",1606 => "11000000",1607 => "11000100",1608 => "00110001",1609 => "11011001",1610 => "10000110",1611 => "10110110",1612 => "01011001",1613 => "10000111",1614 => "01001010",1615 => "11101000",1616 => "11000001",1617 => "00001101",1618 => "10010100",1619 => "00101101",1620 => "00111111",1621 => "01111110",1622 => "11011111",1623 => "00011101",1624 => "11111110",1625 => "01111101",1626 => "01010100",1627 => "11100111",1628 => "01100011",1629 => "00101111",1630 => "10110000",1631 => "10111001",1632 => "01011000",1633 => "11101110",1634 => "10110101",1635 => "00011111",1636 => "01100100",1637 => "11101000",1638 => "00101001",1639 => "10111001",1640 => "00010111",1641 => "11100010",1642 => "01010110",1643 => "11010111",1644 => "10000011",1645 => "10111110",1646 => "00011110",1647 => "00100111",1648 => "00110101",1649 => "10010000",1650 => "10011101",1651 => "11111100",1652 => "01011010",1653 => "00001111",1654 => "10010011",1655 => "01011010",1656 => "01001100",1657 => "00100111",1658 => "10010101",1659 => "10101000",1660 => "01011101",1661 => "00000111",1662 => "10111111",1663 => "11101001",1664 => "01111111",1665 => "00010000",1666 => "11000101",1667 => "10000101",1668 => "11010010",1669 => "01010010",1670 => "11001101",1671 => "11001011",1672 => "10001100",1673 => "00110110",1674 => "01110001",1675 => "01010011",1676 => "00000100",1677 => "10000010",1678 => "10111110",1679 => "10111011",1680 => "00010001",1681 => "01000100",1682 => "00001000",1683 => "01000000",1684 => "01111000",1685 => "11101101",1686 => "10001010",1687 => "00110001",1688 => "01100000",1689 => "01100101",1690 => "01110000",1691 => "10010010",1692 => "10010001",1693 => "00011001",1694 => "01011000",1695 => "00011000",1696 => "11111100",1697 => "00110101",1698 => "00100110",1699 => "10100100",1700 => "00100000",1701 => "01101010",1702 => "00001110",1703 => "10110100",1704 => "01110100",1705 => "10011010",1706 => "10110101",1707 => "11011000",1708 => "10100001",1709 => "01001001",1710 => "10011110",1711 => "01111011",1712 => "01111001",1713 => "11001000",1714 => "00010010",1715 => "11001101",1716 => "01101010",1717 => "01001111",1718 => "00111101",1719 => "01000111",1720 => "01011110",1721 => "10111100",1722 => "11000100",1723 => "00110111",1724 => "00001101",1725 => "01101110",1726 => "01011000",1727 => "00101111",1728 => "01110000",1729 => "11100011",1730 => "01101010",1731 => "01100011",1732 => "10111100",1733 => "01000100",1734 => "01111110",1735 => "01111110",1736 => "01010001",1737 => "00010100",1738 => "11110111",1739 => "10011010",1740 => "01110001",1741 => "10000101",1742 => "00101110",1743 => "10010001",1744 => "01010110",1745 => "00101101",1746 => "10010010",1747 => "01000111",1748 => "00101001",1749 => "11101011",1750 => "00010100",1751 => "01100000",1752 => "01001000",1753 => "11111011",1754 => "01101001",1755 => "10000011",1756 => "01110001",1757 => "10010101",1758 => "01010011",1759 => "01010101",1760 => "01111000",1761 => "10101111",1762 => "00101111",1763 => "10000011",1764 => "01001100",1765 => "00111001",1766 => "01011101",1767 => "00010010",1768 => "01101111",1769 => "01100010",1770 => "00101110",1771 => "00101010",1772 => "00000111",1773 => "10100011",1774 => "11100011",1775 => "00001111",1776 => "01110100",1777 => "01111000",1778 => "10100110",1779 => "11111000",1780 => "00100110",1781 => "00100010",1782 => "11010110",1783 => "00001010",1784 => "00100100",1785 => "11001011",1786 => "01010010",1787 => "11111101",1788 => "01000010",1789 => "00011110",1790 => "11110011",1791 => "10100001",1792 => "10101011",1793 => "00001010",1794 => "00111111",1795 => "00101110",1796 => "01000101",1797 => "00001110",1798 => "10110111",1799 => "01011101",1800 => "11001101",1801 => "11010101",1802 => "01101011",1803 => "10100111",1804 => "10110111",1805 => "01111111",1806 => "10100110",1807 => "00100010",1808 => "00001010",1809 => "10010010",1810 => "10001111",1811 => "10011100",1812 => "00011101",1813 => "00001101",1814 => "11100000",1815 => "10010110",1816 => "01100101",1817 => "00111001",1818 => "00110100",1819 => "00101100",1820 => "01010101",1821 => "01101100",1822 => "10111000",1823 => "00110001",1824 => "11000110",1825 => "01110100",1826 => "10101100",1827 => "01001100",1828 => "01001000",1829 => "01100000",1830 => "10000111",1831 => "00100000",1832 => "11001101",1833 => "01001001",1834 => "10000110",1835 => "01100110",1836 => "11101111",1837 => "10001011",1838 => "00111101",1839 => "11111011",1840 => "01010001",1841 => "11000011",1842 => "11001101",1843 => "10100010",1844 => "11000101",1845 => "00010000",1846 => "10111010",1847 => "10000011",1848 => "01111111",1849 => "11010001",1850 => "10010000",1851 => "01100000",1852 => "10011011",1853 => "10100110",1854 => "11011111",1855 => "01001010",1856 => "00011000",1857 => "11000011",1858 => "00100100",1859 => "01010101",1860 => "11110000",1861 => "10001110",1862 => "01111100",1863 => "00001101",1864 => "00110011",1865 => "01011101",1866 => "10101111",1867 => "01011110",1868 => "10101110",1869 => "01001001",1870 => "11001110",1871 => "10111001",1872 => "00110110",1873 => "01101000",1874 => "10000111",1875 => "11011010",1876 => "11110101",1877 => "11000101",1878 => "10010111",1879 => "01011110",1880 => "01011011",1881 => "11010000",1882 => "00101011",1883 => "01001000",1884 => "11001010",1885 => "01011011",1886 => "10001011",1887 => "10011010",1888 => "11100000",1889 => "11101111",1890 => "00001010",1891 => "11010010",1892 => "01101001",1893 => "11101001",1894 => "01101010",1895 => "11000101",1896 => "10111111",1897 => "11101111",1898 => "01010010",1899 => "10111010",1900 => "10010101",1901 => "10111100",1902 => "01111010",1903 => "11111001",1904 => "00100000",1905 => "00001101",1906 => "00110001",1907 => "01000011",1908 => "11101111",1909 => "10111101",1910 => "10010000",1911 => "11010111",1912 => "11001000",1913 => "11100111",1914 => "01011101",1915 => "00010011",1916 => "01110111",1917 => "10000101",1918 => "10101000",1919 => "10010110",1920 => "01111001",1921 => "10110010",1922 => "11101000",1923 => "10101001",1924 => "00111100",1925 => "11100010",1926 => "00011010",1927 => "01101101",1928 => "00100010",1929 => "11001000",1930 => "01010110",1931 => "10011010",1932 => "01000101",1933 => "11111001",1934 => "01001000",1935 => "11111001",1936 => "10000010",1937 => "10111011",1938 => "01100110",1939 => "01110000",1940 => "01010111",1941 => "10101101",1942 => "00100110",1943 => "00000001",1944 => "10000000",1945 => "00011011",1946 => "11000001",1947 => "01101000",1948 => "11101011",1949 => "10111000",1950 => "00100010",1951 => "10110100",1952 => "01000010",1953 => "10111101",1954 => "01011111",1955 => "10110111",1956 => "11110100",1957 => "10011001",1958 => "01101111",1959 => "00101011",1960 => "01100100",1961 => "00000011",1962 => "10110010",1963 => "10010111",1964 => "10111100",1965 => "00101000",1966 => "11101101",1967 => "11110100",1968 => "01000010",1969 => "01111010",1970 => "00101000",1971 => "00001000",1972 => "00001001",1973 => "00110000",1974 => "10111100",1975 => "00001000",1976 => "01101000",1977 => "00011111",1978 => "00011110",1979 => "10011110",1980 => "11000011",1981 => "11001101",1982 => "11100011",1983 => "11100001",1984 => "11101010",1985 => "10011111",1986 => "11010100",1987 => "11001010",1988 => "11100000",1989 => "10100000",1990 => "01111111",1991 => "10101101",1992 => "11111110",1993 => "00100000",1994 => "01010111",1995 => "11010001",1996 => "01010100",1997 => "10000000",1998 => "11101000",1999 => "10000110",2000 => "01001001",2001 => "00101011",2002 => "10010001",2003 => "10101110",2004 => "10110011",2005 => "00011010",2006 => "11111111",2007 => "00001110",2008 => "10000010",2009 => "01011101",2010 => "11101100",2011 => "10110010",2012 => "10100000",2013 => "00101111",2014 => "00110000",2015 => "00001101",2016 => "11001101",2017 => "10110101",2018 => "00111000",2019 => "11001010",2020 => "01111000",2021 => "10011010",2022 => "11101110",2023 => "11110110",2024 => "00001110",2025 => "01111011",2026 => "01100000",2027 => "00000011",2028 => "00100010",2029 => "01100100",2030 => "11011011",2031 => "01110100",2032 => "10010110",2033 => "00001001",2034 => "01110100",2035 => "01011100",2036 => "10100001",2037 => "11011101",2038 => "00100111",2039 => "10100000",2040 => "00111001",2041 => "11101010",2042 => "01100101",2043 => "00100000",2044 => "01001111",2045 => "11101101",2046 => "00000111",2047 => "10001111",2048 => "01100001",2049 => "11101100",2050 => "00000011",2051 => "01111111",2052 => "11001110",2053 => "01011001",2054 => "00101000",2055 => "01101100",2056 => "10010000",2057 => "11011101",2058 => "10101010",2059 => "01001010",2060 => "01101000",2061 => "00011101",2062 => "01111011",2063 => "10111011",2064 => "00011111",2065 => "11010001",2066 => "00110000",2067 => "11011010",2068 => "11101001",2069 => "01100001",2070 => "01010111",2071 => "11000100",2072 => "10110110",2073 => "11011110",2074 => "00100101",2075 => "00011110",2076 => "10001101",2077 => "10010001",2078 => "01101000",2079 => "00100010",2080 => "10101010",2081 => "01111100",2082 => "10000011",2083 => "00000100",2084 => "11111111",2085 => "11001101",2086 => "00100001",2087 => "11110100",2088 => "01110100",2089 => "01100101",2090 => "00000111",2091 => "01101111",2092 => "01111011",2093 => "00010110",2094 => "01101001",2095 => "00010001",2096 => "11101001",2097 => "01110100",2098 => "11011100",2099 => "00111111",2100 => "11010011",2101 => "10100000",2102 => "00000100",2103 => "11001111",2104 => "00101101",2105 => "10011111",2106 => "10110000",2107 => "01011001",2108 => "10110010",2109 => "01100000",2110 => "10101001",2111 => "00101011",2112 => "00111001",2113 => "11011100",2114 => "00001000",2115 => "01000111",2116 => "11111001",2117 => "11010000",2118 => "10001011",2119 => "11110111",2120 => "11000001",2121 => "10000110",2122 => "01010110",2123 => "00011101",2124 => "10111101",2125 => "01000100",2126 => "10010001",2127 => "11101101",2128 => "11100011",2129 => "10011111",2130 => "10001001",2131 => "10011100",2132 => "10101011",2133 => "11010101",2134 => "00010011",2135 => "11110011",2136 => "01111001",2137 => "00101110",2138 => "01101010",2139 => "01100000",2140 => "00101100",2141 => "00011101",2142 => "00000110",2143 => "10001100",2144 => "10111001",2145 => "10110000",2146 => "01010010",2147 => "10111010",2148 => "00010100",2149 => "01001100",2150 => "10000100",2151 => "11100110",2152 => "01000110",2153 => "01100011",2154 => "11011100",2155 => "00011110",2156 => "00000111",2157 => "10000011",2158 => "01011000",2159 => "00011001",2160 => "00111000",2161 => "01000101",2162 => "01010000",2163 => "00101001",2164 => "00100100",2165 => "01110011",2166 => "01100101",2167 => "10001100",2168 => "10010011",2169 => "10001100",2170 => "10001011",2171 => "00011001",2172 => "10011111",2173 => "10001000",2174 => "01000100",2175 => "11011001",2176 => "11001100",2177 => "10010011",2178 => "00010010",2179 => "11101001",2180 => "01010001",2181 => "10101101",2182 => "11100111",2183 => "11010010",2184 => "00001001",2185 => "10011011",2186 => "00000100",2187 => "00110011",2188 => "01100010",2189 => "01011101",2190 => "01010101",2191 => "01011000",2192 => "01101010",2193 => "11000101",2194 => "00000011",2195 => "01110100",2196 => "01110110",2197 => "01011011",2198 => "01100111",2199 => "10000101",2200 => "10111010",2201 => "01000110",2202 => "11001011",2203 => "11100101",2204 => "11000011",2205 => "11011110",2206 => "10110001",2207 => "11010011",2208 => "11011101",2209 => "10101100",2210 => "00100101",2211 => "10101101",2212 => "11001000",2213 => "11010001",2214 => "11000100",2215 => "01011101",2216 => "00111101",2217 => "11001001",2218 => "10000001",2219 => "11011010",2220 => "01100110",2221 => "00010110",2222 => "10011100",2223 => "00111001",2224 => "00100111",2225 => "01110101",2226 => "11000001",2227 => "10000001",2228 => "01101001",2229 => "00001111",2230 => "00111010",2231 => "11011001",2232 => "10111001",2233 => "10101101",2234 => "10101100",2235 => "11011001",2236 => "00111001",2237 => "01010001",2238 => "10000000",2239 => "00100000",2240 => "01100111",2241 => "01111000",2242 => "01101111",2243 => "10011110",2244 => "01001100",2245 => "11011001",2246 => "11101010",2247 => "11100011",2248 => "00100001",2249 => "11000110",2250 => "00000111",2251 => "11001111",2252 => "10011011",2253 => "01001000",2254 => "11010011",2255 => "01000010",2256 => "00100101",2257 => "10111011",2258 => "00000000",2259 => "00001110",2260 => "11100001",2261 => "01000111",2262 => "10100100",2263 => "00010111",2264 => "11100101",2265 => "10111101",2266 => "10010011",2267 => "01000000",2268 => "00011100",2269 => "01010001",2270 => "10110111",2271 => "01010110",2272 => "01001010",2273 => "10100001",2274 => "11011111",2275 => "10111000",2276 => "10111001",2277 => "00101011",2278 => "00010010",2279 => "00111110",2280 => "11100111",2281 => "10111101",2282 => "11101111",2283 => "10010111",2284 => "10100010",2285 => "00011000",2286 => "10000101",2287 => "01111101",2288 => "01010100",2289 => "00110010",2290 => "10001101",2291 => "10110011",2292 => "10011011",2293 => "10111111",2294 => "11101101",2295 => "10010011",2296 => "11101000",2297 => "11100010",2298 => "10011011",2299 => "11011111",2300 => "00000111",2301 => "00010011",2302 => "11001100",2303 => "01110010",2304 => "01111100",2305 => "11001101",2306 => "00101110",2307 => "00000000",2308 => "11111111",2309 => "00000110",2310 => "10000101",2311 => "10010011",2312 => "11001100",2313 => "10000111",2314 => "11100001",2315 => "01100010",2316 => "01010100",2317 => "00110001",2318 => "00111101",2319 => "10100001",2320 => "00011101",2321 => "10101010",2322 => "11110101",2323 => "01101101",2324 => "00110010",2325 => "10101010",2326 => "01001010",2327 => "10101011",2328 => "00101101",2329 => "01110000",2330 => "01010111",2331 => "11000111",2332 => "00111001",2333 => "01011101",2334 => "00100001",2335 => "01001101",2336 => "01110010",2337 => "11100000",2338 => "11001100",2339 => "11011101",2340 => "10011000",2341 => "10100010",2342 => "01010111",2343 => "00110001",2344 => "10001010",2345 => "00000111",2346 => "11110010",2347 => "10010000",2348 => "11110101",2349 => "11011000",2350 => "11000010",2351 => "01000110",2352 => "11000011",2353 => "10001110",2354 => "11111100",2355 => "11001110",2356 => "11100110",2357 => "01101110",2358 => "11110100",2359 => "11010011",2360 => "00110110",2361 => "10110101",2362 => "10001000",2363 => "10101110",2364 => "01010001",2365 => "01110101",2366 => "10101001",2367 => "01010101",2368 => "11101001",2369 => "00010111",2370 => "00001011",2371 => "11101100",2372 => "01100010",2373 => "10110110",2374 => "10111110",2375 => "10010001",2376 => "00010010",2377 => "11101001",2378 => "11101111",2379 => "00001000",2380 => "10111111",2381 => "10100000",2382 => "10101010",2383 => "01101111",2384 => "10100010",2385 => "01100110",2386 => "10010001",2387 => "00110010",2388 => "00101100",2389 => "01101101",2390 => "11011110",2391 => "01000010",2392 => "00010111",2393 => "10110001",2394 => "10000110",2395 => "10011100",2396 => "01010101",2397 => "00100111",2398 => "11110000",2399 => "11101111",2400 => "01000111",2401 => "00001110",2402 => "00011110",2403 => "11101001",2404 => "01001000",2405 => "01001111",2406 => "01000010",2407 => "00100010",2408 => "10101011",2409 => "10010100",2410 => "11100010",2411 => "00010011",2412 => "10010101",2413 => "11011011",2414 => "10011010",2415 => "01101111",2416 => "10100101",2417 => "10001101",2418 => "00001011",2419 => "01101101",2420 => "10111101",2421 => "11000010",2422 => "00110111",2423 => "00100111",2424 => "11111011",2425 => "01011110",2426 => "00000000",2427 => "10111101",2428 => "01010000",2429 => "11100110",2430 => "01100001",2431 => "00111001",2432 => "00110011",2433 => "11010001",2434 => "10011000",2435 => "11100111",2436 => "00110111",2437 => "11101101",2438 => "00101101",2439 => "01100000",2440 => "11000100",2441 => "00000110",2442 => "01001101",2443 => "00111011",2444 => "01100110",2445 => "00101010",2446 => "00001110",2447 => "10011110",2448 => "11110000",2449 => "01011010",2450 => "10000011",2451 => "11111101",2452 => "11100101",2453 => "11010001",2454 => "00000110",2455 => "11101011",2456 => "11110011",2457 => "00101100",2458 => "11100100",2459 => "11010100",2460 => "01100111",2461 => "01010011",2462 => "01010011",2463 => "11010110",2464 => "11011111",2465 => "11001111",2466 => "10101110",2467 => "01000011",2468 => "10110010",2469 => "11100011",2470 => "11011110",2471 => "01001110",2472 => "10110000",2473 => "11100101",2474 => "01010100",2475 => "00101110",2476 => "01111110",2477 => "10100100",2478 => "11001101",2479 => "10010010",2480 => "11100100",2481 => "00111101",2482 => "10011111",2483 => "00000110",2484 => "01000111",2485 => "11101110",2486 => "10111000",2487 => "11110011",2488 => "00110010",2489 => "10010101",2490 => "10110001",2491 => "01101001",2492 => "10011001",2493 => "00000110",2494 => "00000000",2495 => "10111010",2496 => "00011111",2497 => "10011101",2498 => "11101011",2499 => "11011101",2500 => "00001000",2501 => "10000111",2502 => "00011011",2503 => "10010101",2504 => "10010111",2505 => "11001111",2506 => "10010001",2507 => "01011111",2508 => "10111001",2509 => "11100001",2510 => "10001110",2511 => "00110111",2512 => "01111110",2513 => "01000001",2514 => "10011000",2515 => "01100000",2516 => "10011101",2517 => "00110011",2518 => "01001111",2519 => "11101110",2520 => "11001111",2521 => "11000110",2522 => "10000010",2523 => "00000011",2524 => "10011001",2525 => "00111111",2526 => "11011111",2527 => "11001111",2528 => "01010111",2529 => "00010001",2530 => "10010001",2531 => "01001101",2532 => "11001000",2533 => "01000001",2534 => "10001011",2535 => "11001110",2536 => "00110000",2537 => "10101110",2538 => "00010010",2539 => "00001101",2540 => "11000100",2541 => "01001111",2542 => "01101000",2543 => "10111100",2544 => "10110110",2545 => "00110001",2546 => "00111011",2547 => "11100010",2548 => "10110010",2549 => "01000000",2550 => "01010010",2551 => "00100101",2552 => "10001111",2553 => "10101110",2554 => "00110111",2555 => "10011011",2556 => "10001110",2557 => "10111101",2558 => "01011010",2559 => "01100100",2560 => "00100000",2561 => "11010100",2562 => "10110111",2563 => "01011101",2564 => "00010011",2565 => "10001111",2566 => "11001110",2567 => "00000110",2568 => "11010001",2569 => "11110000",2570 => "10110001",2571 => "11010111",2572 => "10110101",2573 => "11101101",2574 => "01110010",2575 => "00000000",2576 => "11100100",2577 => "11100001",2578 => "00110101",2579 => "11001100",2580 => "10001010",2581 => "11100111",2582 => "10011101",2583 => "01010011",2584 => "10011100",2585 => "10011010",2586 => "10111010",2587 => "11111001",2588 => "11111000",2589 => "11111110",2590 => "10101111",2591 => "11010001",2592 => "10100110",2593 => "01111000",2594 => "10110111",2595 => "01001100",2596 => "10111101",2597 => "10011101",2598 => "10101101",2599 => "00001111",2600 => "10111101",2601 => "00100010",2602 => "11010100",2603 => "00000011",2604 => "11010000",2605 => "11100111",2606 => "11110011",2607 => "01111001",2608 => "11010101",2609 => "11001110",2610 => "10010010",2611 => "00010001",2612 => "00110111",2613 => "10110010",2614 => "00000000",2615 => "00111010",2616 => "10010110",2617 => "00001011",2618 => "11110000",2619 => "10111001",2620 => "00110100",2621 => "10101111",2622 => "00001111",2623 => "11010011",2624 => "01111000",2625 => "00011101",2626 => "01011101",2627 => "11000001",2628 => "10110101",2629 => "10101011",2630 => "01010000",2631 => "10010011",2632 => "01111001",2633 => "00100100",2634 => "11110111",2635 => "01000111",2636 => "10101110",2637 => "00001011",2638 => "10100000",2639 => "00101110",2640 => "01001100",2641 => "00101111",2642 => "10010001",2643 => "10010110",2644 => "11111111",2645 => "10001100",2646 => "00100000",2647 => "00000101",2648 => "10111001",2649 => "10110110",2650 => "00011101",2651 => "00011001",2652 => "00000010",2653 => "11000011",2654 => "11111101",2655 => "10100011",2656 => "11100011",2657 => "00011110",2658 => "10010101",2659 => "10010110",2660 => "11111100",2661 => "10000110",2662 => "10000010",2663 => "11111110",2664 => "00011111",2665 => "00110111",2666 => "11100101",2667 => "10000111",2668 => "10100010",2669 => "00110111",2670 => "00101010",2671 => "01000100",2672 => "11101010",2673 => "01111111",2674 => "01011000",2675 => "10110011",2676 => "10001001",2677 => "11111011",2678 => "10010101",2679 => "01011110",2680 => "00011100",2681 => "10010001",2682 => "00111101",2683 => "00100110",2684 => "01101101",2685 => "00101010",2686 => "10000000",2687 => "01010111",2688 => "01111100",2689 => "10011110",2690 => "11001100",2691 => "11011101",2692 => "01011000",2693 => "01001110",2694 => "01110010",2695 => "00001101",2696 => "00100100",2697 => "00101100",2698 => "00100001",2699 => "00110101",2700 => "10011010",2701 => "11101111",2702 => "00100110",2703 => "00111101",2704 => "10101010",2705 => "11011000",2706 => "11111100",2707 => "01100001",2708 => "00110011",2709 => "10001110",2710 => "10111101",2711 => "10101100",2712 => "11011010",2713 => "00111110",2714 => "01010010",2715 => "11010100",2716 => "10000101",2717 => "01110111",2718 => "10001001",2719 => "10010100",2720 => "01011010",2721 => "00010001",2722 => "00011111",2723 => "00100111",2724 => "01011100",2725 => "01110101",2726 => "10110001",2727 => "10010100",2728 => "00111011",2729 => "11001101",2730 => "10000010",2731 => "01101000",2732 => "01001100",2733 => "00101101",2734 => "00110111",2735 => "00010100",2736 => "00001111",2737 => "11011010",2738 => "00100111",2739 => "10001101",2740 => "11101001",2741 => "00111001",2742 => "00011110",2743 => "11111111",2744 => "10101101",2745 => "00110011",2746 => "10100111",2747 => "11101001",2748 => "10101011",2749 => "11110000",2750 => "00000010",2751 => "11101011",2752 => "10100000",2753 => "01001110",2754 => "01011110",2755 => "01001000",2756 => "00111111",2757 => "10001010",2758 => "00010011",2759 => "11001001",2760 => "10101100",2761 => "01101101",2762 => "11110101",2763 => "00110001",2764 => "01100011",2765 => "00111110",2766 => "00111101",2767 => "01111111",2768 => "11110010",2769 => "00100001",2770 => "11111001",2771 => "00010001",2772 => "10111011",2773 => "10001100",2774 => "01111001",2775 => "00001100",2776 => "01011011",2777 => "10011101",2778 => "10110000",2779 => "01001011",2780 => "01100000",2781 => "01110001",2782 => "11010110",2783 => "10001100",2784 => "10111001",2785 => "01001100",2786 => "01011100",2787 => "00011111",2788 => "10110111",2789 => "10100110",2790 => "10100000",2791 => "01101111",2792 => "10010011",2793 => "10010111",2794 => "11100111",2795 => "10000011",2796 => "00110011",2797 => "11100110",2798 => "11101010",2799 => "01010101",2800 => "11100000",2801 => "01100011",2802 => "10110010",2803 => "11101110",2804 => "11000101",2805 => "00100000",2806 => "11011111",2807 => "01110011",2808 => "10011000",2809 => "11011111",2810 => "11100111",2811 => "01111001",2812 => "00110011",2813 => "10101011",2814 => "10100011",2815 => "11010111",2816 => "00010101",2817 => "01000011",2818 => "10001010",2819 => "10101110",2820 => "10100101",2821 => "00010101",2822 => "11111010",2823 => "10001111",2824 => "00100101",2825 => "10010110",2826 => "10000000",2827 => "00000101",2828 => "01010001",2829 => "00010111",2830 => "01101001",2831 => "00101101",2832 => "11100101",2833 => "11110010",2834 => "01000001",2835 => "01100000",2836 => "01011001",2837 => "10001000",2838 => "01110011",2839 => "11011010",2840 => "01001110",2841 => "01110101",2842 => "10011110",2843 => "01000100",2844 => "00011011",2845 => "11100111",2846 => "01001011",2847 => "10100101",2848 => "11001101",2849 => "01110111",2850 => "10010001",2851 => "10100101",2852 => "11110100",2853 => "11111100",2854 => "01001101",2855 => "11111000",2856 => "10010011",2857 => "11011000",2858 => "00010100",2859 => "01000111",2860 => "00001000",2861 => "10001101",2862 => "10111110",2863 => "10110010",2864 => "11100101",2865 => "11000111",2866 => "11111000",2867 => "00100100",2868 => "01100101",2869 => "01000001",2870 => "10111000",2871 => "01011011",2872 => "00001110",2873 => "01000000",2874 => "01000000",2875 => "10111101",2876 => "11001001",2877 => "11010101",2878 => "10001001",2879 => "11101010",2880 => "10010101",2881 => "00000100",2882 => "01101000",2883 => "10001011",2884 => "11101000",2885 => "10111111",2886 => "10111000",2887 => "11101001",2888 => "01001101",2889 => "00000100",2890 => "11101010",2891 => "01000000",2892 => "00011000",2893 => "11000110",2894 => "00011100",2895 => "11100110",2896 => "10000100",2897 => "01001001",2898 => "01111111",2899 => "00010011",2900 => "01000110",2901 => "01111111",2902 => "01010111",2903 => "11010110",2904 => "10010101",2905 => "10000010",2906 => "00110111",2907 => "01010100",2908 => "00010001",2909 => "11110001",2910 => "10000110",2911 => "00100000",2912 => "10010110",2913 => "11101001",2914 => "00100010",2915 => "10110101",2916 => "00001111",2917 => "01000000",2918 => "01110111",2919 => "10101001",2920 => "01101001",2921 => "11101000",2922 => "01100100",2923 => "10100000",2924 => "11000111",2925 => "10110111",2926 => "10011011",2927 => "11101111",2928 => "00001111",2929 => "01001000",2930 => "01111110",2931 => "00111111",2932 => "01011100",2933 => "01011011",2934 => "00101111",2935 => "10011100",2936 => "00010011",2937 => "00111000",2938 => "00000001",2939 => "10100110",2940 => "00111010",2941 => "00000011",2942 => "11000111",2943 => "01111000",2944 => "00000011",2945 => "10110001",2946 => "00101010",2947 => "00001000",2948 => "01001001",2949 => "01101000",2950 => "01100100",2951 => "10101000",2952 => "11111111",2953 => "00001100",2954 => "10100010",2955 => "00101100",2956 => "11100111",2957 => "00001011",2958 => "11110010",2959 => "11011011",2960 => "01100111",2961 => "01110010",2962 => "00010111",2963 => "00100111",2964 => "00001101",2965 => "10100111",2966 => "11001111",2967 => "11001101",2968 => "11011001",2969 => "11100101",2970 => "01001110",2971 => "10110101",2972 => "10011011",2973 => "11010110",2974 => "10101110",2975 => "00011011",2976 => "00101001",2977 => "11010101",2978 => "00100110",2979 => "01001000",2980 => "11101000",2981 => "00011010",2982 => "10011111",2983 => "10000001",2984 => "11110010",2985 => "11111110",2986 => "01111001",2987 => "00111011",2988 => "11001001",2989 => "10011010",2990 => "01011011",2991 => "11111011",2992 => "00000001",2993 => "00110111",2994 => "00101010",2995 => "00000011",2996 => "11100100",2997 => "00001100",2998 => "10000001",2999 => "11101000",3000 => "00001100",3001 => "11111010",3002 => "00000101",3003 => "01010101",3004 => "00101110",3005 => "01001110",3006 => "10010100",3007 => "01011111",3008 => "11100000",3009 => "01110000",3010 => "01100100",3011 => "01110000",3012 => "10110011",3013 => "11111001",3014 => "01000000",3015 => "00101010",3016 => "01101000",3017 => "11011001",3018 => "10101011",3019 => "01111000",3020 => "10101000",3021 => "01010000",3022 => "01011101",3023 => "01010100",3024 => "11010101",3025 => "11110010",3026 => "11111011",3027 => "10011000",3028 => "10001000",3029 => "10001111",3030 => "11110101",3031 => "01000100",3032 => "10111010",3033 => "01011101",3034 => "00011101",3035 => "10100100",3036 => "11000000",3037 => "00001000",3038 => "00101110",3039 => "00010000",3040 => "00101101",3041 => "10110111",3042 => "11111100",3043 => "00110000",3044 => "10100011",3045 => "11111101",3046 => "01101010",3047 => "10011111",3048 => "01011100",3049 => "11001011",3050 => "00110111",3051 => "11110110",3052 => "11100101",3053 => "10101111",3054 => "00101010",3055 => "11111101",3056 => "01111000",3057 => "11111110",3058 => "00110100",3059 => "01111000",3060 => "00110001",3061 => "00001110",3062 => "11001011",3063 => "00011011",3064 => "00001001",3065 => "11100101",3066 => "10001101",3067 => "10101001",3068 => "01101001",3069 => "11111101",3070 => "01010111",3071 => "01011001",3072 => "01000001",3073 => "00110111",3074 => "10100000",3075 => "00001100",3076 => "01100100",3077 => "11010101",3078 => "10000100",3079 => "01000000",3080 => "11010110",3081 => "10000000",3082 => "00111110",3083 => "10100010",3084 => "10010110",3085 => "01101101",3086 => "10010111",3087 => "10110001",3088 => "10000111",3089 => "10100101",3090 => "11110001",3091 => "00111001",3092 => "11111011",3093 => "11011100",3094 => "10001110",3095 => "00011111",3096 => "01111100",3097 => "00001011",3098 => "01001011",3099 => "01101000",3100 => "11010110",3101 => "01100100",3102 => "11110000",3103 => "11101000",3104 => "11110010",3105 => "11111100",3106 => "01000000",3107 => "10001000",3108 => "10011101",3109 => "01101000",3110 => "11101101",3111 => "10011011",3112 => "01101100",3113 => "11010010",3114 => "10100100",3115 => "01011110",3116 => "00111110",3117 => "01011100",3118 => "00111010",3119 => "01010000",3120 => "00100000",3121 => "11100110",3122 => "10010001",3123 => "00000111",3124 => "11010100",3125 => "00100011",3126 => "11101111",3127 => "01001001",3128 => "00001010",3129 => "11101111",3130 => "11000100",3131 => "10101000",3132 => "01110001",3133 => "00010111",3134 => "11000010",3135 => "01000000",3136 => "11000000",3137 => "10011010",3138 => "11110010",3139 => "11111000",3140 => "11000100",3141 => "00011110",3142 => "11010100",3143 => "00101001",3144 => "00011000",3145 => "11110011",3146 => "10101101",3147 => "11001010",3148 => "00011100",3149 => "10111010",3150 => "00010110",3151 => "01101111",3152 => "00100100",3153 => "11101100",3154 => "11000101",3155 => "00001001",3156 => "11100000",3157 => "11111001",3158 => "01010101",3159 => "10011111",3160 => "01001110",3161 => "11111010",3162 => "10011001",3163 => "10101010",3164 => "11110000",3165 => "10100101",3166 => "10111011",3167 => "01000101",3168 => "00101101",3169 => "11000100",3170 => "11010000",3171 => "11101111",3172 => "01100101",3173 => "01001001",3174 => "10111011",3175 => "11111110",3176 => "00000000",3177 => "01110000",3178 => "11110011",3179 => "00000101",3180 => "01001110",3181 => "11011100",3182 => "00100001",3183 => "10010110",3184 => "10101101",3185 => "11101100",3186 => "10010101",3187 => "00001010",3188 => "00101010",3189 => "00101000",3190 => "11011101",3191 => "01001000",3192 => "00001101",3193 => "11100110",3194 => "10100001",3195 => "01110001",3196 => "11101101",3197 => "10010010",3198 => "10110100",3199 => "11001000",3200 => "00101001",3201 => "10111010",3202 => "10010011",3203 => "00100001",3204 => "10101110",3205 => "11000000",3206 => "00001110",3207 => "10101100",3208 => "01001010",3209 => "00111100",3210 => "00100101",3211 => "01011000",3212 => "00010001",3213 => "00011101",3214 => "10000111",3215 => "00100000",3216 => "01010111",3217 => "11110001",3218 => "00001001",3219 => "10101101",3220 => "01111011",3221 => "00001011",3222 => "10101010",3223 => "11100100",3224 => "10010101",3225 => "00100100",3226 => "01110101",3227 => "00010011",3228 => "11110010",3229 => "11100100",3230 => "01000100",3231 => "10010000",3232 => "10000100",3233 => "10010011",3234 => "11100001",3235 => "01011011",3236 => "11110001",3237 => "10110111",3238 => "11001100",3239 => "00100111",3240 => "11001001",3241 => "01010101",3242 => "11001110",3243 => "10000000",3244 => "10011000",3245 => "00110000",3246 => "10111010",3247 => "01100100",3248 => "01111001",3249 => "11000110",3250 => "11100111",3251 => "01101101",3252 => "11100100",3253 => "10101001",3254 => "00001011",3255 => "00101001",3256 => "01000001",3257 => "10010110",3258 => "01000100",3259 => "01011100",3260 => "10101010",3261 => "11001010",3262 => "10000101",3263 => "10011001",3264 => "11000011",3265 => "01111011",3266 => "01001010",3267 => "11100001",3268 => "01001001",3269 => "10101100",3270 => "00010100",3271 => "00111100",3272 => "01100011",3273 => "10000001",3274 => "11111011",3275 => "01110011",3276 => "10001001",3277 => "10011011",3278 => "00001010",3279 => "01001011",3280 => "01010100",3281 => "11111111",3282 => "00101011",3283 => "10011101",3284 => "00001001",3285 => "10111110",3286 => "11000100",3287 => "01011001",3288 => "11011101",3289 => "00111101",3290 => "00110010",3291 => "01010100",3292 => "11110011",3293 => "01001101",3294 => "11010000",3295 => "10111100",3296 => "00001101",3297 => "11001011",3298 => "00100111",3299 => "11100111",3300 => "10100010",3301 => "01100011",3302 => "00100111",3303 => "11100100",3304 => "11001011",3305 => "10001010",3306 => "10001010",3307 => "11000110",3308 => "01110011",3309 => "10001000",3310 => "10010101",3311 => "00011101",3312 => "10011101",3313 => "01001000",3314 => "00100010",3315 => "01001001",3316 => "10010101",3317 => "00011011",3318 => "10001111",3319 => "01010101",3320 => "11111000",3321 => "00101101",3322 => "00100101",3323 => "01010101",3324 => "11100011",3325 => "10101110",3326 => "01011100",3327 => "11011001",3328 => "01100111",3329 => "11010000",3330 => "01000010",3331 => "00010001",3332 => "01101001",3333 => "11000100",3334 => "01000000",3335 => "10101010",3336 => "10001000",3337 => "00000101",3338 => "00111111",3339 => "01111100",3340 => "01010101",3341 => "11000000",3342 => "10110110",3343 => "01110111",3344 => "10101110",3345 => "00111001",3346 => "01000001",3347 => "10000000",3348 => "00000000",3349 => "01000100",3350 => "11011110",3351 => "11101000",3352 => "10000010",3353 => "00011000",3354 => "00110100",3355 => "11111010",3356 => "11100010",3357 => "10010000",3358 => "10010000",3359 => "10010010",3360 => "11011101",3361 => "00000100",3362 => "10100111",3363 => "01101001",3364 => "01110111",3365 => "00100100",3366 => "11010111",3367 => "00111000",3368 => "10000000",3369 => "01010011",3370 => "11110110",3371 => "01011011",3372 => "11100000",3373 => "10111110",3374 => "11101110",3375 => "00001110",3376 => "01010010",3377 => "10100111",3378 => "11100110",3379 => "10000111",3380 => "00101001",3381 => "00110110",3382 => "00100101",3383 => "11001010",3384 => "01001111",3385 => "01001000",3386 => "11111101",3387 => "00000001",3388 => "01111111",3389 => "01001001",3390 => "11100000",3391 => "01001010",3392 => "00010001",3393 => "10101000",3394 => "00010000",3395 => "11010100",3396 => "01101111",3397 => "10110101",3398 => "00001001",3399 => "11000010",3400 => "01011110",3401 => "01011110",3402 => "11110101",3403 => "10011111",3404 => "11100010",3405 => "01100111",3406 => "01001010",3407 => "01100011",3408 => "11010101",3409 => "01100011",3410 => "11001000",3411 => "11100010",3412 => "11110001",3413 => "10101011",3414 => "10000110",3415 => "01111011",3416 => "00111001",3417 => "11110000",3418 => "01110001",3419 => "10000010",3420 => "01110001",3421 => "10111001",3422 => "10010011",3423 => "00001101",3424 => "11111111",3425 => "01000001",3426 => "00100110",3427 => "11001101",3428 => "01001010",3429 => "10010101",3430 => "10101000",3431 => "10000000",3432 => "10110000",3433 => "00111110",3434 => "01100011",3435 => "01011000",3436 => "10010000",3437 => "11010011",3438 => "10011111",3439 => "01011001",3440 => "01100001",3441 => "11110000",3442 => "00011100",3443 => "11111101",3444 => "10100110",3445 => "11010010",3446 => "10111001",3447 => "00101001",3448 => "11001011",3449 => "11100110",3450 => "01100011",3451 => "01101101",3452 => "10010101",3453 => "10101000",3454 => "00100010",3455 => "01011110",3456 => "01111001",3457 => "01011010",3458 => "11011011",3459 => "10000110",3460 => "10101010",3461 => "01110010",3462 => "00111100",3463 => "10000011",3464 => "10100101",3465 => "11010110",3466 => "10010110",3467 => "00110010",3468 => "11011010",3469 => "01000110",3470 => "00001110",3471 => "00011010",3472 => "00010000",3473 => "00110101",3474 => "11111001",3475 => "11011110",3476 => "11111110",3477 => "00010111",3478 => "10110111",3479 => "10111001",3480 => "11101111",3481 => "10001000",3482 => "00111000",3483 => "00100100",3484 => "10010111",3485 => "11111100",3486 => "01100010",3487 => "10111111",3488 => "01100000",3489 => "01011111",3490 => "11111001",3491 => "00001101",3492 => "01010110",3493 => "00011110",3494 => "01111011",3495 => "11111000",3496 => "01000011",3497 => "01011001",3498 => "10101011",3499 => "11100111",3500 => "01111110",3501 => "01101101",3502 => "11011101",3503 => "11011111",3504 => "10101000",3505 => "00100111",3506 => "10100010",3507 => "10101000",3508 => "01000101",3509 => "11000010",3510 => "00010110",3511 => "10100000",3512 => "01110101",3513 => "10000001",3514 => "01011000",3515 => "10011000",3516 => "11110000",3517 => "00010001",3518 => "00010100",3519 => "10110111",3520 => "01000110",3521 => "10011101",3522 => "10100110",3523 => "11100110",3524 => "11010100",3525 => "11010110",3526 => "00101010",3527 => "11011011",3528 => "10000011",3529 => "11011011",3530 => "11100110",3531 => "11110001",3532 => "11010010",3533 => "11100011",3534 => "10110010",3535 => "10111001",3536 => "10001000",3537 => "00010011",3538 => "10110010",3539 => "00101101",3540 => "10001010",3541 => "01101010",3542 => "11001111",3543 => "11100111",3544 => "10100001",3545 => "00011001",3546 => "01011100",3547 => "10100001",3548 => "10110001",3549 => "11011011",3550 => "10110011",3551 => "00010001",3552 => "00011000",3553 => "01111011",3554 => "01111000",3555 => "00010110",3556 => "00010010",3557 => "10010010",3558 => "10110110",3559 => "10101101",3560 => "10011111",3561 => "00001011",3562 => "01010111",3563 => "10111100",3564 => "00101001",3565 => "10110101",3566 => "10100000",3567 => "00001010",3568 => "10000011",3569 => "10001011",3570 => "10111100",3571 => "00001100",3572 => "10011001",3573 => "01100001",3574 => "10010011",3575 => "11011011",3576 => "01111011",3577 => "11100011",3578 => "01111100",3579 => "10100001",3580 => "11010100",3581 => "01100110",3582 => "01101111",3583 => "01101111",3584 => "00100100",3585 => "11000010",3586 => "10111001",3587 => "10101100",3588 => "00100101",3589 => "10001110",3590 => "11001101",3591 => "00011010",3592 => "01001001",3593 => "01110011",3594 => "00100100",3595 => "10010100",3596 => "11011110",3597 => "01001000",3598 => "10111110",3599 => "10001111",3600 => "00011000",3601 => "11000100",3602 => "11100100",3603 => "11110011",3604 => "11010010",3605 => "11001010",3606 => "00110000",3607 => "00011110",3608 => "10011111",3609 => "01011000",3610 => "00100000",3611 => "11101010",3612 => "01110110",3613 => "11110001",3614 => "00000111",3615 => "11000111",3616 => "01000011",3617 => "01100101",3618 => "10111010",3619 => "00010100",3620 => "11010001",3621 => "01011110",3622 => "10000001",3623 => "00010001",3624 => "11000000",3625 => "10011000",3626 => "00000011",3627 => "11100100",3628 => "10101001",3629 => "00010011",3630 => "00000111",3631 => "00101111",3632 => "11101100",3633 => "10101100",3634 => "00010101",3635 => "10110100",3636 => "11100011",3637 => "00000001",3638 => "00011100",3639 => "00101001",3640 => "10010011",3641 => "11101100",3642 => "11000000",3643 => "11011001",3644 => "10110000",3645 => "10010010",3646 => "00111000",3647 => "00010101",3648 => "10110100",3649 => "11110001",3650 => "01111001",3651 => "00001101",3652 => "00010000",3653 => "00110100",3654 => "10101011",3655 => "11110001",3656 => "01111001",3657 => "00000111",3658 => "11001101",3659 => "00000100",3660 => "11110000",3661 => "01000100",3662 => "10110110",3663 => "10000100",3664 => "11001101",3665 => "10000100",3666 => "10110101",3667 => "00001100",3668 => "00000010",3669 => "10111001",3670 => "11000010",3671 => "10110100",3672 => "01000101",3673 => "11001011",3674 => "00000110",3675 => "01111010",3676 => "10101111",3677 => "00111110",3678 => "10111110",3679 => "10110011",3680 => "11000011",3681 => "11011111",3682 => "01100000",3683 => "11111010",3684 => "11111110",3685 => "01001100",3686 => "11001111",3687 => "10001111",3688 => "11101000",3689 => "11110100",3690 => "00100010",3691 => "11001000",3692 => "10011111",3693 => "00111100",3694 => "10000001",3695 => "00110010",3696 => "11011010",3697 => "00101000",3698 => "01100000",3699 => "00011001",3700 => "01011011",3701 => "10110000",3702 => "00100001",3703 => "11101010",3704 => "01000010",3705 => "01100010",3706 => "01111111",3707 => "10101100",3708 => "00011011",3709 => "10000100",3710 => "00001011",3711 => "00010001",3712 => "10000010",3713 => "00111101",3714 => "10001010",3715 => "10010111",3716 => "10010111",3717 => "01101000",3718 => "00100000",3719 => "01101000",3720 => "01010100",3721 => "01000110",3722 => "00010000",3723 => "00000010",3724 => "10000111",3725 => "01111111",3726 => "10000010",3727 => "01100111",3728 => "11100010",3729 => "01110110",3730 => "11000110",3731 => "00001001",3732 => "00010111",3733 => "10101111",3734 => "11100010",3735 => "01001100",3736 => "10011110",3737 => "10110100",3738 => "11101001",3739 => "10001001",3740 => "10100100",3741 => "00111101",3742 => "00011001",3743 => "00001111",3744 => "00101010",3745 => "10000011",3746 => "11100000",3747 => "10011100",3748 => "00000000",3749 => "10110011",3750 => "00101110",3751 => "10110100",3752 => "01111000",3753 => "10110011",3754 => "00101111",3755 => "10111101",3756 => "01100000",3757 => "11111000",3758 => "01111101",3759 => "01001011",3760 => "11000011",3761 => "10000111",3762 => "00011110",3763 => "10011001",3764 => "10111000",3765 => "11110010",3766 => "01100001",3767 => "00101001",3768 => "10101011",3769 => "00110001",3770 => "01001000",3771 => "00011010",3772 => "00100101",3773 => "01011111",3774 => "01100011",3775 => "00000101",3776 => "00011010",3777 => "01010011",3778 => "11110000",3779 => "00111111",3780 => "10101101",3781 => "00000001",3782 => "10110000",3783 => "10100011",3784 => "01010011",3785 => "00011011",3786 => "01100111",3787 => "01111101",3788 => "10110000",3789 => "10010111",3790 => "10111000",3791 => "01000111",3792 => "01010001",3793 => "00000001",3794 => "00110001",3795 => "01100100",3796 => "00000110",3797 => "10111011",3798 => "00010010",3799 => "00111110",3800 => "10010010",3801 => "10001001",3802 => "11101110",3803 => "01001000",3804 => "11100110",3805 => "01000010",3806 => "00101111",3807 => "11110010",3808 => "11011110",3809 => "10011001",3810 => "11000010",3811 => "11000100",3812 => "00010110",3813 => "00110011",3814 => "01110110",3815 => "11000000",3816 => "11101001",3817 => "10000010",3818 => "11101011",3819 => "01101011",3820 => "00001010",3821 => "10101110",3822 => "01011000",3823 => "01000110",3824 => "01010010",3825 => "11110100",3826 => "01011100",3827 => "10000001",3828 => "10010110",3829 => "11001101",3830 => "11000000",3831 => "11110100",3832 => "11101110",3833 => "00001110",3834 => "11100001",3835 => "00010001",3836 => "01100011",3837 => "10111100",3838 => "00110001",3839 => "00001110",3840 => "01100001",3841 => "01101011",3842 => "01010011",3843 => "01100100",3844 => "00011000",3845 => "10000101",3846 => "00110110",3847 => "01001110",3848 => "01010101",3849 => "11010111",3850 => "00010001",3851 => "00110110",3852 => "00011001",3853 => "10100001",3854 => "01100000",3855 => "10000110",3856 => "01100000",3857 => "11011000",3858 => "11001011",3859 => "10010101",3860 => "10010001",3861 => "10110011",3862 => "00001110",3863 => "01011100",3864 => "11101000",3865 => "00000100",3866 => "01000100",3867 => "10010100",3868 => "00001100",3869 => "11010100",3870 => "00100010",3871 => "00011001",3872 => "10111000",3873 => "11011001",3874 => "10111000",3875 => "01001011",3876 => "11000110",3877 => "10100100",3878 => "10111101",3879 => "10100000",3880 => "01010010",3881 => "11101010",3882 => "10111101",3883 => "11000011",3884 => "00101010",3885 => "01110000",3886 => "01001011",3887 => "10000100",3888 => "10101010",3889 => "00010100",3890 => "10101100",3891 => "11011111",3892 => "00101000",3893 => "01101100",3894 => "01100000",3895 => "11011100",3896 => "11101100",3897 => "00010100",3898 => "10011101",3899 => "01101100",3900 => "01101111",3901 => "10010111",3902 => "00101111",3903 => "10011110",3904 => "10101101",3905 => "11100111",3906 => "10110100",3907 => "01001110",3908 => "11111101",3909 => "10110010",3910 => "11100100",3911 => "11010000",3912 => "11100100",3913 => "00011001",3914 => "01111101",3915 => "00101001",3916 => "10001110",3917 => "01000101",3918 => "10110010",3919 => "10111010",3920 => "00000100",3921 => "00111100",3922 => "00101110",3923 => "01100111",3924 => "10010101",3925 => "00111010",3926 => "10010101",3927 => "10011000",3928 => "10010101",3929 => "00101101",3930 => "01100110",3931 => "00110110",3932 => "11111110",3933 => "00000010",3934 => "10100000",3935 => "00011011",3936 => "00101100",3937 => "01011010",3938 => "01001001",3939 => "00000111",3940 => "01001110",3941 => "11010000",3942 => "11101001",3943 => "11011110",3944 => "11001101",3945 => "01101011",3946 => "10110110",3947 => "00000111",3948 => "10000111",3949 => "11111001",3950 => "00101110",3951 => "00110011",3952 => "10011000",3953 => "10100100",3954 => "11101010",3955 => "10110011",3956 => "01111101",3957 => "11011100",3958 => "01001011",3959 => "10111011",3960 => "10100110",3961 => "01010001",3962 => "00000010",3963 => "11110010",3964 => "01001111",3965 => "00011111",3966 => "00101111",3967 => "00100011",3968 => "00001000",3969 => "01101001",3970 => "01011110",3971 => "00100010",3972 => "10110111",3973 => "00011010",3974 => "00111100",3975 => "11111000",3976 => "01010011",3977 => "11101110",3978 => "01101001",3979 => "01110001",3980 => "11001001",3981 => "10110011",3982 => "11000011",3983 => "11011101",3984 => "11001010",3985 => "01001010",3986 => "10110101",3987 => "11100001",3988 => "00000001",3989 => "00110110",3990 => "00010010",3991 => "11100001",3992 => "11111100",3993 => "01100101",3994 => "01001010",3995 => "10111100",3996 => "00010011",3997 => "00101111",3998 => "10100110",3999 => "10011011",4000 => "00101111",4001 => "01111100",4002 => "00010000",4003 => "00011101",4004 => "10100001",4005 => "00100111",4006 => "11000010",4007 => "11101000",4008 => "01100001",4009 => "00111111",4010 => "01110100",4011 => "00010111",4012 => "11110110",4013 => "01101110",4014 => "10000010",4015 => "00001110",4016 => "11001101",4017 => "00011001",4018 => "11111110",4019 => "01010101",4020 => "00000011",4021 => "10011011",4022 => "00100010",4023 => "11101010",4024 => "11000100",4025 => "00100101",4026 => "11101100",4027 => "01001110",4028 => "10101000",4029 => "01101011",4030 => "11000110",4031 => "01010010",4032 => "01100011",4033 => "00001010",4034 => "10001001",4035 => "10010000",4036 => "00100111",4037 => "00011000",4038 => "01010101",4039 => "11101000",4040 => "01110101",4041 => "01110010",4042 => "00110100",4043 => "11010001",4044 => "00001001",4045 => "11000000",4046 => "01101110",4047 => "00010000",4048 => "10011011",4049 => "00010000",4050 => "10100101",4051 => "01101111",4052 => "11011001",4053 => "11011110",4054 => "10110111",4055 => "01110001",4056 => "10110101",4057 => "00110001",4058 => "00011011",4059 => "11000000",4060 => "00101001",4061 => "10111010",4062 => "11110011",4063 => "11010010",4064 => "01000111",4065 => "10000010",4066 => "11110010",4067 => "11000111",4068 => "10111110",4069 => "01001110",4070 => "11001100",4071 => "01000100",4072 => "11001111",4073 => "01110010",4074 => "01001111",4075 => "00000101",4076 => "01100000",4077 => "10010110",4078 => "01010110",4079 => "00110111",4080 => "10110001",4081 => "10110110",4082 => "01100100",4083 => "11100011",4084 => "10011010",4085 => "11011101",4086 => "11101110",4087 => "10110010",4088 => "01000011",4089 => "00101000",4090 => "11010011",4091 => "00111100",4092 => "10101011",4093 => "01101110",4094 => "10100011",4095 => "00100011",4096 => "01111101",4097 => "10001000",4098 => "10111100",4099 => "11110001",4100 => "11111011",4101 => "11100000",4102 => "00111000",4103 => "01100111",4104 => "10011100",4105 => "11110110",4106 => "00101111",4107 => "01000011",4108 => "10100101",4109 => "01000011",4110 => "11000110",4111 => "10111111",4112 => "10010111",4113 => "11101110",4114 => "10110101",4115 => "11101100",4116 => "00100101",4117 => "10000010",4118 => "11101100",4119 => "01100011",4120 => "00111000",4121 => "01110010",4122 => "10000011",4123 => "10011100",4124 => "11111010",4125 => "10001011",4126 => "10111100",4127 => "01011101",4128 => "00010110",4129 => "01100100",4130 => "01011101",4131 => "10100001",4132 => "10011011",4133 => "10000010",4134 => "00010101",4135 => "10000000",4136 => "00001000",4137 => "11101000",4138 => "10111100",4139 => "00110000",4140 => "00001010",4141 => "01000111",4142 => "01111010",4143 => "10000011",4144 => "00010001",4145 => "00111001",4146 => "10011111",4147 => "11101011",4148 => "00011110",4149 => "11010010",4150 => "10101100",4151 => "00100100",4152 => "10000010",4153 => "11111101",4154 => "10101001",4155 => "10011100",4156 => "11101011",4157 => "01011100",4158 => "01010001",4159 => "00100111",4160 => "11001110",4161 => "10110010",4162 => "00011010",4163 => "00011100",4164 => "00100111",4165 => "00111010",4166 => "11011111",4167 => "00110101",4168 => "01010011",4169 => "11101101",4170 => "00011010",4171 => "11101100",4172 => "00000000",4173 => "11001001",4174 => "10000011",4175 => "01111011",4176 => "11001001",4177 => "11110100",4178 => "10011110",4179 => "01011100",4180 => "10010001",4181 => "10101100",4182 => "01001111",4183 => "01110010",4184 => "01100101",4185 => "00100111",4186 => "01001111",4187 => "11011111",4188 => "00110110",4189 => "11111011",4190 => "01111011",4191 => "10011010",4192 => "10001000",4193 => "00010010",4194 => "10000101",4195 => "01001000",4196 => "10000011",4197 => "11011100",4198 => "11011011",4199 => "10001011",4200 => "00001100",4201 => "00111111",4202 => "00101101",4203 => "00010010",4204 => "11100111",4205 => "11010101",4206 => "10101101",4207 => "11101000",4208 => "01100101",4209 => "10011010",4210 => "11010101",4211 => "10111011",4212 => "10011101",4213 => "01000001",4214 => "10011110",4215 => "00001001",4216 => "10010011",4217 => "01110010",4218 => "01101010",4219 => "11101011",4220 => "10101101",4221 => "01001101",4222 => "00110101",4223 => "11101111",4224 => "00001100",4225 => "10000111",4226 => "10011011",4227 => "10011010",4228 => "00101110",4229 => "00010011",4230 => "01001011",4231 => "11011110",4232 => "11010011",4233 => "01011101",4234 => "01011000",4235 => "01011001",4236 => "00000101",4237 => "11001100",4238 => "10010011",4239 => "01000110",4240 => "10110100",4241 => "00111011",4242 => "01001001",4243 => "10100100",4244 => "11001001",4245 => "11111000",4246 => "01010111",4247 => "11000100",4248 => "00101001",4249 => "00000110",4250 => "00001110",4251 => "00100001",4252 => "00011110",4253 => "10000100",4254 => "01000011",4255 => "01100101",4256 => "11000101",4257 => "01011110",4258 => "10101010",4259 => "01100001",4260 => "11101001",4261 => "01001111",4262 => "01110111",4263 => "00110000",4264 => "11111011",4265 => "01101001",4266 => "10010010",4267 => "10010100",4268 => "01001101",4269 => "10100101",4270 => "11001111",4271 => "11000110",4272 => "10100011",4273 => "11000001",4274 => "00010100",4275 => "01111010",4276 => "11101000",4277 => "11001100",4278 => "11001100",4279 => "01010100",4280 => "11000101",4281 => "11010010",4282 => "10010011",4283 => "11010010",4284 => "10010010",4285 => "01101110",4286 => "01000000",4287 => "10011101",4288 => "11101001",4289 => "10111010",4290 => "00000101",4291 => "10001010",4292 => "11001010",4293 => "01010010",4294 => "11000100",4295 => "10001111",4296 => "11111101",4297 => "00010000",4298 => "10011110",4299 => "11111000",4300 => "10000101",4301 => "11100100",4302 => "01010101",4303 => "00000010",4304 => "11100110",4305 => "11000101",4306 => "10101011",4307 => "01111011",4308 => "10111111",4309 => "01011100",4310 => "11001001",4311 => "10000010",4312 => "10010111",4313 => "10000011",4314 => "11111111",4315 => "10110111",4316 => "10100001",4317 => "11111111",4318 => "01101100",4319 => "11000001",4320 => "11100111",4321 => "01001010",4322 => "10000010",4323 => "00001001",4324 => "10100011",4325 => "01010001",4326 => "11011011",4327 => "10001111",4328 => "01011110",4329 => "00001110",4330 => "10001101",4331 => "10101011",4332 => "00010000",4333 => "11001111",4334 => "01010110",4335 => "00010000",4336 => "00100101",4337 => "01111100",4338 => "00101110",4339 => "00110101",4340 => "00011100",4341 => "10110111",4342 => "01011000",4343 => "00111001",4344 => "01010000",4345 => "11001100",4346 => "10111000",4347 => "10000111",4348 => "01110010",4349 => "01001111",4350 => "00110011",4351 => "11011001",4352 => "00110010",4353 => "01000110",4354 => "00100111",4355 => "11001100",4356 => "10001001",4357 => "00110011",4358 => "11111111",4359 => "01110010",4360 => "11111011",4361 => "00111000",4362 => "10010010",4363 => "00110000",4364 => "01011010",4365 => "10010100",4366 => "10000001",4367 => "11100000",4368 => "10000011",4369 => "10000111",4370 => "11100000",4371 => "00000111",4372 => "10001101",4373 => "11100101",4374 => "00101001",4375 => "11000000",4376 => "10100101",4377 => "11010001",4378 => "11000001",4379 => "11100011",4380 => "01011010",4381 => "00110101",4382 => "11001010",4383 => "10010101",4384 => "00000000",4385 => "10011100",4386 => "01011011",4387 => "11011111",4388 => "00001101",4389 => "10011111",4390 => "00011111",4391 => "10010011",4392 => "01110101",4393 => "11111001",4394 => "11011111",4395 => "01101011",4396 => "00111111",4397 => "11111111",4398 => "00001101",4399 => "10010011",4400 => "10001011",4401 => "00010111",4402 => "00001111",4403 => "11001111",4404 => "10001101",4405 => "11101110",4406 => "10100100",4407 => "00000111",4408 => "01101011",4409 => "01110100",4410 => "00110110",4411 => "00101011",4412 => "01011100",4413 => "00011100",4414 => "10101100",4415 => "01110111",4416 => "00101110",4417 => "10110101",4418 => "00110110",4419 => "11110100",4420 => "11011111",4421 => "11001101",4422 => "01101000",4423 => "10110100",4424 => "01000110",4425 => "11001000",4426 => "00110000",4427 => "01100111",4428 => "11011001",4429 => "10011000",4430 => "10010011",4431 => "01100100",4432 => "01100000",4433 => "00010111",4434 => "10001110",4435 => "11000111",4436 => "10000001",4437 => "10011010",4438 => "10100100",4439 => "11010100",4440 => "01010110",4441 => "00011111",4442 => "00110000",4443 => "00010011",4444 => "01110101",4445 => "01111101",4446 => "11000100",4447 => "11010011",4448 => "01110001",4449 => "10010000",4450 => "00111110",4451 => "00001000",4452 => "01011100",4453 => "01010011",4454 => "11000110",4455 => "11110100",4456 => "10100110",4457 => "01001100",4458 => "10011010",4459 => "00010011",4460 => "10011110",4461 => "01000110",4462 => "11001100",4463 => "01111111",4464 => "00011101",4465 => "01001111",4466 => "01001000",4467 => "00101101",4468 => "00100010",4469 => "10111011",4470 => "10001111",4471 => "10100001",4472 => "01010000",4473 => "00011000",4474 => "01010101",4475 => "00100001",4476 => "01111110",4477 => "11111110",4478 => "00101000",4479 => "01001111",4480 => "00011111",4481 => "10110100",4482 => "01100100",4483 => "00001100",4484 => "00101010",4485 => "11010010",4486 => "10101010",4487 => "10110100",4488 => "10111111",4489 => "10010010",4490 => "11010101",4491 => "10101001",4492 => "11010001",4493 => "10100100",4494 => "10000010",4495 => "10110010",4496 => "10110100",4497 => "10101001",4498 => "00101010",4499 => "00011010",4500 => "00101111",4501 => "10111101",4502 => "11100001",4503 => "10001011",4504 => "11011100",4505 => "00010010",4506 => "00011010",4507 => "11101111",4508 => "11001100",4509 => "00000110",4510 => "01110111",4511 => "01101101",4512 => "00111100",4513 => "00010110",4514 => "01110100",4515 => "10100101",4516 => "00000111",4517 => "10000010",4518 => "01001110",4519 => "10011111",4520 => "10100011",4521 => "11011010",4522 => "10100100",4523 => "10101100",4524 => "11110010",4525 => "10001110",4526 => "00011001",4527 => "10011010",4528 => "10100001",4529 => "00111001",4530 => "11000011",4531 => "01011100",4532 => "01100000",4533 => "11111110",4534 => "10010001",4535 => "11111010",4536 => "01011010",4537 => "01000001",4538 => "00000000",4539 => "11010011",4540 => "10011010",4541 => "00001011",4542 => "11010101",4543 => "11010001",4544 => "00011110",4545 => "00011101",4546 => "00100111",4547 => "01000110",4548 => "10011010",4549 => "10101100",4550 => "10010101",4551 => "01000110",4552 => "11000101",4553 => "00011011",4554 => "10100010",4555 => "00011011",4556 => "11111101",4557 => "00111100",4558 => "10010010",4559 => "10100100",4560 => "11111010",4561 => "01000011",4562 => "00001100",4563 => "10100000",4564 => "10110000",4565 => "11000111",4566 => "11111111",4567 => "10110011",4568 => "01000101",4569 => "00101100",4570 => "01001011",4571 => "11111111",4572 => "10000110",4573 => "01011000",4574 => "11111011",4575 => "01010111",4576 => "00101110",4577 => "00011100",4578 => "11101110",4579 => "11101000",4580 => "10110100",4581 => "10100111",4582 => "00011011",4583 => "00011100",4584 => "10000000",4585 => "10010001",4586 => "10111011",4587 => "11011000",4588 => "10001111",4589 => "01111001",4590 => "01001101",4591 => "00100001",4592 => "01111000",4593 => "00010001",4594 => "01000000",4595 => "10011010",4596 => "01110101",4597 => "11011010",4598 => "11111100",4599 => "00001011",4600 => "11001010",4601 => "00101010",4602 => "00110100",4603 => "11101110",4604 => "00111001",4605 => "11010000",4606 => "11011100",4607 => "00101100",4608 => "11010100",4609 => "01100110",4610 => "01101110",4611 => "11001101",4612 => "00101000",4613 => "01101101",4614 => "01100011",4615 => "10110100",4616 => "01100000",4617 => "11111000",4618 => "10001100",4619 => "11110001",4620 => "01000001",4621 => "10010000",4622 => "00001001",4623 => "11101101",4624 => "01000001",4625 => "10000000",4626 => "01101100",4627 => "11000011",4628 => "10110111",4629 => "01001010",4630 => "11001100",4631 => "00001101",4632 => "01011011",4633 => "10010100",4634 => "11010101",4635 => "11110100",4636 => "10001100",4637 => "01010110",4638 => "11111010",4639 => "00000011",4640 => "01011011",4641 => "11100010",4642 => "00111010",4643 => "10100010",4644 => "10011101",4645 => "01101000",4646 => "01110100",4647 => "10101001",4648 => "11001100",4649 => "11111111",4650 => "00100111",4651 => "00000111",4652 => "01000111",4653 => "11110110",4654 => "01011100",4655 => "00011001",4656 => "10110110",4657 => "10011100",4658 => "01001100",4659 => "11001101",4660 => "11100100",4661 => "00010010",4662 => "10111110",4663 => "10011001",4664 => "11111101",4665 => "11001000",4666 => "01000101",4667 => "01100101",4668 => "00010001",4669 => "01000110",4670 => "11111001",4671 => "01000101",4672 => "01111000",4673 => "11101100",4674 => "11100110",4675 => "11000001",4676 => "11001001",4677 => "00000000",4678 => "01100111",4679 => "10001000",4680 => "10001011",4681 => "01101101",4682 => "10110100",4683 => "10000110",4684 => "11101010",4685 => "11001001",4686 => "01001101",4687 => "01001101",4688 => "00111101",4689 => "10101100",4690 => "11101000",4691 => "00000010",4692 => "11110111",4693 => "00010001",4694 => "01110101",4695 => "10100000",4696 => "00010000",4697 => "00011111",4698 => "00100100",4699 => "00110000",4700 => "10001011",4701 => "00010010",4702 => "01100100",4703 => "01010111",4704 => "10011111",4705 => "10110000",4706 => "11011011",4707 => "10110000",4708 => "00111000",4709 => "11001011",4710 => "00101000",4711 => "00000110",4712 => "10110011",4713 => "11100001",4714 => "00011000",4715 => "00110011",4716 => "11100101",4717 => "10001011",4718 => "11110001",4719 => "11101101",4720 => "00101100",4721 => "01111110",4722 => "10110000",4723 => "10111000",4724 => "00011011",4725 => "11011011",4726 => "10000001",4727 => "01001001",4728 => "11111100",4729 => "00010010",4730 => "00000011",4731 => "11111010",4732 => "11010110",4733 => "01101010",4734 => "10100001",4735 => "01101010",4736 => "00101010",4737 => "01110110",4738 => "11100110",4739 => "11111011",4740 => "00011010",4741 => "00001010",4742 => "01100110",4743 => "10100000",4744 => "11111101",4745 => "11011000",4746 => "01110001",4747 => "10101001",4748 => "00110000",4749 => "10101101",4750 => "10110011",4751 => "01010100",4752 => "10100111",4753 => "11000011",4754 => "01111101",4755 => "01010111",4756 => "00000011",4757 => "00111100",4758 => "01010100",4759 => "10101000",4760 => "00101110",4761 => "10011110",4762 => "00011010",4763 => "10001001",4764 => "00011110",4765 => "10000100",4766 => "11101101",4767 => "00111100",4768 => "11110101",4769 => "11111000",4770 => "10010001",4771 => "11000001",4772 => "00011001",4773 => "00011111",4774 => "00110111",4775 => "10101110",4776 => "11010110",4777 => "11110000",4778 => "10010110",4779 => "00000001",4780 => "01010011",4781 => "10001011",4782 => "10101111",4783 => "01001011",4784 => "10111111",4785 => "01100001",4786 => "10110011",4787 => "00100110",4788 => "01000110",4789 => "01101010",4790 => "01101101",4791 => "10011110",4792 => "00100111",4793 => "00101101",4794 => "10110001",4795 => "10011110",4796 => "10011010",4797 => "11100010",4798 => "10001111",4799 => "10000000",4800 => "00100001",4801 => "00110010",4802 => "00010001",4803 => "01110000",4804 => "11000110",4805 => "01011001",4806 => "00010100",4807 => "10001101",4808 => "11011111",4809 => "00010110",4810 => "10010010",4811 => "10001000",4812 => "10001100",4813 => "01101001",4814 => "01100101",4815 => "10110100",4816 => "00010111",4817 => "10000010",4818 => "11000101",4819 => "00110001",4820 => "01111010",4821 => "10011110",4822 => "00110111",4823 => "10000101",4824 => "10010011",4825 => "00011010",4826 => "00111110",4827 => "00000110",4828 => "01101001",4829 => "11111000",4830 => "11111010",4831 => "11101111",4832 => "10011100",4833 => "11111001",4834 => "11010100",4835 => "01011001",4836 => "00000001",4837 => "01000100",4838 => "00010110",4839 => "11001100",4840 => "10100101",4841 => "10101011",4842 => "00111111",4843 => "11010111",4844 => "10110110",4845 => "00100110",4846 => "01101010",4847 => "10110011",4848 => "01011111",4849 => "00010000",4850 => "11000000",4851 => "11011000",4852 => "10100100",4853 => "11111100",4854 => "10100111",4855 => "00110111",4856 => "11101101",4857 => "10101010",4858 => "01010110",4859 => "10000111",4860 => "01101010",4861 => "01000011",4862 => "01001110",4863 => "10001111",4864 => "10111011",4865 => "01010111",4866 => "00001110",4867 => "01110001",4868 => "10101110",4869 => "11100011",4870 => "01000101",4871 => "10111001",4872 => "01101001",4873 => "00111001",4874 => "10100101",4875 => "10001001",4876 => "00010001",4877 => "00010011",4878 => "11100110",4879 => "01100011",4880 => "00111100",4881 => "00100101",4882 => "11001100",4883 => "00010111",4884 => "00001110",4885 => "00000001",4886 => "10101010",4887 => "11111100",4888 => "11100010",4889 => "00110100",4890 => "00110100",4891 => "01111101",4892 => "11101100",4893 => "00000000",4894 => "10101100",4895 => "00101101",4896 => "10010011",4897 => "01011111",4898 => "10010100",4899 => "01001111",4900 => "01000111",4901 => "10001110",4902 => "11110111",4903 => "11100011",4904 => "10001001",4905 => "00100110",4906 => "00111001",4907 => "00010011",4908 => "00010011",4909 => "10111101",4910 => "00100100",4911 => "00111001",4912 => "00101100",4913 => "10100011",4914 => "00011001",4915 => "11100101",4916 => "11000000",4917 => "11000011",4918 => "11001111",4919 => "11011110",4920 => "10000111",4921 => "00001001",4922 => "01110111",4923 => "01100110",4924 => "10001111",4925 => "01011100",4926 => "00010101",4927 => "10101110",4928 => "10011000",4929 => "10110100",4930 => "01001101",4931 => "11011110",4932 => "10101000",4933 => "11000110",4934 => "11001101",4935 => "11001011",4936 => "11011011",4937 => "11001110",4938 => "00111011",4939 => "10000000",4940 => "10101000",4941 => "00011111",4942 => "10101101",4943 => "11111111",4944 => "11011101",4945 => "10111110",4946 => "10011111",4947 => "01000100",4948 => "01000110",4949 => "10111001",4950 => "10111101",4951 => "10011111",4952 => "10001011",4953 => "00000011",4954 => "00110100",4955 => "01010001",4956 => "10100111",4957 => "00011111",4958 => "01100111",4959 => "00011111",4960 => "11100101",4961 => "01111011",4962 => "01100010",4963 => "01010010",4964 => "11001110",4965 => "01011110",4966 => "10000101",4967 => "11010110",4968 => "10000000",4969 => "11010000",4970 => "10111000",4971 => "11000011",4972 => "11001110",4973 => "10100100",4974 => "11001000",4975 => "11100011",4976 => "10110100",4977 => "00100100",4978 => "11011101",4979 => "10111110",4980 => "10011000",4981 => "00110110",4982 => "01110000",4983 => "11001110",4984 => "11011010",4985 => "11111110",4986 => "10111001",4987 => "01110010",4988 => "01110011",4989 => "00011000",4990 => "01011111",4991 => "00011101",4992 => "00010001",4993 => "11101110",4994 => "11000011",4995 => "00000000",4996 => "01100010",4997 => "10111111",4998 => "10110011",4999 => "01111101",5000 => "01101010",5001 => "10111110",5002 => "01000011",5003 => "00001001",5004 => "10110101",5005 => "10001000",5006 => "00110101",5007 => "01001000",5008 => "01001101",5009 => "00100010",5010 => "00101000",5011 => "11001011",5012 => "10101000",5013 => "00100001",5014 => "11110010",5015 => "10100001",5016 => "11011001",5017 => "10100101",5018 => "11101011",5019 => "10001100",5020 => "01000101",5021 => "00110101",5022 => "10111110",5023 => "10010010",5024 => "11100110",5025 => "11010110",5026 => "11111000",5027 => "01010000",5028 => "11101011",5029 => "11001101",5030 => "00100000",5031 => "00011011",5032 => "00101010",5033 => "10110001",5034 => "01100010",5035 => "00111100",5036 => "11101111",5037 => "00110110",5038 => "00110101",5039 => "00110000",5040 => "00001101",5041 => "10100011",5042 => "10010001",5043 => "11100011",5044 => "01011011",5045 => "11011001",5046 => "11010011",5047 => "01111101",5048 => "00101011",5049 => "10001000",5050 => "10001101",5051 => "11111011",5052 => "11101100",5053 => "00000111",5054 => "00100111",5055 => "11111111",5056 => "10001100",5057 => "00000001",5058 => "11010111",5059 => "01111110",5060 => "10100100",5061 => "11110011",5062 => "00010100",5063 => "10110111",5064 => "00101111",5065 => "10101100",5066 => "00001011",5067 => "10000110",5068 => "00101000",5069 => "01110010",5070 => "00100000",5071 => "10000010",5072 => "00000100",5073 => "10001100",5074 => "00101111",5075 => "01110011",5076 => "11101010",5077 => "01111010",5078 => "01011110",5079 => "01011000",5080 => "11010000",5081 => "10111010",5082 => "00001111",5083 => "10000110",5084 => "01110100",5085 => "00100100",5086 => "00001111",5087 => "01001000",5088 => "10101111",5089 => "00010111",5090 => "10011110",5091 => "10011011",5092 => "00110011",5093 => "11100100",5094 => "01000101",5095 => "11000010",5096 => "11110000",5097 => "10110101",5098 => "01011110",5099 => "00001101",5100 => "01111000",5101 => "11011110",5102 => "11101101",5103 => "10010011",5104 => "11000101",5105 => "01010010",5106 => "10110011",5107 => "11110010",5108 => "11101011",5109 => "10011010",5110 => "00001111",5111 => "11011100",5112 => "11100000",5113 => "00100001",5114 => "11111011",5115 => "01001001",5116 => "10010010",5117 => "00100011",5118 => "11100011",5119 => "00000110",5120 => "11110110",5121 => "11111011",5122 => "01011110",5123 => "00010110",5124 => "00101101",5125 => "01110001",5126 => "00001101",5127 => "11010000",5128 => "11100011",5129 => "10111010",5130 => "11101010",5131 => "01001011",5132 => "10001000",5133 => "11110100",5134 => "11101101",5135 => "10111010",5136 => "11111100",5137 => "10000000",5138 => "01110011",5139 => "10011011",5140 => "10110001",5141 => "01000100",5142 => "01110000",5143 => "00110101",5144 => "01001001",5145 => "11001101",5146 => "10000001",5147 => "11010101",5148 => "01110010",5149 => "01011001",5150 => "00110001",5151 => "11000010",5152 => "11001100",5153 => "10000101",5154 => "10010110",5155 => "01110001",5156 => "01000101",5157 => "11111111",5158 => "10010111",5159 => "01111001",5160 => "00011010",5161 => "00111110",5162 => "11110010",5163 => "01001010",5164 => "00100110",5165 => "10110010",5166 => "10111010",5167 => "10111100",5168 => "11111011",5169 => "11110100",5170 => "10010000",5171 => "00001110",5172 => "01111000",5173 => "10011101",5174 => "11100000",5175 => "11100010",5176 => "11011011",5177 => "11010010",5178 => "00001001",5179 => "01110100",5180 => "00001110",5181 => "10101110",5182 => "01000110",5183 => "11101010",5184 => "11011111",5185 => "00000100",5186 => "01010011",5187 => "11100110",5188 => "01000101",5189 => "01100111",5190 => "11011100",5191 => "00011111",5192 => "01001111",5193 => "00010111",5194 => "11011010",5195 => "11000000",5196 => "11000110",5197 => "00101001",5198 => "10110111",5199 => "01000011",5200 => "01011000",5201 => "10001011",5202 => "11110111",5203 => "11111100",5204 => "10101110",5205 => "01000001",5206 => "10011010",5207 => "11010101",5208 => "00011100",5209 => "00001110",5210 => "10000111",5211 => "01101011",5212 => "11101101",5213 => "00101110",5214 => "01000011",5215 => "11111011",5216 => "10001000",5217 => "01011101",5218 => "01001010",5219 => "11010000",5220 => "01100011",5221 => "11001001",5222 => "11000101",5223 => "11111000",5224 => "11000011",5225 => "11100101",5226 => "10010011",5227 => "01000001",5228 => "10001101",5229 => "11100011",5230 => "00101101",5231 => "00001111",5232 => "01110111",5233 => "11010010",5234 => "01000001",5235 => "11100001",5236 => "10010010",5237 => "10101011",5238 => "10101110",5239 => "01010001",5240 => "00011011",5241 => "10111111",5242 => "11111100",5243 => "11100110",5244 => "11000011",5245 => "11000001",5246 => "01100010",5247 => "01010110",5248 => "11100110",5249 => "10101011",5250 => "01111011",5251 => "00100000",5252 => "10110001",5253 => "11111010",5254 => "10111101",5255 => "01011000",5256 => "00100011",5257 => "11010011",5258 => "10100101",5259 => "00111100",5260 => "00011001",5261 => "00011001",5262 => "01111000",5263 => "00101100",5264 => "01110110",5265 => "00010001",5266 => "10111011",5267 => "00010111",5268 => "01000000",5269 => "00101001",5270 => "11010111",5271 => "11001111",5272 => "10000110",5273 => "01101001",5274 => "00000101",5275 => "11101100",5276 => "01110111",5277 => "01100011",5278 => "11110101",5279 => "10111010",5280 => "10110110",5281 => "00010011",5282 => "11111101",5283 => "10001111",5284 => "00001010",5285 => "00000010",5286 => "00010001",5287 => "00010010",5288 => "00110001",5289 => "00100000",5290 => "10011000",5291 => "10001001",5292 => "01011010",5293 => "00110011",5294 => "10001101",5295 => "10010100",5296 => "10100000",5297 => "00100000",5298 => "10111000",5299 => "00011000",5300 => "11110101",5301 => "10011000",5302 => "10110000",5303 => "10110100",5304 => "00001111",5305 => "01101000",5306 => "00010001",5307 => "01011101",5308 => "10001010",5309 => "11110101",5310 => "10001100",5311 => "10100000",5312 => "00010101",5313 => "01010101",5314 => "11010001",5315 => "01110010",5316 => "01101111",5317 => "10001001",5318 => "01010111",5319 => "10110111",5320 => "00111110",5321 => "01011000",5322 => "00100100",5323 => "11001111",5324 => "11100110",5325 => "00000000",5326 => "11010001",5327 => "01110011",5328 => "11000000",5329 => "11001110",5330 => "10110110",5331 => "01100111",5332 => "01000101",5333 => "00101000",5334 => "00111111",5335 => "11011110",5336 => "00101100",5337 => "00111111",5338 => "00100000",5339 => "10110010",5340 => "00100000",5341 => "00001110",5342 => "00000011",5343 => "00011111",5344 => "11001111",5345 => "01110111",5346 => "10101101",5347 => "00000010",5348 => "11100110",5349 => "11100001",5350 => "10100000",5351 => "01101000",5352 => "10111101",5353 => "00010101",5354 => "10111010",5355 => "00110101",5356 => "11101111",5357 => "10110110",5358 => "00001001",5359 => "10110001",5360 => "00010111",5361 => "10101011",5362 => "01001111",5363 => "11110010",5364 => "11101100",5365 => "01111100",5366 => "10001100",5367 => "10000011",5368 => "10000000",5369 => "10010100",5370 => "00111010",5371 => "00111011",5372 => "11100100",5373 => "01100110",5374 => "00101001",5375 => "11100111",5376 => "00100101",5377 => "11000110",5378 => "00011001",5379 => "10000001",5380 => "10101001",5381 => "00101101",5382 => "10001100",5383 => "11101110",5384 => "11110010",5385 => "00000100",5386 => "10001000",5387 => "01110110",5388 => "01100010",5389 => "10000010",5390 => "01110000",5391 => "01100101",5392 => "10011000",5393 => "00110011",5394 => "10110000",5395 => "01111010",5396 => "01110010",5397 => "11011001",5398 => "11100011",5399 => "00110011",5400 => "10111011",5401 => "11000111",5402 => "00000011",5403 => "01010001",5404 => "01000011",5405 => "00001011",5406 => "01111001",5407 => "11010010",5408 => "00001001",5409 => "00100110",5410 => "01111100",5411 => "01111101",5412 => "10101000",5413 => "11001100",5414 => "10001100",5415 => "01111101",5416 => "00101001",5417 => "00100111",5418 => "01111110",5419 => "01010111",5420 => "00011011",5421 => "01001011",5422 => "11111110",5423 => "10011100",5424 => "10111010",5425 => "10001010",5426 => "01010000",5427 => "00000010",5428 => "00011001",5429 => "00000001",5430 => "01111000",5431 => "10000111",5432 => "01110000",5433 => "10111001",5434 => "01101001",5435 => "01111011",5436 => "11101100",5437 => "11101101",5438 => "01101100",5439 => "01100011",5440 => "00011000",5441 => "11010110",5442 => "00010000",5443 => "00011011",5444 => "01000111",5445 => "01001100",5446 => "10111100",5447 => "10101111",5448 => "11010110",5449 => "10000011",5450 => "00100010",5451 => "10100011",5452 => "01100010",5453 => "10100001",5454 => "01110001",5455 => "00000000",5456 => "00100001",5457 => "10110000",5458 => "11111001",5459 => "00100011",5460 => "11001101",5461 => "11011000",5462 => "01111110",5463 => "10000100",5464 => "00111010",5465 => "10100110",5466 => "10010010",5467 => "10110100",5468 => "10110011",5469 => "10111010",5470 => "11111101",5471 => "11110011",5472 => "11100011",5473 => "00101111",5474 => "01001100",5475 => "00101111",5476 => "10010100",5477 => "00110100",5478 => "00001011",5479 => "01110001",5480 => "00101100",5481 => "00011010",5482 => "00111100",5483 => "11011000",5484 => "10100010",5485 => "01000000",5486 => "00101010",5487 => "00001110",5488 => "01011000",5489 => "10101011",5490 => "00100111",5491 => "11101001",5492 => "11111010",5493 => "00001101",5494 => "01111001",5495 => "10111011",5496 => "01000111",5497 => "11011110",5498 => "01101000",5499 => "11100011",5500 => "11101101",5501 => "10000101",5502 => "11010001",5503 => "01100100",5504 => "01000111",5505 => "00000101",5506 => "00011101",5507 => "01001100",5508 => "01100111",5509 => "11111010",5510 => "01000000",5511 => "10001110",5512 => "00110100",5513 => "11011011",5514 => "01000110",5515 => "01011101",5516 => "11100100",5517 => "11100111",5518 => "10010011",5519 => "01101000",5520 => "00111000",5521 => "01001100",5522 => "11010101",5523 => "11000011",5524 => "11111010",5525 => "10101011",5526 => "11110001",5527 => "01101111",5528 => "01011011",5529 => "00011111",5530 => "10101110",5531 => "11101101",5532 => "00011000",5533 => "01011100",5534 => "00100101",5535 => "01101000",5536 => "01111010",5537 => "00111101",5538 => "10100110",5539 => "10100010",5540 => "11001110",5541 => "01101100",5542 => "11101111",5543 => "10110011",5544 => "00010000",5545 => "00001001",5546 => "10010001",5547 => "00010101",5548 => "00110001",5549 => "01011000",5550 => "00111100",5551 => "01110100",5552 => "01010100",5553 => "11000110",5554 => "11110100",5555 => "01111010",5556 => "10111011",5557 => "00100011",5558 => "00001100",5559 => "11111001",5560 => "11001100",5561 => "01000101",5562 => "10001001",5563 => "00010000",5564 => "11111001",5565 => "01100000",5566 => "01110110",5567 => "00111011",5568 => "11111111",5569 => "01101101",5570 => "10001100",5571 => "11010000",5572 => "10101111",5573 => "00101111",5574 => "10110111",5575 => "00111111",5576 => "10001101",5577 => "10000010",5578 => "00011110",5579 => "00101111",5580 => "10000010",5581 => "00110100",5582 => "01100001",5583 => "10100010",5584 => "01010001",5585 => "00100110",5586 => "01001100",5587 => "10101011",5588 => "11011011",5589 => "11011101",5590 => "00101101",5591 => "10110100",5592 => "11011110",5593 => "10101011",5594 => "00101011",5595 => "11101100",5596 => "10100011",5597 => "10111100",5598 => "10000011",5599 => "00100000",5600 => "11011101",5601 => "10101100",5602 => "10100111",5603 => "10111010",5604 => "00100110",5605 => "10010111",5606 => "11100100",5607 => "11111111",5608 => "00101001",5609 => "10100110",5610 => "11000000",5611 => "10000000",5612 => "00000011",5613 => "11100000",5614 => "11011110",5615 => "11101110",5616 => "00110000",5617 => "10000101",5618 => "01000011",5619 => "10011001",5620 => "11000001",5621 => "10011100",5622 => "10011011",5623 => "10010000",5624 => "00101000",5625 => "11000101",5626 => "11011010",5627 => "11111111",5628 => "00111111",5629 => "01010110",5630 => "00111011",5631 => "10111100",5632 => "01100101",5633 => "01110100",5634 => "10101010",5635 => "01110101",5636 => "00010110",5637 => "11101010",5638 => "11010001",5639 => "00010001",5640 => "00110100",5641 => "11011001",5642 => "10101110",5643 => "11001001",5644 => "00100111",5645 => "11010111",5646 => "00111000",5647 => "11111011",5648 => "00100011",5649 => "01010010",5650 => "01001001",5651 => "11001100",5652 => "01011000",5653 => "00101110",5654 => "11111110",5655 => "11111011",5656 => "01100000",5657 => "00111100",5658 => "10011010",5659 => "11100101",5660 => "00110100",5661 => "11000000",5662 => "00111111",5663 => "00111110",5664 => "11111101",5665 => "11111101",5666 => "01100000",5667 => "01001000",5668 => "11100001",5669 => "01100000",5670 => "11001110",5671 => "00100101",5672 => "01001000",5673 => "01011000",5674 => "11001011",5675 => "01010100",5676 => "10011110",5677 => "01010111",5678 => "11100011",5679 => "00110010",5680 => "10101010",5681 => "00010110",5682 => "00100001",5683 => "00100100",5684 => "01001001",5685 => "00011010",5686 => "01001110",5687 => "10000001",5688 => "00101100",5689 => "11001011",5690 => "10001100",5691 => "00000100",5692 => "11101001",5693 => "10100101",5694 => "00000010",5695 => "00011000",5696 => "01101010",5697 => "10001110",5698 => "01001111",5699 => "00010100",5700 => "01110010",5701 => "11110010",5702 => "00101100",5703 => "10100011",5704 => "11101001",5705 => "10010000",5706 => "00100101",5707 => "00001000",5708 => "01000101",5709 => "01100111",5710 => "00100011",5711 => "01000000",5712 => "01011000",5713 => "01010110",5714 => "01001000",5715 => "10011001",5716 => "11010010",5717 => "11011011",5718 => "10011110",5719 => "00100100",5720 => "10111001",5721 => "10100000",5722 => "11100101",5723 => "01000111",5724 => "00100001",5725 => "10011111",5726 => "11110011",5727 => "11010111",5728 => "11110010",5729 => "10100110",5730 => "01111111",5731 => "00001001",5732 => "01110111",5733 => "11110000",5734 => "11000000",5735 => "00010100",5736 => "11000110",5737 => "10101011",5738 => "00010100",5739 => "11100100",5740 => "01001010",5741 => "00000011",5742 => "00101111",5743 => "01101001",5744 => "11011011",5745 => "01100111",5746 => "01110011",5747 => "01010110",5748 => "11101111",5749 => "00010000",5750 => "00110000",5751 => "01010000",5752 => "01100101",5753 => "11011111",5754 => "01011110",5755 => "10001000",5756 => "01111110",5757 => "01110101",5758 => "10011100",5759 => "00011101",5760 => "10110111",5761 => "10110111",5762 => "01010101",5763 => "11100101",5764 => "10110110",5765 => "01110111",5766 => "00011011",5767 => "10111101",5768 => "01010000",5769 => "00100010",5770 => "01001010",5771 => "11000101",5772 => "11100111",5773 => "10111110",5774 => "11100010",5775 => "01101000",5776 => "10100011",5777 => "01011001",5778 => "00111011",5779 => "01110101",5780 => "01000110",5781 => "11111011",5782 => "00000010",5783 => "11111000",5784 => "01011000",5785 => "01001111",5786 => "00000110",5787 => "00000000",5788 => "00010001",5789 => "11101000",5790 => "00100010",5791 => "00000011",5792 => "10010001",5793 => "11011110",5794 => "10011111",5795 => "01110000",5796 => "00101111",5797 => "01001011",5798 => "00000000",5799 => "01011001",5800 => "01000101",5801 => "01011110",5802 => "01110101",5803 => "00101110",5804 => "00101011",5805 => "01110110",5806 => "01101010",5807 => "10110010",5808 => "10111001",5809 => "10111110",5810 => "10110101",5811 => "01001100",5812 => "11000100",5813 => "00111011",5814 => "10110000",5815 => "10010001",5816 => "01110110",5817 => "10110001",5818 => "01111100",5819 => "01101000",5820 => "11101101",5821 => "11010111",5822 => "11101011",5823 => "10101000",5824 => "10111011",5825 => "10010111",5826 => "10110101",5827 => "01110001",5828 => "01010010",5829 => "01011101",5830 => "10001001",5831 => "10111010",5832 => "01111111",5833 => "00000000",5834 => "00101110",5835 => "11101010",5836 => "11010110",5837 => "01011111",5838 => "10010011",5839 => "11001000",5840 => "11001111",5841 => "11101001",5842 => "01000001",5843 => "11011010",5844 => "11001010",5845 => "00001100",5846 => "01001100",5847 => "01101111",5848 => "10100100",5849 => "11100000",5850 => "11110001",5851 => "10111111",5852 => "00101101",5853 => "01001100",5854 => "10001110",5855 => "11101101",5856 => "01010110",5857 => "00101100",5858 => "00111101",5859 => "10100110",5860 => "00000011",5861 => "01011010",5862 => "10110100",5863 => "00110110",5864 => "10101001",5865 => "01000110",5866 => "11010110",5867 => "10101100",5868 => "00001001",5869 => "10011110",5870 => "01110110",5871 => "01010000",5872 => "00011000",5873 => "11111000",5874 => "10101001",5875 => "11101010",5876 => "11101100",5877 => "01010001",5878 => "10111101",5879 => "01000001",5880 => "10001101",5881 => "11111010",5882 => "10110001",5883 => "11000000",5884 => "00110100",5885 => "10111101",5886 => "11111000",5887 => "10001101",5888 => "11111001",5889 => "01100010",5890 => "00110001",5891 => "11111011",5892 => "11101001",5893 => "10101100",5894 => "00000100",5895 => "10011100",5896 => "01101111",5897 => "00010011",5898 => "00011111",5899 => "00000100",5900 => "11001101",5901 => "10001010",5902 => "00010110",5903 => "00011110",5904 => "10001101",5905 => "11111011",5906 => "01010111",5907 => "01000110",5908 => "00010011",5909 => "00000011",5910 => "00011001",5911 => "01010110",5912 => "11011000",5913 => "00101001",5914 => "11010111",5915 => "10101001",5916 => "10110100",5917 => "10101101",5918 => "10101110",5919 => "01101101",5920 => "10111010",5921 => "00111011",5922 => "00010010",5923 => "10000111",5924 => "10000111",5925 => "10000000",5926 => "11111101",5927 => "11010011",5928 => "10011100",5929 => "10011101",5930 => "10100101",5931 => "11111001",5932 => "10010001",5933 => "01110100",5934 => "10101000",5935 => "00011101",5936 => "01000110",5937 => "01100100",5938 => "01101100",5939 => "10011010",5940 => "11110000",5941 => "01110001",5942 => "01111111",5943 => "01110101",5944 => "10001100",5945 => "00001110",5946 => "11111000",5947 => "00010010",5948 => "11011101",5949 => "10110101",5950 => "10101111",5951 => "00011010",5952 => "10111010",5953 => "00101001",5954 => "01101011",5955 => "01110111",5956 => "10000010",5957 => "00110000",5958 => "10011011",5959 => "01001001",5960 => "01111011",5961 => "11000010",5962 => "01011101",5963 => "10101011",5964 => "10110110",5965 => "00001010",5966 => "01001100",5967 => "11101011",5968 => "01010111",5969 => "10000001",5970 => "01110100",5971 => "10000100",5972 => "00000000",5973 => "00001010",5974 => "01000000",5975 => "10000100",5976 => "01111111",5977 => "11100000",5978 => "11111111",5979 => "11010000",5980 => "10111101",5981 => "11010001",5982 => "10111101",5983 => "10110111",5984 => "11100000",5985 => "01010110",5986 => "01111001",5987 => "10111011",5988 => "00001011",5989 => "11010010",5990 => "01010110",5991 => "01100010",5992 => "11100100",5993 => "01110001",5994 => "01111100",5995 => "01011100",5996 => "10111111",5997 => "01010011",5998 => "10011100",5999 => "00100111",6000 => "10011010",6001 => "00001011",6002 => "00000000",6003 => "01110001",6004 => "01110001",6005 => "11000010",6006 => "00101010",6007 => "11110001",6008 => "11001111",6009 => "10110101",6010 => "10100111",6011 => "10011101",6012 => "00001000",6013 => "00100110",6014 => "10111111",6015 => "01101001",6016 => "00101101",6017 => "10010101",6018 => "01100001",6019 => "11101010",6020 => "11101100",6021 => "11011010",6022 => "10110011",6023 => "00000101",6024 => "11000000",6025 => "01010111",6026 => "00000011",6027 => "11011011",6028 => "10001010",6029 => "01011010",6030 => "01101111",6031 => "01100000",6032 => "10100011",6033 => "01101011",6034 => "01011010",6035 => "01111010",6036 => "11001110",6037 => "10101101",6038 => "00001111",6039 => "11100111",6040 => "10001110",6041 => "11101101",6042 => "00010000",6043 => "01111110",6044 => "10010011",6045 => "01011101",6046 => "00010100",6047 => "00110000",6048 => "10111111",6049 => "11001000",6050 => "00000111",6051 => "00110100",6052 => "11011101",6053 => "10110000",6054 => "00011100",6055 => "01110000",6056 => "11110101",6057 => "10001010",6058 => "01001011",6059 => "00101011",6060 => "01100000",6061 => "00000000",6062 => "01000110",6063 => "10000100",6064 => "11000011",6065 => "10110100",6066 => "00011001",6067 => "00111010",6068 => "10100001",6069 => "00010011",6070 => "01110001",6071 => "01010001",6072 => "11110011",6073 => "11011010",6074 => "10001111",6075 => "11101011",6076 => "01100111",6077 => "01000011",6078 => "10011011",6079 => "11010101",6080 => "10101101",6081 => "11101000",6082 => "11111110",6083 => "10000010",6084 => "00010011",6085 => "10000101",6086 => "00111101",6087 => "01001101",6088 => "01011101",6089 => "00010000",6090 => "11110001",6091 => "11011101",6092 => "01010010",6093 => "00000100",6094 => "01000100",6095 => "11101000",6096 => "01000010",6097 => "11101010",6098 => "00010100",6099 => "01111100",6100 => "11111101",6101 => "01110111",6102 => "01101111",6103 => "01011101",6104 => "10000111",6105 => "10101011",6106 => "10100111",6107 => "10010110",6108 => "01011010",6109 => "01110011",6110 => "01101110",6111 => "11010010",6112 => "00001100",6113 => "00110001",6114 => "10100010",6115 => "11000101",6116 => "00000100",6117 => "01111011",6118 => "00111111",6119 => "01001000",6120 => "01111111",6121 => "10001100",6122 => "10000100",6123 => "11001100",6124 => "01001001",6125 => "10100001",6126 => "10111001",6127 => "11111110",6128 => "10001001",6129 => "01011011",6130 => "11111001",6131 => "10000001",6132 => "01000001",6133 => "00101110",6134 => "01111001",6135 => "00010001",6136 => "01011001",6137 => "10010000",6138 => "10100101",6139 => "00100101",6140 => "01101000",6141 => "10000100",6142 => "11101111",6143 => "11101100",6144 => "10101001",6145 => "00001000",6146 => "10111111",6147 => "11000110",6148 => "11111111",6149 => "10011000",6150 => "00011011",6151 => "00000010",6152 => "10010111",6153 => "01110010",6154 => "10110100",6155 => "00111101",6156 => "01011110",6157 => "10010001",6158 => "11011111",6159 => "11001000",6160 => "10010110",6161 => "11010001",6162 => "01100111",6163 => "11111001",6164 => "10000110",6165 => "01101001",6166 => "00000110",6167 => "00101001",6168 => "10111111",6169 => "01001100",6170 => "10010101",6171 => "01000101",6172 => "01101011",6173 => "10011110",6174 => "10000000",6175 => "10101001",6176 => "11001000",6177 => "10000101",6178 => "11010001",6179 => "01000101",6180 => "11110110",6181 => "01110110",6182 => "01000101",6183 => "00100001",6184 => "01100101",6185 => "00111010",6186 => "01100001",6187 => "11000100",6188 => "11111000",6189 => "10110100",6190 => "10100110",6191 => "11110001",6192 => "10110011",6193 => "00001011",6194 => "01111100",6195 => "00011101",6196 => "00101011",6197 => "01011010",6198 => "00100000",6199 => "11110111",6200 => "10101011",6201 => "00111001",6202 => "10010001",6203 => "10001011",6204 => "11101011",6205 => "11100111",6206 => "00011110",6207 => "00010111",6208 => "11100100",6209 => "11000011",6210 => "00010111",6211 => "00111111",6212 => "11010001",6213 => "10100101",6214 => "00001100",6215 => "00110111",6216 => "01100011",6217 => "01111110",6218 => "11011010",6219 => "10101001",6220 => "00100001",6221 => "00110100",6222 => "11000011",6223 => "11000111",6224 => "00001111",6225 => "00111111",6226 => "01000101",6227 => "11110000",6228 => "01000001",6229 => "11011000",6230 => "10111101",6231 => "01001111",6232 => "00010101",6233 => "01010001",6234 => "11001011",6235 => "00111011",6236 => "11110111",6237 => "11100000",6238 => "10010000",6239 => "00110100",6240 => "01110001",6241 => "00010000",6242 => "01111110",6243 => "01001010",6244 => "10111000",6245 => "01101010",6246 => "01011101",6247 => "11010101",6248 => "10011010",6249 => "10101011",6250 => "01011000",6251 => "01111000",6252 => "10110000",6253 => "00100101",6254 => "11001110",6255 => "10011110",6256 => "10110101",6257 => "11010001",6258 => "11110011",6259 => "11110011",6260 => "10000101",6261 => "11011001",6262 => "00110010",6263 => "11000110",6264 => "10101110",6265 => "10110110",6266 => "10000101",6267 => "11111011",6268 => "11000110",6269 => "00111100",6270 => "11100101",6271 => "10000100",6272 => "01111111",6273 => "10001011",6274 => "10101011",6275 => "00100001",6276 => "11011000",6277 => "11011100",6278 => "01010000",6279 => "00011000",6280 => "01110110",6281 => "11101001",6282 => "10101001",6283 => "10000110",6284 => "10000110",6285 => "01110001",6286 => "11010111",6287 => "01100010",6288 => "11100101",6289 => "00011000",6290 => "01011111",6291 => "01010101",6292 => "00100010",6293 => "10010000",6294 => "11101011",6295 => "10101111",6296 => "01001011",6297 => "00001011",6298 => "00001011",6299 => "01110100",6300 => "10001100",6301 => "01110001",6302 => "10110101",6303 => "00010111",6304 => "10000101",6305 => "10010100",6306 => "01110101",6307 => "01110011",6308 => "10101000",6309 => "01100111",6310 => "00000100",6311 => "10100010",6312 => "01010101",6313 => "10001111",6314 => "10000101",6315 => "10111101",6316 => "00110000",6317 => "01110000",6318 => "11111000",6319 => "11000100",6320 => "00010001",6321 => "01111111",6322 => "01010100",6323 => "11001010",6324 => "11101110",6325 => "11000101",6326 => "00000101",6327 => "00100101",6328 => "10010110",6329 => "01011101",6330 => "01001010",6331 => "10110101",6332 => "01101011",6333 => "11011000",6334 => "00010011",6335 => "10100100",6336 => "00110001",6337 => "00100000",6338 => "10011110",6339 => "11010001",6340 => "01011110",6341 => "10010110",6342 => "10001110",6343 => "10111010",6344 => "01100000",6345 => "10111010",6346 => "01000010",6347 => "10000011",6348 => "10010101",6349 => "11011010",6350 => "01101010",6351 => "10101100",6352 => "10010011",6353 => "01011000",6354 => "10001000",6355 => "00110001",6356 => "01100001",6357 => "10110000",6358 => "11111001",6359 => "11111101",6360 => "01111100",6361 => "00000100",6362 => "10101101",6363 => "11100000",6364 => "01111011",6365 => "01011010",6366 => "01111001",6367 => "00110100",6368 => "11111100",6369 => "01001100",6370 => "01111100",6371 => "10111100",6372 => "10011101",6373 => "11011011",6374 => "11111111",6375 => "11000100",6376 => "00010011",6377 => "00110000",6378 => "01101010",6379 => "10101111",6380 => "00011101",6381 => "01001000",6382 => "10101001",6383 => "11000001",6384 => "01111100",6385 => "00011110",6386 => "10000011",6387 => "10100110",6388 => "11000001",6389 => "11101001",6390 => "10011110",6391 => "10000111",6392 => "11000011",6393 => "11000110",6394 => "01000011",6395 => "10111110",6396 => "10011001",6397 => "00101111",6398 => "01100011",6399 => "01010000",6400 => "11001110",6401 => "10110100",6402 => "01110101",6403 => "00001110",6404 => "01000101",6405 => "10000101",6406 => "00011011",6407 => "10110110",6408 => "01011010",6409 => "00010000",6410 => "00001101",6411 => "01010011",6412 => "10011110",6413 => "01100111",6414 => "00001000",6415 => "10011111",6416 => "00110010",6417 => "11011010",6418 => "10100011",6419 => "01101101",6420 => "00111110",6421 => "00111110",6422 => "01001110",6423 => "11011100",6424 => "11001001",6425 => "10011101",6426 => "00001111",6427 => "00011010",6428 => "11010000",6429 => "10011010",6430 => "11111100",6431 => "10111011",6432 => "01010100",6433 => "10110100",6434 => "00110110",6435 => "11101110",6436 => "00010010",6437 => "11010100",6438 => "01010001",6439 => "11001101",6440 => "01100101",6441 => "01001110",6442 => "11111111",6443 => "00100011",6444 => "11000100",6445 => "10101000",6446 => "00100101",6447 => "00100001",6448 => "00100000",6449 => "10100011",6450 => "10111111",6451 => "00100000",6452 => "00010111",6453 => "01011100",6454 => "11100001",6455 => "10011000",6456 => "00010001",6457 => "11011010",6458 => "10101001",6459 => "01010001",6460 => "01001110",6461 => "11001101",6462 => "01010100",6463 => "00111101",6464 => "10011111",6465 => "11101001",6466 => "11000000",6467 => "10001000",6468 => "01011001",6469 => "10110101",6470 => "01101110",6471 => "01101010",6472 => "01100001",6473 => "11000110",6474 => "01111001",6475 => "00000101",6476 => "00111111",6477 => "10111001",6478 => "01111000",6479 => "00001100",6480 => "10111100",6481 => "01101010",6482 => "01101100",6483 => "11001111",6484 => "10111001",6485 => "01001110",6486 => "01111001",6487 => "11110000",6488 => "10000100",6489 => "11010010",6490 => "10001111",6491 => "11001001",6492 => "11000000",6493 => "01000001",6494 => "01001000",6495 => "00101000",6496 => "10111001",6497 => "00110011",6498 => "00000011",6499 => "11110000",6500 => "00100011",6501 => "10111101",6502 => "10011111",6503 => "11010110",6504 => "11100101",6505 => "00101111",6506 => "01010000",6507 => "10000010",6508 => "11000011",6509 => "11011100",6510 => "11010100",6511 => "01110011",6512 => "11100100",6513 => "00110011",6514 => "00111011",6515 => "01011011",6516 => "10001110",6517 => "00010110",6518 => "01111001",6519 => "10000010",6520 => "11110001",6521 => "10100001",6522 => "11101001",6523 => "01000001",6524 => "11101101",6525 => "10101001",6526 => "11001010",6527 => "10000000",6528 => "10000110",6529 => "10001001",6530 => "01101001",6531 => "11100101",6532 => "11100011",6533 => "10011101",6534 => "11100111",6535 => "11001110",6536 => "11110010",6537 => "01001011",6538 => "10011111",6539 => "00101110",6540 => "01010000",6541 => "10001001",6542 => "01101010",6543 => "11111110",6544 => "10010000",6545 => "00001001",6546 => "01111010",6547 => "01110110",6548 => "11111001",6549 => "01111110",6550 => "01010011",6551 => "00010100",6552 => "01101001",6553 => "11011011",6554 => "01011110",6555 => "00101010",6556 => "00001000",6557 => "11100000",6558 => "01101001",6559 => "00100100",6560 => "10011111",6561 => "10100101",6562 => "11011101",6563 => "10010100",6564 => "00111100",6565 => "00001111",6566 => "01011111",6567 => "10011111",6568 => "10000000",6569 => "00101000",6570 => "10001010",6571 => "11111100",6572 => "01101101",6573 => "11010111",6574 => "01000011",6575 => "10010111",6576 => "10111011",6577 => "10110011",6578 => "00001011",6579 => "11011101",6580 => "01010001",6581 => "11011100",6582 => "11010111",6583 => "01011001",6584 => "11100001",6585 => "10000111",6586 => "10010000",6587 => "10100011",6588 => "00111010",6589 => "00010110",6590 => "01000100",6591 => "00001101",6592 => "00111011",6593 => "11111010",6594 => "10111110",6595 => "00001011",6596 => "00100110",6597 => "10110101",6598 => "00101011",6599 => "01111000",6600 => "10000011",6601 => "10011100",6602 => "00000110",6603 => "00010010",6604 => "10100110",6605 => "00101111",6606 => "01100001",6607 => "00000010",6608 => "00110011",6609 => "00011011",6610 => "10000101",6611 => "10100010",6612 => "00110111",6613 => "10110100",6614 => "00000000",6615 => "10000100",6616 => "11111111",6617 => "11101100",6618 => "01101101",6619 => "00101011",6620 => "10001110",6621 => "01111101",6622 => "00011011",6623 => "11001001",6624 => "11111001",6625 => "01010001",6626 => "10111010",6627 => "00010010",6628 => "01100111",6629 => "10001000",6630 => "00001001",6631 => "11101001",6632 => "01111000",6633 => "01111010",6634 => "11010010",6635 => "01011101",6636 => "11000100",6637 => "00000100",6638 => "00100111",6639 => "11001101",6640 => "00001101",6641 => "10100110",6642 => "10111000",6643 => "01101011",6644 => "01110011",6645 => "01010010",6646 => "10001111",6647 => "10000000",6648 => "00011001",6649 => "00101100",6650 => "11011100",6651 => "10110101",6652 => "10011100",6653 => "10101011",6654 => "10101100",6655 => "10101000",6656 => "11101110",6657 => "00000100",6658 => "11001101",6659 => "10111000",6660 => "10101111",6661 => "10001111",6662 => "00011001",6663 => "00001011",6664 => "00010000",6665 => "10000101",6666 => "00011111",6667 => "10110011",6668 => "11111100",6669 => "00100111",6670 => "01010101",6671 => "10100111",6672 => "01100100",6673 => "01100010",6674 => "10001011",6675 => "01110110",6676 => "10000100",6677 => "11101011",6678 => "00110110",6679 => "11110011",6680 => "01000111",6681 => "11011100",6682 => "01111001",6683 => "00100011",6684 => "10111100",6685 => "11011100",6686 => "01001101",6687 => "11001111",6688 => "11111011",6689 => "10110010",6690 => "10011001",6691 => "11010110",6692 => "11110100",6693 => "01000000",6694 => "11101111",6695 => "00100111",6696 => "10101011",6697 => "10100111",6698 => "01011101",6699 => "10011111",6700 => "10100010",6701 => "10100100",6702 => "10011001",6703 => "01010000",6704 => "11101000",6705 => "11110111",6706 => "00001111",6707 => "10100000",6708 => "10101011",6709 => "00111011",6710 => "10010000",6711 => "01010001",6712 => "01100010",6713 => "01001001",6714 => "11110101",6715 => "00010101",6716 => "01110111",6717 => "01100001",6718 => "11000101",6719 => "10010001",6720 => "10101000",6721 => "00001001",6722 => "10100001",6723 => "01101011",6724 => "11001100",6725 => "01001010",6726 => "00101100",6727 => "11101110",6728 => "10011011",6729 => "11010101",6730 => "00100111",6731 => "01100111",6732 => "10001011",6733 => "01100011",6734 => "11110010",6735 => "00100001",6736 => "01110000",6737 => "11010111",6738 => "11101110",6739 => "00110001",6740 => "11010001",6741 => "11000111",6742 => "10101011",6743 => "10110000",6744 => "10100001",6745 => "00100111",6746 => "11010000",6747 => "10101010",6748 => "10110011",6749 => "01110010",6750 => "01101101",6751 => "01101010",6752 => "11010110",6753 => "10001110",6754 => "00101000",6755 => "00011010",6756 => "01110000",6757 => "00100100",6758 => "10011011",6759 => "10111010",6760 => "11001100",6761 => "10101001",6762 => "10001001",6763 => "11001110",6764 => "10000011",6765 => "00000000",6766 => "00101100",6767 => "10100101",6768 => "01110101",6769 => "00011101",6770 => "11111110",6771 => "01101101",6772 => "01110000",6773 => "01000110",6774 => "00001110",6775 => "00000010",6776 => "01111010",6777 => "10010101",6778 => "01010000",6779 => "00000010",6780 => "10000010",6781 => "01100100",6782 => "01101101",6783 => "01010101",6784 => "01100101",6785 => "11111101",6786 => "10110011",6787 => "00100100",6788 => "01011001",6789 => "01001101",6790 => "11011101",6791 => "11010101",6792 => "00100101",6793 => "11100001",6794 => "10001001",6795 => "10110010",6796 => "10110100",6797 => "11010001",6798 => "00110110",6799 => "11110001",6800 => "01001010",6801 => "11110011",6802 => "00100010",6803 => "11001101",6804 => "10000010",6805 => "01001010",6806 => "10010110",6807 => "00101101",6808 => "10101101",6809 => "01110100",6810 => "00010110",6811 => "00010100",6812 => "00110100",6813 => "11011110",6814 => "10110100",6815 => "01110001",6816 => "10100000",6817 => "00011001",6818 => "00101011",6819 => "11010010",6820 => "11000111",6821 => "11110001",6822 => "11011001",6823 => "00000001",6824 => "11010110",6825 => "01101010",6826 => "10010101",6827 => "11011110",6828 => "11101110",6829 => "01000111",6830 => "01011101",6831 => "10001010",6832 => "00100110",6833 => "00100111",6834 => "10000111",6835 => "01010001",6836 => "11010111",6837 => "10101010",6838 => "10001101",6839 => "01100110",6840 => "10010100",6841 => "00011001",6842 => "00010010",6843 => "01100011",6844 => "00011111",6845 => "11000101",6846 => "00011111",6847 => "10010001",6848 => "10011101",6849 => "10010101",6850 => "00101101",6851 => "01011010",6852 => "01110000",6853 => "00001010",6854 => "11111101",6855 => "11001000",6856 => "00110000",6857 => "10000000",6858 => "10101100",6859 => "01000010",6860 => "10110000",6861 => "01111101",6862 => "00000100",6863 => "01100010",6864 => "10001000",6865 => "10111011",6866 => "10001000",6867 => "01100111",6868 => "11110000",6869 => "10001010",6870 => "11011101",6871 => "01100001",6872 => "00100110",6873 => "11010100",6874 => "10001101",6875 => "11010101",6876 => "11111001",6877 => "11010110",6878 => "00000110",6879 => "11001011",6880 => "00101110",6881 => "11101111",6882 => "10000010",6883 => "11100101",6884 => "11100001",6885 => "01011000",6886 => "11000111",6887 => "11101110",6888 => "11010110",6889 => "10111000",6890 => "00101100",6891 => "11101011",6892 => "10111011",6893 => "10010011",6894 => "01011110",6895 => "00110111",6896 => "11100111",6897 => "01100000",6898 => "10101111",6899 => "00011001",6900 => "01110110",6901 => "10001111",6902 => "11111110",6903 => "11100100",6904 => "10000001",6905 => "00110110",6906 => "01000110",6907 => "10101101",6908 => "00010101",6909 => "01011101",6910 => "00001000",6911 => "10100100",6912 => "10001001",6913 => "01011111",6914 => "01100010",6915 => "01111100",6916 => "00101100",6917 => "00010011",6918 => "10110110",6919 => "01011001",6920 => "11100001",6921 => "01010111",6922 => "01101110",6923 => "00111100",6924 => "10100110",6925 => "11101100",6926 => "00000111",6927 => "00001110",6928 => "10001000",6929 => "00011010",6930 => "11010000",6931 => "11001111",6932 => "11000101",6933 => "11010011",6934 => "01010101",6935 => "10011111",6936 => "01010100",6937 => "01111001",6938 => "01001010",6939 => "10010110",6940 => "10000001",6941 => "01110011",6942 => "11100000",6943 => "11010111",6944 => "10000101",6945 => "01000010",6946 => "11110111",6947 => "01000101",6948 => "01100000",6949 => "10101101",6950 => "00100101",6951 => "11001010",6952 => "11100110",6953 => "11100100",6954 => "11001101",6955 => "10111111",6956 => "01000111",6957 => "01100010",6958 => "00010110",6959 => "11100000",6960 => "11000110",6961 => "11010110",6962 => "00100011",6963 => "00001011",6964 => "00010110",6965 => "01100110",6966 => "10100101",6967 => "10111111",6968 => "11101001",6969 => "10001011",6970 => "00001011",6971 => "01110010",6972 => "01100000",6973 => "00110101",6974 => "01111111",6975 => "00111010",6976 => "11100100",6977 => "01011000",6978 => "11101111",6979 => "01011110",6980 => "01010000",6981 => "10100000",6982 => "10011111",6983 => "10001101",6984 => "11011101",6985 => "01100100",6986 => "01111100",6987 => "11001000",6988 => "10111001",6989 => "00001111",6990 => "00110110",6991 => "11011010",6992 => "01000010",6993 => "11001010",6994 => "11100101",6995 => "11011000",6996 => "10010111",6997 => "01000101",6998 => "00010001",6999 => "10010110",7000 => "00100101",7001 => "11101110",7002 => "00100100",7003 => "00011000",7004 => "01011111",7005 => "00011100",7006 => "10011101",7007 => "00101010",7008 => "11100100",7009 => "11010101",7010 => "10010010",7011 => "01100111",7012 => "11110010",7013 => "00100100",7014 => "01100010",7015 => "00011001",7016 => "00101110",7017 => "11100010",7018 => "01011000",7019 => "00001101",7020 => "01100111",7021 => "10111101",7022 => "11010000",7023 => "01000000",7024 => "01110110",7025 => "00101000",7026 => "01111000",7027 => "00001110",7028 => "10110011",7029 => "11010110",7030 => "00000001",7031 => "10110101",7032 => "10110011",7033 => "11101111",7034 => "11101010",7035 => "01111100",7036 => "11111110",7037 => "00101011",7038 => "00000101",7039 => "11111110",7040 => "00000001",7041 => "10001000",7042 => "00101110",7043 => "00010110",7044 => "01101010",7045 => "11101000",7046 => "10001111",7047 => "00110010",7048 => "10111110",7049 => "11000100",7050 => "11001001",7051 => "00111001",7052 => "11100011",7053 => "11010011",7054 => "01110011",7055 => "10010101",7056 => "01110011",7057 => "01011100",7058 => "10111001",7059 => "01011101",7060 => "00101110",7061 => "11000111",7062 => "11100011",7063 => "00100101",7064 => "01001100",7065 => "11101110",7066 => "01000100",7067 => "11000110",7068 => "00000010",7069 => "11110101",7070 => "11111001",7071 => "01110010",7072 => "00100010",7073 => "10000010",7074 => "11011111",7075 => "01000100",7076 => "10000011",7077 => "11011111",7078 => "10001111",7079 => "00010100",7080 => "00101011",7081 => "11000100",7082 => "01011011",7083 => "10001000",7084 => "00010100",7085 => "11000110",7086 => "00000101",7087 => "00100011",7088 => "10100000",7089 => "11011011",7090 => "11111010",7091 => "11111101",7092 => "11110100",7093 => "01000111",7094 => "11010010",7095 => "00101001",7096 => "10011110",7097 => "11011110",7098 => "10010001",7099 => "10110100",7100 => "00011110",7101 => "00101100",7102 => "01111100",7103 => "01111110",7104 => "01011100",7105 => "11110100",7106 => "01000001",7107 => "00110000",7108 => "01001101",7109 => "01110011",7110 => "01110001",7111 => "11111101",7112 => "01100110",7113 => "10000010",7114 => "10011100",7115 => "01100001",7116 => "00000110",7117 => "01100101",7118 => "10111001",7119 => "01111010",7120 => "01010000",7121 => "01011000",7122 => "00001110",7123 => "01110111",7124 => "00110111",7125 => "01110010",7126 => "00101000",7127 => "11100000",7128 => "11000111",7129 => "00111010",7130 => "00011110",7131 => "11010100",7132 => "10111101",7133 => "10001011",7134 => "01001100",7135 => "10001100",7136 => "01110011",7137 => "10110010",7138 => "10101010",7139 => "00000010",7140 => "11111100",7141 => "00001101",7142 => "01100101",7143 => "00111110",7144 => "11110110",7145 => "11110011",7146 => "11110110",7147 => "10010011",7148 => "01011011",7149 => "11101111",7150 => "01101011",7151 => "01010011",7152 => "00010011",7153 => "10011001",7154 => "11010111",7155 => "11101001",7156 => "11011111",7157 => "11110110",7158 => "10011100",7159 => "00000001",7160 => "00000001",7161 => "01010000",7162 => "00001101",7163 => "00010001",7164 => "10010110",7165 => "10101001",7166 => "01101011",7167 => "11000011",7168 => "00001001",7169 => "01000010",7170 => "11111010",7171 => "00100000",7172 => "10000110",7173 => "00000001",7174 => "00100110",7175 => "10001101",7176 => "00001100",7177 => "01011111",7178 => "11000001",7179 => "01000010",7180 => "01000001",7181 => "11010010",7182 => "00101100",7183 => "00000110",7184 => "00001111",7185 => "00101100",7186 => "11101000",7187 => "10001101",7188 => "01010111",7189 => "01010101",7190 => "01101010",7191 => "00001010",7192 => "00101010",7193 => "11111011",7194 => "10001100",7195 => "01001101",7196 => "10010001",7197 => "00001111",7198 => "01100000",7199 => "10110111",7200 => "00000111",7201 => "01100011",7202 => "10000011",7203 => "10101101",7204 => "10011101",7205 => "00011001",7206 => "11011101",7207 => "01100001",7208 => "10011011",7209 => "01111010",7210 => "10000100",7211 => "11000010",7212 => "00011110",7213 => "11010110",7214 => "00100010",7215 => "11011001",7216 => "01010101",7217 => "00101111",7218 => "10001001",7219 => "00101100",7220 => "00000000",7221 => "01010101",7222 => "11000111",7223 => "01101010",7224 => "01101000",7225 => "00100000",7226 => "11010100",7227 => "10110001",7228 => "11010101",7229 => "00100111",7230 => "01100011",7231 => "11010111",7232 => "00010101",7233 => "00011101",7234 => "00101110",7235 => "00101100",7236 => "01001110",7237 => "11000100",7238 => "01110011",7239 => "10010111",7240 => "01110011",7241 => "10000001",7242 => "10101000",7243 => "00010010",7244 => "10111101",7245 => "10010101",7246 => "10010001",7247 => "00110110",7248 => "01110000",7249 => "01100110",7250 => "01001111",7251 => "10010110",7252 => "01001010",7253 => "01010100",7254 => "01100000",7255 => "11111011",7256 => "00000001",7257 => "10000110",7258 => "11100100",7259 => "00111010",7260 => "10011100",7261 => "01101011",7262 => "01010001",7263 => "11100110",7264 => "01011110",7265 => "11100001",7266 => "01001011",7267 => "11101000",7268 => "10100011",7269 => "01110110",7270 => "10011111",7271 => "11101001",7272 => "11010110",7273 => "11100101",7274 => "10111001",7275 => "11101011",7276 => "01011001",7277 => "00111110",7278 => "11111100",7279 => "11100010",7280 => "10011000",7281 => "00001011",7282 => "10101100",7283 => "11101101",7284 => "11100010",7285 => "00101001",7286 => "11111111",7287 => "11011011",7288 => "01010000",7289 => "01011001",7290 => "11010010",7291 => "00100100",7292 => "10110001",7293 => "10110000",7294 => "11110010",7295 => "10111111",7296 => "00000010",7297 => "11110101",7298 => "00111011",7299 => "10111100",7300 => "11000010",7301 => "01100110",7302 => "10001101",7303 => "11111110",7304 => "10010111",7305 => "11100000",7306 => "01101110",7307 => "00111111",7308 => "11111001",7309 => "00000101",7310 => "10110000",7311 => "00001010",7312 => "01000101",7313 => "00100010",7314 => "00111001",7315 => "11000000",7316 => "01001101",7317 => "00011100",7318 => "00111101",7319 => "01010000",7320 => "11110001",7321 => "10001110",7322 => "01111001",7323 => "11010101",7324 => "10000010",7325 => "10111010",7326 => "00101001",7327 => "01001111",7328 => "00100000",7329 => "00111011",7330 => "00100111",7331 => "00111101",7332 => "11011001",7333 => "10100001",7334 => "01010000",7335 => "00100100",7336 => "01011001",7337 => "01000011",7338 => "01100000",7339 => "10100000",7340 => "11011111",7341 => "10001111",7342 => "01010000",7343 => "10000011",7344 => "11100001",7345 => "00001100",7346 => "00100010",7347 => "11111110",7348 => "11110100",7349 => "10011010",7350 => "00001001",7351 => "01011100",7352 => "00011010",7353 => "00100101",7354 => "10010100",7355 => "01101111",7356 => "00101111",7357 => "11101011",7358 => "01000111",7359 => "11000110",7360 => "10001110",7361 => "00001000",7362 => "10110011",7363 => "00111000",7364 => "00110110",7365 => "10001000",7366 => "10110111",7367 => "10110011",7368 => "00001111",7369 => "11011010",7370 => "01101010",7371 => "01111101",7372 => "10111001",7373 => "01110011",7374 => "01110010",7375 => "01011011",7376 => "00101000",7377 => "01010000",7378 => "01000000",7379 => "11000000",7380 => "10110110",7381 => "01000100",7382 => "10010100",7383 => "01100001",7384 => "11111101",7385 => "01100000",7386 => "10001111",7387 => "00101001",7388 => "11010010",7389 => "01111100",7390 => "01101111",7391 => "11111010",7392 => "01111011",7393 => "11001100",7394 => "00101100",7395 => "01011011",7396 => "11011011",7397 => "00101100",7398 => "01001111",7399 => "01001100",7400 => "00101111",7401 => "11011111",7402 => "01100111",7403 => "11101011",7404 => "00100010",7405 => "11000001",7406 => "00110000",7407 => "10011011",7408 => "00100101",7409 => "10101011",7410 => "11110010",7411 => "11100000",7412 => "01110101",7413 => "01010110",7414 => "10100101",7415 => "10010111",7416 => "11101000",7417 => "00110001",7418 => "01110000",7419 => "10111010",7420 => "10000100",7421 => "11000101",7422 => "11001010",7423 => "00110000",7424 => "10110111",7425 => "00111010",7426 => "00101100",7427 => "10010011",7428 => "01101111",7429 => "00000011",7430 => "11110111",7431 => "00110001",7432 => "00010010",7433 => "10001110",7434 => "10100000",7435 => "10101000",7436 => "00101010",7437 => "11000101",7438 => "00000011",7439 => "11000100",7440 => "01010111",7441 => "01101101",7442 => "10001111",7443 => "10100010",7444 => "01010101",7445 => "00101010",7446 => "00100111",7447 => "01100010",7448 => "01110100",7449 => "01010000",7450 => "01111001",7451 => "01011101",7452 => "00001010",7453 => "11100011",7454 => "01111001",7455 => "10100001",7456 => "01111110",7457 => "00001110",7458 => "10010110",7459 => "11011110",7460 => "01000110",7461 => "01000001",7462 => "01000111",7463 => "10010110",7464 => "01001101",7465 => "10101001",7466 => "11000000",7467 => "10010100",7468 => "10000010",7469 => "11011001",7470 => "11011110",7471 => "01010001",7472 => "01110111",7473 => "10100101",7474 => "10010111",7475 => "11001110",7476 => "01000010",7477 => "10010010",7478 => "10101101",7479 => "01011001",7480 => "01100111",7481 => "11110001",7482 => "11111000",7483 => "01111000",7484 => "01101111",7485 => "11001000",7486 => "00101100",7487 => "01000011",7488 => "01010101",7489 => "01110101",7490 => "01010011",7491 => "10110010",7492 => "10110101",7493 => "10010111",7494 => "11100110",7495 => "10011101",7496 => "10011010",7497 => "00101101",7498 => "11110001",7499 => "01000101",7500 => "11101011",7501 => "11111100",7502 => "11010110",7503 => "11111001",7504 => "11100011",7505 => "01000101",7506 => "00001000",7507 => "00110000",7508 => "01101000",7509 => "00111111",7510 => "01111100",7511 => "00001110",7512 => "11011000",7513 => "11111001",7514 => "00000001",7515 => "11001101",7516 => "00010001",7517 => "00001110",7518 => "01001101",7519 => "11010111",7520 => "01111100",7521 => "01001010",7522 => "11011100",7523 => "10010000",7524 => "11011010",7525 => "01000110",7526 => "11110100",7527 => "00101111",7528 => "00101000",7529 => "11000011",7530 => "00111100",7531 => "11010011",7532 => "01011101",7533 => "00010110",7534 => "10100000",7535 => "11100110",7536 => "00101010",7537 => "11011000",7538 => "00101100",7539 => "01001101",7540 => "10110110",7541 => "01011111",7542 => "01100111",7543 => "11001110",7544 => "11011000",7545 => "01110010",7546 => "10100111",7547 => "10001100",7548 => "01110101",7549 => "10111011",7550 => "11010000",7551 => "00110001",7552 => "01110111",7553 => "01001100",7554 => "11111011",7555 => "01010111",7556 => "10011000",7557 => "01000000",7558 => "00010001",7559 => "10111000",7560 => "00000001",7561 => "00111010",7562 => "01011111",7563 => "10001101",7564 => "01110100",7565 => "11111110",7566 => "11011101",7567 => "10010001",7568 => "11110110",7569 => "00000000",7570 => "10111001",7571 => "00011011",7572 => "00101011",7573 => "00010111",7574 => "10111111",7575 => "10000100",7576 => "11111001",7577 => "11100110",7578 => "11111000",7579 => "11110001",7580 => "00110000",7581 => "11010001",7582 => "10111110",7583 => "11001111",7584 => "00101001",7585 => "11010100",7586 => "11111001",7587 => "00011010",7588 => "01101000",7589 => "01000000",7590 => "11101100",7591 => "01010111",7592 => "00110110",7593 => "00000011",7594 => "10010000",7595 => "11111011",7596 => "11011111",7597 => "10110001",7598 => "01001000",7599 => "01110101",7600 => "10110111",7601 => "01110010",7602 => "01111001",7603 => "10011010",7604 => "01101011",7605 => "11111011",7606 => "11100110",7607 => "01110101",7608 => "00000011",7609 => "01101011",7610 => "01101110",7611 => "11100100",7612 => "11101010",7613 => "11101011",7614 => "01100110",7615 => "01010100",7616 => "00110000",7617 => "10010100",7618 => "10110000",7619 => "11100101",7620 => "00101011",7621 => "00110111",7622 => "10011011",7623 => "10000001",7624 => "01111101",7625 => "00000001",7626 => "11010110",7627 => "10110110",7628 => "10101111",7629 => "10110000",7630 => "00111111",7631 => "11000101",7632 => "10100011",7633 => "10010100",7634 => "01111010",7635 => "11111100",7636 => "10101101",7637 => "01101101",7638 => "10110010",7639 => "00010101",7640 => "11000011",7641 => "01110000",7642 => "11100110",7643 => "00101111",7644 => "10010000",7645 => "10001110",7646 => "00010000",7647 => "01001110",7648 => "01001111",7649 => "01011001",7650 => "01011011",7651 => "10010111",7652 => "11000001",7653 => "11010111",7654 => "01110011",7655 => "00000101",7656 => "11101111",7657 => "10111110",7658 => "00001000",7659 => "01001010",7660 => "01011101",7661 => "01100001",7662 => "00110001",7663 => "01100101",7664 => "11010010",7665 => "11111011",7666 => "00011000",7667 => "00100010",7668 => "11110011",7669 => "01100011",7670 => "00101110",7671 => "11101001",7672 => "00011000",7673 => "11001111",7674 => "10110110",7675 => "01100111",7676 => "10111110",7677 => "11000011",7678 => "10011111",7679 => "01111000",7680 => "11101111",7681 => "10000010",7682 => "01010000",7683 => "01111000",7684 => "10111101",7685 => "10100101",7686 => "01111000",7687 => "10001000",7688 => "00110110",7689 => "10100010",7690 => "01111000",7691 => "11100110",7692 => "10001001",7693 => "01010001",7694 => "10010100",7695 => "11111111",7696 => "00000111",7697 => "11011110",7698 => "10010100",7699 => "11111000",7700 => "11010100",7701 => "10001010",7702 => "00010010",7703 => "00001100",7704 => "01111111",7705 => "10001011",7706 => "01011100",7707 => "10010001",7708 => "01111101",7709 => "10101000",7710 => "01100000",7711 => "01100011",7712 => "11111001",7713 => "00101111",7714 => "00011001",7715 => "00101100",7716 => "00011101",7717 => "10010111",7718 => "10001001",7719 => "10101100",7720 => "11101010",7721 => "00010110",7722 => "00111011",7723 => "01011011",7724 => "11010010",7725 => "10001111",7726 => "10010010",7727 => "00011111",7728 => "00011101",7729 => "10010100",7730 => "11000111",7731 => "10010001",7732 => "00100011",7733 => "01100011",7734 => "01001100",7735 => "11101000",7736 => "10100011",7737 => "10010111",7738 => "11010000",7739 => "10010011",7740 => "01001110",7741 => "10011110",7742 => "10000011",7743 => "11101000",7744 => "11010011",7745 => "01011111",7746 => "10100100",7747 => "11000010",7748 => "00100011",7749 => "01010101",7750 => "11110001",7751 => "00100010",7752 => "01001100",7753 => "00101101",7754 => "00011100",7755 => "11111111",7756 => "11101111",7757 => "00010100",7758 => "01001011",7759 => "10000010",7760 => "11101101",7761 => "11000001",7762 => "01010101",7763 => "00011100",7764 => "01000010",7765 => "10101110",7766 => "00110001",7767 => "00010101",7768 => "11101110",7769 => "00011000",7770 => "10101101",7771 => "11010111",7772 => "10011101",7773 => "11100111",7774 => "11101101",7775 => "11001111",7776 => "00011101",7777 => "11010010",7778 => "11010110",7779 => "10010000",7780 => "00001101",7781 => "11011011",7782 => "00101011",7783 => "11101010",7784 => "10001100",7785 => "11000010",7786 => "00011111",7787 => "01001001",7788 => "00111100",7789 => "01101010",7790 => "00001100",7791 => "01001001",7792 => "11011001",7793 => "01111111",7794 => "10111011",7795 => "11100110",7796 => "10110011",7797 => "00111100",7798 => "01110001",7799 => "11111111",7800 => "01011110",7801 => "00100111",7802 => "00000111",7803 => "11001011",7804 => "10000011",7805 => "00111010",7806 => "01010011",7807 => "10001110",7808 => "00110110",7809 => "10110101",7810 => "00111110",7811 => "11110010",7812 => "10010010",7813 => "00100010",7814 => "01111011",7815 => "10011100",7816 => "01011001",7817 => "00110100",7818 => "00111100",7819 => "10000010",7820 => "11111111",7821 => "00000101",7822 => "10010010",7823 => "00001010",7824 => "10110101",7825 => "11010010",7826 => "10011000",7827 => "10000010",7828 => "00001110",7829 => "10001001",7830 => "11001100",7831 => "10111000",7832 => "01010100",7833 => "01110100",7834 => "11110001",7835 => "00000110",7836 => "01000100",7837 => "01001101",7838 => "01010110",7839 => "10001111",7840 => "01100001",7841 => "00000111",7842 => "01001100",7843 => "00100001",7844 => "01000010",7845 => "01101011",7846 => "01101101",7847 => "10000111",7848 => "01111011",7849 => "11110010",7850 => "01101111",7851 => "10101001",7852 => "11000101",7853 => "11100001",7854 => "00000111",7855 => "11111011",7856 => "10001110",7857 => "01000011",7858 => "00010100",7859 => "10001111",7860 => "11011000",7861 => "10001100",7862 => "10001101",7863 => "11111011",7864 => "11100110",7865 => "00010000",7866 => "01000100",7867 => "11100101",7868 => "01111111",7869 => "00000011",7870 => "11011111",7871 => "11111100",7872 => "01000100",7873 => "01001100",7874 => "01110011",7875 => "01000000",7876 => "01101100",7877 => "10110000",7878 => "00101001",7879 => "10110010",7880 => "01101101",7881 => "10111001",7882 => "11101110",7883 => "11000110",7884 => "10011110",7885 => "00010000",7886 => "10101110",7887 => "00011011",7888 => "01101000",7889 => "00001111",7890 => "11011000",7891 => "01101001",7892 => "11000100",7893 => "11011011",7894 => "10101100",7895 => "10111011",7896 => "01001110",7897 => "10001111",7898 => "00010001",7899 => "00010110",7900 => "00001010",7901 => "10110110",7902 => "01000011",7903 => "11100000",7904 => "10101001",7905 => "01000011",7906 => "00010001",7907 => "00101111",7908 => "01111101",7909 => "10111101",7910 => "01111000",7911 => "10000000",7912 => "10000010",7913 => "11011000",7914 => "00111110",7915 => "10100111",7916 => "00010000",7917 => "10001111",7918 => "11101010",7919 => "11110100",7920 => "00100010",7921 => "00111111",7922 => "01010110",7923 => "11011011",7924 => "10111001",7925 => "10101010",7926 => "01011100",7927 => "01101101",7928 => "10111110",7929 => "00110010",7930 => "11011100",7931 => "11111001",7932 => "11111000",7933 => "00111101",7934 => "01110110",7935 => "11101100",7936 => "11000011",7937 => "10011000",7938 => "00001010",7939 => "10001111",7940 => "01111011",7941 => "00101100",7942 => "00111001",7943 => "01000110",7944 => "11101100",7945 => "10101101",7946 => "00110111",7947 => "01000010",7948 => "10110010",7949 => "01011010",7950 => "10101001",7951 => "01111000",7952 => "01100100",7953 => "00011001",7954 => "10111000",7955 => "11001100",7956 => "11000001",7957 => "10110101",7958 => "01111111",7959 => "10001100",7960 => "10111001",7961 => "11011011",7962 => "00001001",7963 => "00110110",7964 => "11010100",7965 => "10101011",7966 => "00011101",7967 => "10011100",7968 => "11101110",7969 => "01001100",7970 => "01111011",7971 => "10000001",7972 => "11010111",7973 => "11010010",7974 => "00110010",7975 => "10011110",7976 => "10001011",7977 => "10000111",7978 => "01101011",7979 => "00101001",7980 => "01010000",7981 => "01001101",7982 => "00010111",7983 => "01000101",7984 => "10000001",7985 => "10100100",7986 => "00010100",7987 => "10101011",7988 => "00100010",7989 => "00111000",7990 => "10101001",7991 => "00101111",7992 => "10100110",7993 => "00001111",7994 => "01101111",7995 => "00110000",7996 => "01100011",7997 => "00101010",7998 => "11111100",7999 => "00110101",8000 => "00001111",8001 => "00111111",8002 => "01111011",8003 => "00001100",8004 => "10001110",8005 => "01111110",8006 => "01101001",8007 => "01111001",8008 => "10101001",8009 => "11100011",8010 => "00010101",8011 => "01001001",8012 => "01011000",8013 => "10101010",8014 => "01000101",8015 => "10111011",8016 => "10101110",8017 => "00110010",8018 => "10010001",8019 => "10001011",8020 => "00001000",8021 => "10111000",8022 => "10111010",8023 => "11011011",8024 => "10010101",8025 => "01101011",8026 => "01011010",8027 => "10111111",8028 => "00011011",8029 => "11111010",8030 => "11110111",8031 => "01011001",8032 => "00110010",8033 => "11101101",8034 => "00011100",8035 => "01101010",8036 => "00010011",8037 => "00011000",8038 => "01010100",8039 => "10100001",8040 => "00010110",8041 => "00011111",8042 => "10001011",8043 => "10001101",8044 => "11101101",8045 => "01111001",8046 => "01011010",8047 => "00001011",8048 => "11010111",8049 => "11011111",8050 => "10101110",8051 => "11001110",8052 => "00110000",8053 => "00101001",8054 => "01101000",8055 => "11000100",8056 => "00011001",8057 => "00010101",8058 => "00000101",8059 => "01010101",8060 => "11110010",8061 => "10110011",8062 => "11100100",8063 => "11110011",8064 => "01110001",8065 => "11010100",8066 => "11101100",8067 => "01000101",8068 => "01111110",8069 => "00101011",8070 => "00011001",8071 => "11110001",8072 => "10101101",8073 => "00010110",8074 => "00011011",8075 => "01101100",8076 => "00101011",8077 => "01000110",8078 => "01111100",8079 => "10011100",8080 => "00111011",8081 => "00001001",8082 => "01010100",8083 => "01100001",8084 => "00101001",8085 => "01001010",8086 => "00001001",8087 => "00011101",8088 => "11101000",8089 => "00110100",8090 => "00011001",8091 => "00000000",8092 => "11011110",8093 => "11111001",8094 => "10100101",8095 => "00011010",8096 => "10011010",8097 => "10011111",8098 => "00011010",8099 => "11111011",8100 => "00111101",8101 => "00001011",8102 => "11111001",8103 => "01010000",8104 => "00000110",8105 => "01111100",8106 => "11110001",8107 => "00010111",8108 => "01000100",8109 => "11110000",8110 => "11011101",8111 => "11111011",8112 => "01001001",8113 => "00000100",8114 => "11001101",8115 => "01101011",8116 => "10111110",8117 => "10110111",8118 => "00111101",8119 => "00111000",8120 => "00010011",8121 => "11110110",8122 => "10000101",8123 => "10110100",8124 => "11111001",8125 => "11110001",8126 => "00111001",8127 => "01101100",8128 => "01000010",8129 => "11101001",8130 => "00101001",8131 => "00000011",8132 => "00011010",8133 => "10111011",8134 => "01011110",8135 => "01111100",8136 => "00011000",8137 => "01011011",8138 => "10011110",8139 => "01100101",8140 => "00100100",8141 => "10101110",8142 => "01101001",8143 => "11000001",8144 => "01110011",8145 => "10111001",8146 => "10110110",8147 => "00111011",8148 => "00011110",8149 => "10000011",8150 => "11101001",8151 => "10000011",8152 => "01000011",8153 => "01001010",8154 => "00010000",8155 => "10010100",8156 => "01110100",8157 => "10001011",8158 => "01100011",8159 => "01001111",8160 => "01011110",8161 => "10000110",8162 => "00101000",8163 => "01101010",8164 => "10001100",8165 => "10001100",8166 => "11100000",8167 => "11001101",8168 => "11001100",8169 => "00111110",8170 => "00000011",8171 => "10101100",8172 => "10111110",8173 => "10010100",8174 => "00010010",8175 => "11100011",8176 => "11011011",8177 => "01011110",8178 => "00001100",8179 => "00010111",8180 => "00101111",8181 => "10101001",8182 => "01011001",8183 => "01011001",8184 => "00110100",8185 => "00000100",8186 => "10010111",8187 => "01000000",8188 => "01100011",8189 => "10011100",8190 => "00101100",8191 => "01000011",8192 => "10100101",8193 => "00000010",8194 => "10101001",8195 => "10100011",8196 => "00001101",8197 => "10100111",8198 => "10100100",8199 => "01111011",8200 => "10010100",8201 => "01010110",8202 => "11101000",8203 => "00010101",8204 => "01000110",8205 => "10101000",8206 => "11101110",8207 => "11100100",8208 => "01011110",8209 => "01100101",8210 => "10000001",8211 => "10111001",8212 => "00110101",8213 => "10001010",8214 => "10010011",8215 => "11001001",8216 => "11000011",8217 => "11110110",8218 => "10101101",8219 => "11001110",8220 => "10101001",8221 => "00011111",8222 => "10011000",8223 => "01000100",8224 => "00000001",8225 => "11111011",8226 => "01110100",8227 => "10010001",8228 => "00110000",8229 => "11000100",8230 => "10110011",8231 => "01101101",8232 => "10101101",8233 => "01010101",8234 => "00111110",8235 => "01010011",8236 => "11010011",8237 => "10000000",8238 => "11010111",8239 => "10001111",8240 => "10010001",8241 => "10011111",8242 => "00001111",8243 => "11110100",8244 => "11010000",8245 => "00101110",8246 => "00010110",8247 => "01011010",8248 => "01101110",8249 => "10101100",8250 => "11100011",8251 => "01011101",8252 => "10000110",8253 => "00010001",8254 => "00011000",8255 => "10100011",8256 => "01000010",8257 => "01011010",8258 => "11110111",8259 => "11111101",8260 => "01111101",8261 => "11000111",8262 => "10010100",8263 => "00100011",8264 => "01100011",8265 => "10101100",8266 => "11011100",8267 => "01100101",8268 => "01110101",8269 => "11111011",8270 => "00101010",8271 => "01001110",8272 => "10111000",8273 => "00101100",8274 => "10011110",8275 => "10101110",8276 => "10110000",8277 => "11111110",8278 => "11110100",8279 => "00010011",8280 => "10110001",8281 => "01001010",8282 => "11101000",8283 => "00100110",8284 => "11111111",8285 => "00011100",8286 => "00110101",8287 => "11011001",8288 => "00000011",8289 => "00110010",8290 => "00010001",8291 => "00100000",8292 => "01110111",8293 => "11001100",8294 => "01110001",8295 => "11100011",8296 => "11010101",8297 => "11001100",8298 => "00110101",8299 => "01000000",8300 => "11010001",8301 => "11100111",8302 => "01010111",8303 => "10010111",8304 => "11000011",8305 => "10100010",8306 => "10011010",8307 => "11001111",8308 => "00001111",8309 => "01101101",8310 => "01111110",8311 => "00100010",8312 => "00001010",8313 => "10011011",8314 => "10111001",8315 => "11101000",8316 => "10110100",8317 => "10001011",8318 => "00101001",8319 => "01110011",8320 => "00110100",8321 => "00101000",8322 => "00000110",8323 => "01001000",8324 => "01011110",8325 => "11011000",8326 => "11010001",8327 => "11001111",8328 => "11001010",8329 => "01000101",8330 => "11101110",8331 => "01110110",8332 => "11000111",8333 => "00000011",8334 => "11001100",8335 => "11111000",8336 => "11111101",8337 => "00100101",8338 => "01001101",8339 => "11011110",8340 => "10010111",8341 => "00001100",8342 => "11111011",8343 => "10000100",8344 => "11000110",8345 => "11111011",8346 => "01011001",8347 => "00110111",8348 => "10111010",8349 => "00010110",8350 => "00110110",8351 => "01110111",8352 => "01010101",8353 => "10101010",8354 => "11111111",8355 => "11110101",8356 => "00011000",8357 => "00001001",8358 => "11111100",8359 => "00010001",8360 => "01001010",8361 => "10000000",8362 => "11111010",8363 => "10000111",8364 => "01011100",8365 => "01000010",8366 => "01000000",8367 => "10001100",8368 => "10111000",8369 => "10011110",8370 => "00011101",8371 => "00101011",8372 => "11110010",8373 => "01001001",8374 => "00110000",8375 => "00001011",8376 => "11111011",8377 => "11010110",8378 => "11101100",8379 => "11110000",8380 => "01010100",8381 => "00101110",8382 => "11110000",8383 => "10100110",8384 => "00011101",8385 => "00110010",8386 => "11010000",8387 => "10000000",8388 => "01011111",8389 => "11101100",8390 => "01011000",8391 => "00110111",8392 => "10101001",8393 => "01000110",8394 => "11011011",8395 => "10100111",8396 => "11001101",8397 => "01010101",8398 => "00111111",8399 => "11010011",8400 => "10011111",8401 => "01111000",8402 => "10110000",8403 => "01111100",8404 => "11101010",8405 => "01110111",8406 => "00001001",8407 => "00001100",8408 => "00011011",8409 => "10111100",8410 => "00000001",8411 => "10110100",8412 => "10111000",8413 => "11100011",8414 => "00010100",8415 => "11000011",8416 => "00011011",8417 => "01001101",8418 => "11110001",8419 => "11101110",8420 => "00110111",8421 => "11101011",8422 => "00110110",8423 => "10101111",8424 => "10011011",8425 => "10001110",8426 => "01110011",8427 => "11111101",8428 => "10011010",8429 => "01111001",8430 => "11010000",8431 => "00111101",8432 => "10001011",8433 => "11111101",8434 => "11001011",8435 => "10111100",8436 => "00001101",8437 => "10110011",8438 => "01111000",8439 => "11001010",8440 => "11101010",8441 => "10110001",8442 => "11011110",8443 => "01100101",8444 => "00100101",8445 => "00000100",8446 => "01111101",8447 => "11011000",8448 => "10001010",8449 => "01110001",8450 => "01011010",8451 => "11000010",8452 => "01001010",8453 => "01101100",8454 => "10011100",8455 => "11110110",8456 => "01011100",8457 => "00000010",8458 => "01100011",8459 => "11110001",8460 => "00001000",8461 => "01101110",8462 => "01011011",8463 => "00111101",8464 => "10000001",8465 => "11001110",8466 => "11000000",8467 => "01111010",8468 => "01011101",8469 => "10010101",8470 => "00011001",8471 => "10110000",8472 => "10011101",8473 => "11111010",8474 => "01101110",8475 => "10001001",8476 => "11011011",8477 => "10001111",8478 => "11010000",8479 => "10001001",8480 => "00010110",8481 => "11000011",8482 => "00011001",8483 => "00011110",8484 => "00010011",8485 => "01001010",8486 => "01010000",8487 => "00100000",8488 => "01011010",8489 => "10101101",8490 => "11010011",8491 => "01100101",8492 => "10000101",8493 => "11010010",8494 => "10100011",8495 => "01110110",8496 => "00110000",8497 => "10011001",8498 => "10111010",8499 => "10010011",8500 => "00010000",8501 => "01011111",8502 => "01010110",8503 => "10111100",8504 => "10001110",8505 => "10110011",8506 => "01011110",8507 => "00111101",8508 => "11010110",8509 => "10011100",8510 => "00101001",8511 => "10011100",8512 => "11101001",8513 => "00011010",8514 => "11100011",8515 => "00110010",8516 => "01111000",8517 => "01111111",8518 => "00101101",8519 => "11011000",8520 => "10000011",8521 => "11111110",8522 => "10010110",8523 => "01000110",8524 => "00101001",8525 => "10010100",8526 => "01010111",8527 => "00101100",8528 => "01010001",8529 => "01010110",8530 => "01100011",8531 => "11001010",8532 => "00110000",8533 => "01101100",8534 => "01110000",8535 => "01111111",8536 => "01010001",8537 => "11101010",8538 => "10101001",8539 => "11101100",8540 => "11111000",8541 => "10110110",8542 => "00100111",8543 => "11101010",8544 => "10011010",8545 => "11010000",8546 => "11011010",8547 => "11101111",8548 => "11001111",8549 => "00001101",8550 => "11000000",8551 => "01111101",8552 => "00111001",8553 => "01000111",8554 => "01100110",8555 => "11111110",8556 => "10111010",8557 => "10011101",8558 => "01111000",8559 => "11111111",8560 => "01111111",8561 => "11101111",8562 => "01101110",8563 => "10101100",8564 => "00110111",8565 => "11111111",8566 => "00001000",8567 => "01001010",8568 => "11110110",8569 => "01100111",8570 => "01010010",8571 => "10001010",8572 => "11110111",8573 => "00001101",8574 => "01110110",8575 => "11011101",8576 => "01111011",8577 => "01010111",8578 => "00100001",8579 => "00111101",8580 => "11101111",8581 => "00011111",8582 => "11100100",8583 => "00011111",8584 => "00101001",8585 => "11110100",8586 => "00101000",8587 => "01100111",8588 => "00000000",8589 => "00101011",8590 => "11100100",8591 => "11110000",8592 => "00001001",8593 => "11111010",8594 => "10000010",8595 => "10001110",8596 => "00000111",8597 => "00000000",8598 => "11011100",8599 => "11111010",8600 => "10001110",8601 => "11101011",8602 => "01000000",8603 => "01100000",8604 => "00110011",8605 => "01010100",8606 => "10100011",8607 => "01011101",8608 => "10001010",8609 => "10101111",8610 => "11010000",8611 => "11100101",8612 => "10001110",8613 => "10011100",8614 => "00001101",8615 => "10101101",8616 => "11000111",8617 => "00101000",8618 => "01000101",8619 => "11110111",8620 => "11001100",8621 => "00101111",8622 => "01100111",8623 => "10100101",8624 => "01001101",8625 => "00001000",8626 => "10010011",8627 => "00001001",8628 => "00100011",8629 => "10100110",8630 => "00101111",8631 => "11110010",8632 => "10101000",8633 => "10110100",8634 => "10001010",8635 => "11000000",8636 => "00110100",8637 => "10101101",8638 => "01010011",8639 => "10000010",8640 => "10001001",8641 => "11100001",8642 => "00000101",8643 => "01000110",8644 => "01011011",8645 => "00100101",8646 => "11111010",8647 => "10101111",8648 => "01001001",8649 => "01011001",8650 => "11111010",8651 => "00011000",8652 => "01101110",8653 => "01011010",8654 => "10000111",8655 => "01011110",8656 => "00100111",8657 => "00000101",8658 => "01001110",8659 => "01010101",8660 => "00010111",8661 => "10110110",8662 => "10010010",8663 => "11100011",8664 => "01010100",8665 => "10100100",8666 => "01110100",8667 => "00110011",8668 => "01100111",8669 => "10111000",8670 => "01001011",8671 => "01000111",8672 => "10000011",8673 => "01100101",8674 => "10000010",8675 => "01110101",8676 => "01101111",8677 => "00110101",8678 => "11000111",8679 => "01100111",8680 => "01011011",8681 => "00000101",8682 => "01100100",8683 => "00100110",8684 => "11000100",8685 => "01000000",8686 => "01111001",8687 => "00101010",8688 => "10100011",8689 => "11000010",8690 => "00001110",8691 => "11101000",8692 => "11110101",8693 => "01101100",8694 => "00000101",8695 => "11000101",8696 => "11100001",8697 => "00101100",8698 => "10111100",8699 => "10001110",8700 => "01011001",8701 => "11001110",8702 => "11011000",8703 => "11000011",8704 => "10000111",8705 => "01001000",8706 => "00111110",8707 => "00101110",8708 => "01000111",8709 => "11001111",8710 => "10110011",8711 => "01011000",8712 => "11101111",8713 => "11101100",8714 => "11100000",8715 => "00000111",8716 => "00011101",8717 => "01110110",8718 => "11111000",8719 => "11101010",8720 => "00001011",8721 => "11001110",8722 => "01000010",8723 => "01100100",8724 => "01101001",8725 => "10000011",8726 => "11001100",8727 => "11001100",8728 => "10011000",8729 => "11110101",8730 => "10101110",8731 => "11000000",8732 => "01111100",8733 => "11000011",8734 => "10010101",8735 => "11011100",8736 => "11110010",8737 => "00010111",8738 => "11000100",8739 => "11000110",8740 => "10010101",8741 => "11001101",8742 => "01110110",8743 => "11001111",8744 => "01011111",8745 => "11101000",8746 => "10100111",8747 => "01110011",8748 => "01110001",8749 => "11000110",8750 => "01101110",8751 => "01101011",8752 => "11000001",8753 => "00110110",8754 => "01001111",8755 => "00110011",8756 => "11111010",8757 => "01000100",8758 => "00111100",8759 => "00111001",8760 => "10001000",8761 => "11100001",8762 => "01011100",8763 => "00011011",8764 => "11101010",8765 => "11001110",8766 => "00101110",8767 => "11100000",8768 => "00101110",8769 => "01000110",8770 => "10001000",8771 => "10110010",8772 => "01011100",8773 => "00100110",8774 => "01110110",8775 => "01101101",8776 => "00011100",8777 => "10110010",8778 => "01101001",8779 => "11100101",8780 => "10110101",8781 => "11101000",8782 => "01001000",8783 => "01000010",8784 => "00101000",8785 => "00011111",8786 => "11001000",8787 => "10010000",8788 => "00011000",8789 => "10100111",8790 => "00101010",8791 => "00001001",8792 => "01001110",8793 => "11010000",8794 => "10010110",8795 => "10010101",8796 => "10010111",8797 => "10000101",8798 => "11001101",8799 => "11001000",8800 => "10111010",8801 => "01010010",8802 => "01011000",8803 => "11000111",8804 => "10111100",8805 => "00001011",8806 => "01000000",8807 => "10100111",8808 => "11001111",8809 => "10101110",8810 => "11100001",8811 => "11110001",8812 => "11101001",8813 => "00101000",8814 => "00101000",8815 => "00001001",8816 => "00110110",8817 => "00010101",8818 => "10101110",8819 => "01001001",8820 => "10101100",8821 => "10010110",8822 => "01101111",8823 => "10001101",8824 => "10001110",8825 => "00010001",8826 => "01011101",8827 => "00100001",8828 => "00000111",8829 => "01001100",8830 => "01010001",8831 => "01001101",8832 => "11101110",8833 => "01010010",8834 => "01101110",8835 => "10101001",8836 => "00111010",8837 => "01011001",8838 => "00001001",8839 => "10100001",8840 => "11010111",8841 => "00110000",8842 => "10001001",8843 => "10010101",8844 => "01011101",8845 => "01010000",8846 => "11101010",8847 => "01100100",8848 => "10010011",8849 => "10000101",8850 => "11001000",8851 => "00000010",8852 => "01011100",8853 => "01000011",8854 => "01001101",8855 => "10110010",8856 => "00001010",8857 => "01010000",8858 => "01111010",8859 => "01110011",8860 => "00001111",8861 => "10111101",8862 => "01101100",8863 => "11100010",8864 => "01011000",8865 => "01011110",8866 => "11000101",8867 => "11001111",8868 => "10001000",8869 => "10110011",8870 => "00111110",8871 => "00001110",8872 => "01100010",8873 => "01001100",8874 => "00001100",8875 => "01111111",8876 => "11011010",8877 => "11111100",8878 => "01110100",8879 => "11101001",8880 => "10010001",8881 => "11000100",8882 => "11110110",8883 => "00111111",8884 => "01000000",8885 => "01001010",8886 => "11001000",8887 => "01010001",8888 => "11101101",8889 => "10011101",8890 => "10011000",8891 => "00000110",8892 => "10111001",8893 => "00010001",8894 => "11101110",8895 => "00001011",8896 => "11111011",8897 => "10011010",8898 => "00000110",8899 => "01111000",8900 => "01010000",8901 => "11110011",8902 => "10100101",8903 => "01101000",8904 => "00010111",8905 => "11110101",8906 => "00111010",8907 => "11000000",8908 => "01111100",8909 => "01111111",8910 => "10100001",8911 => "10101011",8912 => "01010000",8913 => "10100010",8914 => "01010100",8915 => "00011111",8916 => "10110000",8917 => "01010111",8918 => "00000100",8919 => "01010101",8920 => "10010101",8921 => "10000100",8922 => "01100110",8923 => "10001111",8924 => "01011101",8925 => "11111000",8926 => "00111111",8927 => "01111011",8928 => "01100101",8929 => "11101100",8930 => "00000000",8931 => "10111010",8932 => "10001001",8933 => "11101001",8934 => "00111010",8935 => "01001101",8936 => "11001100",8937 => "00110011",8938 => "00011000",8939 => "01100101",8940 => "01100110",8941 => "11000101",8942 => "10100000",8943 => "01011111",8944 => "01010100",8945 => "10000111",8946 => "00011110",8947 => "10100101",8948 => "00101000",8949 => "00111101",8950 => "01001001",8951 => "11101111",8952 => "00110110",8953 => "10101110",8954 => "01101001",8955 => "00001000",8956 => "00111000",8957 => "11100000",8958 => "11110110",8959 => "10010101",8960 => "10110110",8961 => "01110001",8962 => "00010001",8963 => "10111111",8964 => "11101110",8965 => "10010100",8966 => "11110101",8967 => "00001010",8968 => "11110000",8969 => "01010100",8970 => "01100101",8971 => "00011000",8972 => "00010100",8973 => "01011010",8974 => "10100001",8975 => "00110111",8976 => "01100000",8977 => "10100000",8978 => "11110010",8979 => "10110011",8980 => "00010001",8981 => "10001101",8982 => "11001000",8983 => "00110010",8984 => "01011110",8985 => "01010000",8986 => "01010101",8987 => "11110110",8988 => "01101000",8989 => "10011101",8990 => "01100111",8991 => "10111011",8992 => "11010100",8993 => "10100100",8994 => "10100000",8995 => "10011001",8996 => "11111111",8997 => "11110101",8998 => "10001100",8999 => "11010100",9000 => "00111000",9001 => "01111110",9002 => "10110010",9003 => "00000100",9004 => "11110101",9005 => "00100110",9006 => "11100011",9007 => "00101010",9008 => "00010010",9009 => "00100101",9010 => "10001110",9011 => "11111001",9012 => "01110100",9013 => "10100010",9014 => "11010011",9015 => "01001110",9016 => "00001001",9017 => "00011110",9018 => "10010010",9019 => "01101000",9020 => "01011101",9021 => "11111100",9022 => "01011101",9023 => "11101100",9024 => "10110010",9025 => "01111101",9026 => "11010100",9027 => "11111111",9028 => "01011011",9029 => "01110001",9030 => "01100101",9031 => "01001111",9032 => "01110010",9033 => "01101111",9034 => "00100001",9035 => "00111011",9036 => "11011101",9037 => "00000100",9038 => "00010001",9039 => "00011110",9040 => "11101001",9041 => "11010010",9042 => "00011000",9043 => "00101101",9044 => "11000000",9045 => "01101011",9046 => "10100111",9047 => "10010000",9048 => "10100101",9049 => "11111001",9050 => "11011001",9051 => "10101101",9052 => "10111111",9053 => "11011000",9054 => "11000001",9055 => "00110000",9056 => "01100101",9057 => "10110100",9058 => "01001000",9059 => "01011110",9060 => "11111100",9061 => "11111000",9062 => "11001110",9063 => "01101001",9064 => "10111100",9065 => "11011110",9066 => "11110001",9067 => "00011110",9068 => "11100010",9069 => "11101101",9070 => "01000111",9071 => "01111011",9072 => "01001001",9073 => "00000111",9074 => "10000110",9075 => "00001010",9076 => "00110100",9077 => "00000000",9078 => "10011011",9079 => "00110000",9080 => "10111001",9081 => "11000100",9082 => "00001100",9083 => "11110111",9084 => "00000101",9085 => "11000001",9086 => "10011110",9087 => "10011000",9088 => "01000111",9089 => "00011111",9090 => "01110110",9091 => "00000100",9092 => "11111101",9093 => "01101111",9094 => "10111001",9095 => "01010110",9096 => "01101000",9097 => "10001011",9098 => "10000101",9099 => "10111010",9100 => "01111001",9101 => "01011010",9102 => "00010001",9103 => "00011001",9104 => "10110111",9105 => "11110011",9106 => "11011100",9107 => "00010010",9108 => "01010101",9109 => "01110010",9110 => "00110001",9111 => "01001101",9112 => "10110010",9113 => "10111001",9114 => "00010010",9115 => "11000011",9116 => "11101001",9117 => "01100101",9118 => "01010001",9119 => "11011111",9120 => "01101011",9121 => "11111110",9122 => "11001001",9123 => "00000111",9124 => "10001011",9125 => "11000111",9126 => "01110110",9127 => "01111010",9128 => "10000111",9129 => "00011101",9130 => "01101001",9131 => "01000110",9132 => "00110001",9133 => "00001110",9134 => "01001001",9135 => "01000011",9136 => "10011111",9137 => "11001001",9138 => "10001001",9139 => "00010011",9140 => "10000101",9141 => "01100011",9142 => "11000000",9143 => "10101000",9144 => "10110101",9145 => "11100000",9146 => "11010000",9147 => "00010010",9148 => "10101111",9149 => "00110000",9150 => "00010110",9151 => "00101111",9152 => "11101001",9153 => "11011010",9154 => "00011011",9155 => "00101101",9156 => "00001100",9157 => "10110100",9158 => "11000110",9159 => "00101011",9160 => "01110001",9161 => "00011111",9162 => "10000001",9163 => "11010110",9164 => "00110101",9165 => "11000011",9166 => "11001110",9167 => "11011101",9168 => "11101110",9169 => "00100010",9170 => "10111001",9171 => "01001010",9172 => "10010000",9173 => "10010010",9174 => "11101011",9175 => "11100001",9176 => "00010100",9177 => "01000100",9178 => "10101111",9179 => "11111001",9180 => "00111001",9181 => "00101011",9182 => "10100000",9183 => "01101010",9184 => "10101011",9185 => "00001000",9186 => "11001111",9187 => "01011010",9188 => "01110011",9189 => "00111100",9190 => "11000110",9191 => "11111010",9192 => "11001100",9193 => "10101011",9194 => "11011100",9195 => "11110010",9196 => "01100010",9197 => "00001000",9198 => "01110000",9199 => "10111111",9200 => "01011001",9201 => "00101111",9202 => "10010001",9203 => "10011000",9204 => "11010100",9205 => "11110101",9206 => "11110001",9207 => "01101101",9208 => "01001001",9209 => "10010100",9210 => "01000000",9211 => "10011111",9212 => "01011100",9213 => "10010110",9214 => "10010101",9215 => "11011111",9216 => "10010100",9217 => "00010000",9218 => "11000111",9219 => "01111101",9220 => "01101011",9221 => "01011100",9222 => "11011100",9223 => "11011110",9224 => "10101001",9225 => "11101100",9226 => "11010100",9227 => "11111000",9228 => "11101010",9229 => "10001011",9230 => "00100000",9231 => "00100101",9232 => "10100010",9233 => "10011110",9234 => "11000100",9235 => "01111111",9236 => "11100010",9237 => "11110010",9238 => "10100101",9239 => "01101000",9240 => "10001000",9241 => "11010010",9242 => "10100001",9243 => "00110100",9244 => "10000100",9245 => "01101001",9246 => "00000100",9247 => "10110011",9248 => "01011101",9249 => "11000101",9250 => "11010101",9251 => "00010001",9252 => "00101011",9253 => "10001101",9254 => "11001010",9255 => "10010001",9256 => "10110100",9257 => "00001011",9258 => "00000101",9259 => "01011010",9260 => "00111011",9261 => "11010001",9262 => "01111110",9263 => "00110111",9264 => "01011110",9265 => "00110111",9266 => "01001001",9267 => "01100011",9268 => "10011101",9269 => "11001011",9270 => "01010110",9271 => "00011100",9272 => "01010100",9273 => "01000010",9274 => "00011001",9275 => "10101001",9276 => "00100110",9277 => "11100011",9278 => "01101101",9279 => "00010010",9280 => "00010111",9281 => "00010010",9282 => "10001011",9283 => "11110110",9284 => "00001010",9285 => "10111100",9286 => "10110111",9287 => "00111111",9288 => "00100001",9289 => "01110011",9290 => "11101011",9291 => "10100101",9292 => "00101110",9293 => "01110001",9294 => "10001000",9295 => "10111010",9296 => "10110111",9297 => "00100100",9298 => "01111011",9299 => "10000010",9300 => "00100000",9301 => "10000000",9302 => "01100001",9303 => "01010101",9304 => "00101010",9305 => "11101000",9306 => "11101001",9307 => "01110001",9308 => "11111101",9309 => "00001001",9310 => "00111101",9311 => "11001100",9312 => "00101000",9313 => "11010010",9314 => "11001101",9315 => "11110000",9316 => "01101101",9317 => "00011100",9318 => "00001011",9319 => "01001011",9320 => "11011110",9321 => "10001001",9322 => "10011011",9323 => "11101011",9324 => "01110111",9325 => "10001100",9326 => "00000010",9327 => "11100110",9328 => "01100100",9329 => "10010100",9330 => "10010001",9331 => "11101110",9332 => "00000010",9333 => "00100111",9334 => "11001001",9335 => "00011000",9336 => "00110100",9337 => "11001101",9338 => "00011101",9339 => "01011010",9340 => "00000001",9341 => "00100110",9342 => "00000110",9343 => "00000001",9344 => "01110011",9345 => "00010110",9346 => "00111001",9347 => "11001010",9348 => "11100000",9349 => "10101110",9350 => "01011101",9351 => "01110011",9352 => "11000110",9353 => "11111111",9354 => "00000011",9355 => "11100011",9356 => "00010011",9357 => "10011001",9358 => "10100001",9359 => "01101110",9360 => "01000101",9361 => "00001010",9362 => "00001110",9363 => "10010101",9364 => "00011001",9365 => "11001011",9366 => "10100111",9367 => "11111001",9368 => "10111111",9369 => "01000010",9370 => "00101000",9371 => "01110110",9372 => "11001000",9373 => "11101001",9374 => "11010100",9375 => "00110001",9376 => "10111101",9377 => "00101111",9378 => "10010001",9379 => "10000111",9380 => "00111110",9381 => "11001101",9382 => "01101010",9383 => "10011110",9384 => "11010110",9385 => "10011010",9386 => "11000000",9387 => "10101000",9388 => "10100111",9389 => "11010000",9390 => "11011001",9391 => "00111010",9392 => "10101110",9393 => "10001000",9394 => "01001011",9395 => "10000111",9396 => "11110111",9397 => "01100011",9398 => "10010110",9399 => "11000101",9400 => "10010100",9401 => "01100111",9402 => "00001010",9403 => "10000011",9404 => "00010001",9405 => "00110111",9406 => "11101110",9407 => "00101000",9408 => "00010111",9409 => "11000100",9410 => "10011110",9411 => "01100010",9412 => "00001110",9413 => "11010010",9414 => "10101011",9415 => "00101001",9416 => "10000011",9417 => "01110001",9418 => "11001001",9419 => "01111100",9420 => "01000111",9421 => "10011011",9422 => "01010000",9423 => "00011111",9424 => "10001110",9425 => "11110110",9426 => "11110111",9427 => "11000010",9428 => "01001000",9429 => "01100110",9430 => "01111011",9431 => "10101000",9432 => "11010111",9433 => "00111010",9434 => "01100111",9435 => "01100110",9436 => "10011100",9437 => "11101011",9438 => "10011011",9439 => "01010101",9440 => "10111111",9441 => "11000011",9442 => "01101101",9443 => "10100011",9444 => "11001001",9445 => "10110010",9446 => "11001100",9447 => "01111110",9448 => "11101001",9449 => "11101001",9450 => "10010100",9451 => "01010101",9452 => "11110100",9453 => "11101110",9454 => "01110110",9455 => "10011000",9456 => "10100010",9457 => "11011110",9458 => "00011110",9459 => "11110001",9460 => "11011101",9461 => "10110001",9462 => "11001000",9463 => "00100100",9464 => "11001001",9465 => "10100111",9466 => "01001000",9467 => "00110000",9468 => "00100100",9469 => "10101001",9470 => "00011000",9471 => "00010010",9472 => "01001001",9473 => "00011111",9474 => "01100100",9475 => "10011011",9476 => "11110100",9477 => "01000001",9478 => "10100000",9479 => "10001111",9480 => "00011000",9481 => "11101001",9482 => "10110000",9483 => "01000110",9484 => "11100111",9485 => "01111011",9486 => "11100100",9487 => "01010011",9488 => "00110010",9489 => "01010101",9490 => "10011110",9491 => "10000011",9492 => "11000100",9493 => "00011100",9494 => "10110000",9495 => "01101101",9496 => "01111000",9497 => "10000000",9498 => "10110101",9499 => "10100100",9500 => "10101001",9501 => "01101011",9502 => "11101100",9503 => "11100100",9504 => "01000111",9505 => "00011000",9506 => "01100011",9507 => "10011000",9508 => "00111110",9509 => "11100100",9510 => "00011111",9511 => "00110110",9512 => "11010001",9513 => "10101011",9514 => "00101110",9515 => "10001000",9516 => "01001110",9517 => "00010100",9518 => "11110100",9519 => "00101100",9520 => "10101100",9521 => "00010101",9522 => "11110010",9523 => "00101010",9524 => "10010111",9525 => "00011100",9526 => "00110010",9527 => "00011101",9528 => "11011010",9529 => "01111000",9530 => "00010001",9531 => "00100011",9532 => "01000011",9533 => "11100100",9534 => "01101011",9535 => "01111100",9536 => "01110101",9537 => "00111110",9538 => "10110010",9539 => "11101010",9540 => "11100000",9541 => "11001001",9542 => "01001100",9543 => "11100111",9544 => "11111011",9545 => "00011101",9546 => "10111010",9547 => "11001001",9548 => "01110010",9549 => "10010011",9550 => "10111110",9551 => "00001110",9552 => "10101000",9553 => "10011000",9554 => "00111111",9555 => "11101111",9556 => "11000001",9557 => "10111110",9558 => "00110101",9559 => "01000111",9560 => "10100101",9561 => "01001001",9562 => "01110000",9563 => "11001001",9564 => "01000111",9565 => "01000000",9566 => "10011011",9567 => "01010100",9568 => "10011100",9569 => "01100101",9570 => "01100000",9571 => "11101011",9572 => "10111011",9573 => "11000011",9574 => "10010111",9575 => "11000111",9576 => "11011101",9577 => "01101100",9578 => "01011100",9579 => "10101010",9580 => "00001110",9581 => "11100111",9582 => "11001000",9583 => "10110110",9584 => "11101110",9585 => "11111010",9586 => "01000100",9587 => "11111010",9588 => "11001100",9589 => "01011111",9590 => "00100100",9591 => "10010111",9592 => "11011010",9593 => "10101101",9594 => "00011010",9595 => "01010100",9596 => "00010100",9597 => "11101011",9598 => "01010011",9599 => "00101111",9600 => "10010010",9601 => "10101001",9602 => "10100111",9603 => "10011110",9604 => "01010001",9605 => "01101101",9606 => "11001011",9607 => "00100100",9608 => "11010010",9609 => "01110111",9610 => "00101000",9611 => "00001110",9612 => "01111111",9613 => "11100110",9614 => "00010010",9615 => "01110000",9616 => "01101100",9617 => "11001111",9618 => "11101000",9619 => "11011111",9620 => "01001000",9621 => "00011100",9622 => "10010000",9623 => "10111110",9624 => "00001000",9625 => "11011111",9626 => "01100010",9627 => "00110101",9628 => "11011111",9629 => "01001101",9630 => "01100111",9631 => "00101101",9632 => "00111110",9633 => "00010001",9634 => "11001110",9635 => "01000100",9636 => "01000111",9637 => "01101101",9638 => "10101000",9639 => "00100110",9640 => "00001100",9641 => "00010011",9642 => "00010010",9643 => "10011000",9644 => "01101101",9645 => "10000100",9646 => "11100001",9647 => "00101011",9648 => "11001111",9649 => "01111110",9650 => "00000100",9651 => "01100100",9652 => "01101010",9653 => "00110111",9654 => "01101110",9655 => "01000001",9656 => "10011101",9657 => "01001110",9658 => "11101110",9659 => "01101110",9660 => "10110001",9661 => "01100101",9662 => "10010111",9663 => "00101101",9664 => "00111100",9665 => "10001110",9666 => "01111101",9667 => "01011010",9668 => "10110100",9669 => "10100110",9670 => "11011000",9671 => "11111010",9672 => "01100101",9673 => "00001001",9674 => "01011001",9675 => "10000110",9676 => "00000001",9677 => "00101010",9678 => "00011100",9679 => "00101110",9680 => "01010000",9681 => "01101001",9682 => "11010010",9683 => "10101011",9684 => "10010001",9685 => "10010001",9686 => "00110110",9687 => "01110110",9688 => "01100000",9689 => "00111010",9690 => "11100001",9691 => "10111000",9692 => "00011110",9693 => "11111100",9694 => "10110101",9695 => "11101100",9696 => "10001001",9697 => "10000111",9698 => "01111110",9699 => "10000010",9700 => "01010111",9701 => "00000010",9702 => "10111111",9703 => "00101011",9704 => "00111100",9705 => "10111011",9706 => "11000001",9707 => "10000001",9708 => "01101101",9709 => "01110110",9710 => "10010111",9711 => "00000101",9712 => "11010101",9713 => "01011011",9714 => "10011000",9715 => "10111011",9716 => "11111111",9717 => "01100111",9718 => "00100110",9719 => "10110011",9720 => "01101100",9721 => "00010111",9722 => "10011100",9723 => "10001001",9724 => "01101000",9725 => "10010010",9726 => "01111110",9727 => "01110101",9728 => "01100100",9729 => "00011000",9730 => "11010100",9731 => "01000100",9732 => "00101111",9733 => "01000011",9734 => "11011001",9735 => "01010111",9736 => "11100001",9737 => "01101110",9738 => "00111001",9739 => "10100001",9740 => "01000000",9741 => "01000101",9742 => "10001101",9743 => "01111111",9744 => "10010010",9745 => "01101111",9746 => "11111101",9747 => "01001000",9748 => "10100001",9749 => "10111011",9750 => "11101101",9751 => "00010010",9752 => "10111010",9753 => "10000101",9754 => "01000111",9755 => "01010110",9756 => "10011100",9757 => "11100100",9758 => "00101111",9759 => "00000100",9760 => "01010100",9761 => "01100101",9762 => "01101111",9763 => "11000101",9764 => "11000110",9765 => "11001111",9766 => "00110000",9767 => "00111111",9768 => "01000110",9769 => "11110111",9770 => "00001001",9771 => "10101111",9772 => "11100001",9773 => "10100100",9774 => "00110010",9775 => "11010110",9776 => "10001010",9777 => "01011010",9778 => "11100110",9779 => "10010110",9780 => "01100111",9781 => "11001011",9782 => "01000100",9783 => "10101100",9784 => "11101100",9785 => "11111011",9786 => "10100001",9787 => "01110011",9788 => "10010010",9789 => "10111001",9790 => "01100011",9791 => "11100010",9792 => "11111100",9793 => "00110100",9794 => "01111001",9795 => "11010101",9796 => "01000001",9797 => "01111101",9798 => "10000111",9799 => "01011110",9800 => "00111011",9801 => "11110101",9802 => "00011100",9803 => "11100000",9804 => "00101101",9805 => "10001001",9806 => "01011101",9807 => "10101110",9808 => "01110001",9809 => "01110110",9810 => "10100111",9811 => "00001110",9812 => "01000111",9813 => "01100111",9814 => "00111110",9815 => "11111111",9816 => "10100100",9817 => "01110011",9818 => "10100001",9819 => "00001110",9820 => "01010101",9821 => "11110010",9822 => "10010010",9823 => "10000001",9824 => "00011100",9825 => "00110011",9826 => "11101110",9827 => "01011010",9828 => "01010111",9829 => "10011001",9830 => "11101101",9831 => "00001101",9832 => "00111010",9833 => "11000011",9834 => "10101001",9835 => "01000011",9836 => "00011011",9837 => "00111100",9838 => "11110010",9839 => "10001100",9840 => "10011000",9841 => "11111001",9842 => "11010010",9843 => "10110110",9844 => "00001101",9845 => "11111100",9846 => "01110101",9847 => "10101011",9848 => "00111110",9849 => "10001011",9850 => "01111011",9851 => "00011011",9852 => "01110000",9853 => "11101110",9854 => "00001000",9855 => "00000100",9856 => "11010011",9857 => "00100111",9858 => "11110101",9859 => "11010110",9860 => "01111000",9861 => "00001100",9862 => "01010001",9863 => "00100001",9864 => "01001101",9865 => "00110010",9866 => "01101010",9867 => "11100100",9868 => "10101111",9869 => "00001110",9870 => "00110100",9871 => "11101001",9872 => "00101010",9873 => "00011100",9874 => "11000101",9875 => "01110000",9876 => "11111110",9877 => "01110000",9878 => "01001110",9879 => "01001011",9880 => "01011110",9881 => "00011111",9882 => "10011010",9883 => "10001100",9884 => "01010000",9885 => "10000011",9886 => "11001111",9887 => "11111000",9888 => "10101010",9889 => "00010010",9890 => "01111100",9891 => "01101010",9892 => "10101011",9893 => "01110101",9894 => "01100001",9895 => "01000100",9896 => "00010101",9897 => "10011011",9898 => "11100000",9899 => "00001110",9900 => "00100001",9901 => "10100010",9902 => "00101111",9903 => "01011101",9904 => "10101010",9905 => "00101100",9906 => "11000001",9907 => "00000100",9908 => "00100101",9909 => "10110100",9910 => "00001101",9911 => "11101101",9912 => "10001111",9913 => "11101000",9914 => "00001101",9915 => "00110010",9916 => "00000110",9917 => "00011101",9918 => "01011011",9919 => "11101001",9920 => "00011100",9921 => "00000011",9922 => "11001111",9923 => "00011100",9924 => "00011111",9925 => "10010110",9926 => "10100101",9927 => "11010100",9928 => "10111110",9929 => "11001011",9930 => "00111011",9931 => "10011001",9932 => "10110110",9933 => "01010001",9934 => "11111101",9935 => "11010011",9936 => "01101111",9937 => "00101100",9938 => "10001110",9939 => "01000010",9940 => "01011101",9941 => "11110011",9942 => "11110010",9943 => "10101000",9944 => "10011000",9945 => "01101000",9946 => "11101011",9947 => "11000011",9948 => "01011001",9949 => "10111011",9950 => "11010110",9951 => "11110111",9952 => "01011011",9953 => "11110101",9954 => "11001101",9955 => "11101111",9956 => "00101110",9957 => "10011101",9958 => "11100111",9959 => "11100110",9960 => "00111100",9961 => "01110001",9962 => "00001101",9963 => "10010001",9964 => "10110000",9965 => "10111101",9966 => "00110000",9967 => "00011110",9968 => "00100111",9969 => "10001101",9970 => "10101111",9971 => "01110000",9972 => "10110110",9973 => "00011100",9974 => "01011111",9975 => "00100010",9976 => "00001110",9977 => "00111000",9978 => "10011000",9979 => "10001000",9980 => "01100111",9981 => "00111000",9982 => "10001011",9983 => "10100111",9984 => "10111001",9985 => "11101000",9986 => "10011110",9987 => "00100000",9988 => "10001110",9989 => "10010110",9990 => "11110111",9991 => "10011000",9992 => "10101110",9993 => "01011011",9994 => "01100001",9995 => "11101010",9996 => "10001000",9997 => "10001111",9998 => "10001011",9999 => "11011011",10000 => "00001100",10001 => "10000001",10002 => "11000100",10003 => "00000111",10004 => "00000111",10005 => "10111101",10006 => "00100001",10007 => "10100000",10008 => "00001100",10009 => "11000000",10010 => "11011010",10011 => "00010001",10012 => "10100100",10013 => "10101111",10014 => "10100010",10015 => "01101011",10016 => "01010100",10017 => "00011011",10018 => "10110111",10019 => "11010000",10020 => "11001011",10021 => "00001110",10022 => "10110100",10023 => "10000000",10024 => "00101010",10025 => "11011010",10026 => "00100110",10027 => "10011110",10028 => "11000011",10029 => "10110111",10030 => "00100101",10031 => "00000001",10032 => "00111100",10033 => "10011010",10034 => "10010101",10035 => "11010000",10036 => "00111001",10037 => "11100000",10038 => "11010111",10039 => "01110011",10040 => "00011111",10041 => "01011001",10042 => "00110011",10043 => "10111000",10044 => "01101000",10045 => "01100001",10046 => "00100101",10047 => "01110100",10048 => "00111010",10049 => "11111110",10050 => "01110000",10051 => "00110010",10052 => "10000111",10053 => "00111001",10054 => "01111000",10055 => "00110110",10056 => "01010100",10057 => "00001111",10058 => "10011110",10059 => "11011111",10060 => "01111001",10061 => "00010011",10062 => "10111000",10063 => "01001101",10064 => "11011011",10065 => "01010011",10066 => "01001101",10067 => "11011100",10068 => "01100000",10069 => "11001110",10070 => "10010010",10071 => "00101010",10072 => "00001100",10073 => "10110010",10074 => "00100001",10075 => "10010101",10076 => "00100000",10077 => "11110100",10078 => "00000101",10079 => "11011101",10080 => "01011011",10081 => "00101011",10082 => "00001111",10083 => "11011001",10084 => "10010011",10085 => "10001011",10086 => "01100011",10087 => "11001010",10088 => "10101001",10089 => "00000001",10090 => "11010001",10091 => "01011001",10092 => "00101011",10093 => "00111111",10094 => "11110111",10095 => "00000001",10096 => "01001101",10097 => "10111110",10098 => "10101101",10099 => "10111111",10100 => "11100000",10101 => "00111100",10102 => "00000111",10103 => "01010001",10104 => "10110110",10105 => "11011011",10106 => "00000111",10107 => "00010101",10108 => "00000010",10109 => "00001001",10110 => "10010011",10111 => "11001000",10112 => "01100010",10113 => "01111001",10114 => "01010101",10115 => "10001100",10116 => "10111001",10117 => "00011011",10118 => "10001011",10119 => "11111110",10120 => "11010010",10121 => "01011100",10122 => "01000111",10123 => "00011100",10124 => "10101111",10125 => "01101111",10126 => "01101111",10127 => "10101101",10128 => "01101010",10129 => "00000101",10130 => "11001101",10131 => "00001011",10132 => "11101010",10133 => "01110110",10134 => "01110001",10135 => "11111000",10136 => "10110010",10137 => "11110000",10138 => "11001110",10139 => "00000011",10140 => "11010010",10141 => "10010101",10142 => "11001011",10143 => "00111001",10144 => "11111001",10145 => "11110010",10146 => "10001100",10147 => "11011101",10148 => "10101110",10149 => "11010101",10150 => "00110011",10151 => "10001001",10152 => "10111000",10153 => "10110011",10154 => "10101011",10155 => "01010001",10156 => "10110110",10157 => "10010101",10158 => "10001001",10159 => "00000010",10160 => "00111001",10161 => "11110011",10162 => "00000100",10163 => "10001001",10164 => "00110000",10165 => "00100011",10166 => "11001100",10167 => "10100011",10168 => "01101001",10169 => "00010110",10170 => "11110010",10171 => "01111111",10172 => "10100010",10173 => "00100001",10174 => "10010111",10175 => "00001000",10176 => "11110010",10177 => "00011011",10178 => "11000001",10179 => "01010001",10180 => "01011111",10181 => "11011011",10182 => "11110011",10183 => "00111001",10184 => "00001110",10185 => "00000001",10186 => "01000001",10187 => "11000000",10188 => "00000010",10189 => "00000101",10190 => "01110001",10191 => "11101101",10192 => "11111101",10193 => "00010101",10194 => "01000111",10195 => "01010010",10196 => "10011000",10197 => "00110100",10198 => "11100100",10199 => "00100010",10200 => "00101001",10201 => "11101011",10202 => "01101100",10203 => "11000010",10204 => "10011001",10205 => "11110011",10206 => "01010110",10207 => "00111000",10208 => "10010011",10209 => "01110100",10210 => "01000110",10211 => "10001111",10212 => "11110001",10213 => "10101110",10214 => "11001011",10215 => "00111101",10216 => "01110100",10217 => "10110010",10218 => "01101101",10219 => "01100001",10220 => "11001001",10221 => "00110010",10222 => "11011110",10223 => "01000000",10224 => "10110100",10225 => "00000001",10226 => "10111101",10227 => "11110110",10228 => "01111001",10229 => "11111100",10230 => "11011111",10231 => "10110110",10232 => "00101101",10233 => "01011011",10234 => "01001111",10235 => "10100111",10236 => "00010100",10237 => "11010011",10238 => "10100011",10239 => "10000001",10240 => "11010001",10241 => "01111111",10242 => "11101011",10243 => "10111010",10244 => "11010111",10245 => "01100001",10246 => "10110100",10247 => "10101110",10248 => "01010001",10249 => "10101101",10250 => "01111101",10251 => "00000100",10252 => "10010010",10253 => "00000001",10254 => "11001100",10255 => "11011000",10256 => "01110011",10257 => "01000010",10258 => "11101011",10259 => "00100000",10260 => "11101111",10261 => "00110001",10262 => "10000010",10263 => "01001110",10264 => "10111110",10265 => "00100010",10266 => "01011101",10267 => "01100110",10268 => "00000110",10269 => "11110000",10270 => "01000100",10271 => "11101010",10272 => "01011101",10273 => "01111101",10274 => "10110101",10275 => "01101111",10276 => "01001001",10277 => "00000001",10278 => "11000100",10279 => "00101011",10280 => "00000011",10281 => "00010000",10282 => "10001011",10283 => "01111111",10284 => "00001100",10285 => "01111001",10286 => "11001010",10287 => "11100101",10288 => "00011001",10289 => "00001110",10290 => "11000010",10291 => "11100000",10292 => "11000110",10293 => "10111000",10294 => "00011001",10295 => "11001100",10296 => "10110001",10297 => "01111000",10298 => "00011100",10299 => "10011111",10300 => "10000110",10301 => "00001110",10302 => "01101010",10303 => "01000100",10304 => "11011001",10305 => "10110010",10306 => "10011110",10307 => "01010101",10308 => "11111001",10309 => "00111010",10310 => "11110111",10311 => "01000111",10312 => "11110111",10313 => "10111101",10314 => "11000111",10315 => "00001011",10316 => "01101010",10317 => "10010110",10318 => "11011110",10319 => "01000111",10320 => "00000001",10321 => "00110000",10322 => "10100100",10323 => "10110110",10324 => "01100110",10325 => "00000000",10326 => "10010101",10327 => "10100101",10328 => "01000111",10329 => "00110001",10330 => "10010010",10331 => "11100111",10332 => "00110001",10333 => "00111101",10334 => "01111011",10335 => "10011011",10336 => "00101011",10337 => "00101001",10338 => "00010011",10339 => "01000111",10340 => "01011000",10341 => "01110010",10342 => "11000100",10343 => "11000111",10344 => "11110111",10345 => "01011101",10346 => "01011001",10347 => "11001101",10348 => "01111101",10349 => "10100011",10350 => "10110110",10351 => "00011101",10352 => "01010100",10353 => "11100000",10354 => "01001110",10355 => "01000010",10356 => "10000101",10357 => "00001100",10358 => "10110001",10359 => "01101010",10360 => "10110111",10361 => "10001101",10362 => "11100110",10363 => "11100100",10364 => "00010010",10365 => "00110110",10366 => "00011100",10367 => "01100001",10368 => "01000001",10369 => "01110011",10370 => "10101001",10371 => "11011000",10372 => "00011101",10373 => "00000100",10374 => "10010000",10375 => "11100010",10376 => "01101100",10377 => "10101101",10378 => "10010101",10379 => "10011110",10380 => "10000111",10381 => "01010001",10382 => "00011111",10383 => "01011101",10384 => "01111111",10385 => "11111011",10386 => "10101010",10387 => "01001110",10388 => "10100010",10389 => "10111010",10390 => "10111001",10391 => "10011111",10392 => "11111100",10393 => "01110110",10394 => "10011111",10395 => "01111000",10396 => "11100101",10397 => "10110100",10398 => "00000101",10399 => "11101011",10400 => "11011011",10401 => "01010000",10402 => "01110100",10403 => "10011000",10404 => "00110111",10405 => "11011010",10406 => "00000001",10407 => "11000000",10408 => "00110100",10409 => "11111100",10410 => "11011101",10411 => "01110110",10412 => "00111001",10413 => "11101000",10414 => "01111001",10415 => "10001010",10416 => "00001010",10417 => "00010101",10418 => "01011011",10419 => "10001001",10420 => "01011010",10421 => "00110011",10422 => "00000110",10423 => "00100110",10424 => "10101100",10425 => "11111011",10426 => "10111001",10427 => "01111001",10428 => "11000011",10429 => "01001111",10430 => "00000001",10431 => "10100010",10432 => "11111000",10433 => "10100010",10434 => "01011101",10435 => "10110110",10436 => "10011000",10437 => "00010100",10438 => "10110010",10439 => "01111110",10440 => "01011100",10441 => "01110111",10442 => "01011001",10443 => "00101011",10444 => "00101100",10445 => "10011110",10446 => "10010100",10447 => "00100110",10448 => "01000000",10449 => "11010011",10450 => "00110011",10451 => "11001001",10452 => "11000111",10453 => "00010001",10454 => "11111000",10455 => "11101110",10456 => "10010010",10457 => "00101111",10458 => "01101000",10459 => "01101111",10460 => "11000001",10461 => "00000011",10462 => "11101100",10463 => "01010000",10464 => "10111100",10465 => "10111100",10466 => "00010100",10467 => "00100111",10468 => "01100101",10469 => "10100010",10470 => "00110001",10471 => "10110000",10472 => "01011101",10473 => "10011110",10474 => "00011000",10475 => "11110001",10476 => "10011101",10477 => "11101011",10478 => "11110100",10479 => "01101010",10480 => "10011101",10481 => "10000111",10482 => "11011001",10483 => "10011001",10484 => "10010111",10485 => "10010010",10486 => "01101110",10487 => "01101010",10488 => "01000010",10489 => "00010011",10490 => "01100001",10491 => "10100010",10492 => "01110000",10493 => "01100001",10494 => "00001100",10495 => "10111001",10496 => "10111010",10497 => "00000011",10498 => "01000101",10499 => "10111111",10500 => "00011111",10501 => "00011101",10502 => "01001100",10503 => "10110100",10504 => "00010010",10505 => "01010011",10506 => "11101011",10507 => "11001010",10508 => "10010100",10509 => "01000110",10510 => "11100101",10511 => "01110111",10512 => "11000011",10513 => "10111111",10514 => "00010001",10515 => "00001110",10516 => "10001111",10517 => "00000001",10518 => "00101011",10519 => "11001110",10520 => "00010110",10521 => "10000011",10522 => "01000100",10523 => "11001001",10524 => "11111110",10525 => "01000010",10526 => "11111011",10527 => "00111000",10528 => "11100100",10529 => "01001101",10530 => "01001001",10531 => "10111111",10532 => "11001010",10533 => "00001111",10534 => "10111110",10535 => "01100100",10536 => "01111110",10537 => "01010001",10538 => "11001010",10539 => "11100101",10540 => "00100010",10541 => "10100000",10542 => "11110111",10543 => "00100111",10544 => "11011100",10545 => "01011101",10546 => "01010110",10547 => "10100100",10548 => "00111000",10549 => "11000101",10550 => "00010001",10551 => "11001111",10552 => "10001110",10553 => "10110111",10554 => "01101010",10555 => "10110111",10556 => "01100110",10557 => "10010000",10558 => "01011011",10559 => "00000010",10560 => "11001000",10561 => "00111010",10562 => "00100001",10563 => "00010100",10564 => "00101110",10565 => "01001011",10566 => "01001001",10567 => "01001110",10568 => "00100010",10569 => "01010000",10570 => "00001011",10571 => "00101101",10572 => "10111000",10573 => "01010101",10574 => "10001111",10575 => "00111110",10576 => "10010100",10577 => "01001011",10578 => "10110100",10579 => "01100111",10580 => "00011101",10581 => "01010001",10582 => "11011001",10583 => "11011101",10584 => "11000110",10585 => "11100000",10586 => "01011011",10587 => "01110100",10588 => "01110010",10589 => "11011001",10590 => "01001111",10591 => "10100001",10592 => "10110000",10593 => "11001110",10594 => "10010011",10595 => "00111110",10596 => "10000011",10597 => "10000000",10598 => "11001110",10599 => "01111000",10600 => "11000010",10601 => "01111111",10602 => "11001000",10603 => "11011001",10604 => "11110011",10605 => "01100100",10606 => "01011000",10607 => "10000000",10608 => "00010111",10609 => "01111100",10610 => "10001000",10611 => "11010000",10612 => "00111010",10613 => "10100101",10614 => "00001010",10615 => "00100101",10616 => "01110001",10617 => "00001101",10618 => "11011010",10619 => "11111000",10620 => "11001000",10621 => "01011111",10622 => "11111000",10623 => "01111110",10624 => "10101100",10625 => "10101111",10626 => "10100000",10627 => "00101000",10628 => "00101111",10629 => "01000001",10630 => "01110000",10631 => "00001010",10632 => "00101101",10633 => "11101011",10634 => "11010111",10635 => "11101010",10636 => "10011100",10637 => "01111110",10638 => "01010011",10639 => "01000111",10640 => "01101010",10641 => "00110001",10642 => "10100110",10643 => "11011011",10644 => "00001111",10645 => "10011100",10646 => "00011010",10647 => "00000001",10648 => "10101010",10649 => "00000001",10650 => "00010010",10651 => "11110001",10652 => "00010010",10653 => "00000101",10654 => "11011000",10655 => "11000111",10656 => "10000110",10657 => "11110101",10658 => "00000001",10659 => "10100100",10660 => "00111110",10661 => "10101010",10662 => "11101000",10663 => "00101101",10664 => "01000111",10665 => "10001100",10666 => "11111011",10667 => "11000100",10668 => "11010111",10669 => "01111010",10670 => "10001001",10671 => "10110000",10672 => "01011001",10673 => "01000110",10674 => "01100011",10675 => "01111110",10676 => "10110010",10677 => "11000110",10678 => "11101010",10679 => "01110000",10680 => "00000011",10681 => "01100100",10682 => "01111111",10683 => "11000011",10684 => "01000111",10685 => "10101100",10686 => "10100000",10687 => "00111010",10688 => "11110011",10689 => "01100000",10690 => "01000001",10691 => "11101100",10692 => "00011111",10693 => "01111100",10694 => "10101011",10695 => "01100011",10696 => "10111001",10697 => "11111100",10698 => "01011000",10699 => "10100110",10700 => "01101111",10701 => "11110010",10702 => "10001010",10703 => "00110001",10704 => "11000011",10705 => "00110010",10706 => "11101100",10707 => "10100001",10708 => "11011101",10709 => "10000001",10710 => "00110001",10711 => "00001010",10712 => "11101001",10713 => "00111110",10714 => "10111100",10715 => "01011100",10716 => "10111011",10717 => "01010110",10718 => "00010001",10719 => "00000000",10720 => "01111100",10721 => "10001000",10722 => "01010111",10723 => "10100001",10724 => "11000000",10725 => "11111000",10726 => "01011101",10727 => "10100100",10728 => "00010100",10729 => "00100001",10730 => "01010000",10731 => "10001001",10732 => "11101100",10733 => "00010100",10734 => "11011010",10735 => "10110101",10736 => "00001110",10737 => "10001101",10738 => "00100011",10739 => "00100110",10740 => "01010010",10741 => "11111000",10742 => "10101010",10743 => "11001110",10744 => "01000111",10745 => "11001010",10746 => "00110100",10747 => "11010010",10748 => "10010101",10749 => "01111000",10750 => "10100011",10751 => "00100000",10752 => "01001110",10753 => "10000000",10754 => "10101111",10755 => "11111011",10756 => "10110000",10757 => "00100000",10758 => "00001000",10759 => "10000000",10760 => "10110101",10761 => "10110001",10762 => "11110011",10763 => "00111100",10764 => "11001000",10765 => "11101101",10766 => "11110011",10767 => "01110111",10768 => "01100011",10769 => "11000100",10770 => "10101100",10771 => "01010000",10772 => "01111110",10773 => "01101011",10774 => "00010010",10775 => "11011110",10776 => "01111100",10777 => "10011001",10778 => "11101110",10779 => "00001101",10780 => "01100101",10781 => "01010101",10782 => "11010000",10783 => "11000111",10784 => "01000000",10785 => "01110101",10786 => "01110111",10787 => "11000011",10788 => "10010101",10789 => "10110111",10790 => "11101111",10791 => "10100101",10792 => "10111100",10793 => "10100010",10794 => "01110011",10795 => "11011001",10796 => "01111100",10797 => "01111001",10798 => "10010001",10799 => "00110100",10800 => "10001001",10801 => "00010100",10802 => "10111011",10803 => "01100010",10804 => "10111011",10805 => "11111010",10806 => "01011010",10807 => "11111010",10808 => "01100111",10809 => "10000101",10810 => "00010100",10811 => "10101000",10812 => "00000101",10813 => "00110010",10814 => "10101111",10815 => "10100110",10816 => "11011010",10817 => "01011000",10818 => "00001001",10819 => "11101100",10820 => "11100111",10821 => "00101011",10822 => "10110101",10823 => "10110000",10824 => "01011100",10825 => "00100000",10826 => "00010111",10827 => "11100110",10828 => "11101011",10829 => "01101111",10830 => "11100111",10831 => "01010111",10832 => "01010011",10833 => "00101111",10834 => "10110110",10835 => "01100111",10836 => "01001001",10837 => "11001000",10838 => "00101101",10839 => "11011011",10840 => "10111110",10841 => "01010100",10842 => "00110111",10843 => "00000010",10844 => "01101000",10845 => "10000010",10846 => "00100010",10847 => "00010011",10848 => "10001101",10849 => "10010010",10850 => "11101011",10851 => "10011000",10852 => "11000010",10853 => "01110100",10854 => "00001100",10855 => "10100100",10856 => "10010000",10857 => "10100111",10858 => "10001011",10859 => "01110010",10860 => "01001101",10861 => "00011001",10862 => "11100011",10863 => "00010011",10864 => "10111101",10865 => "00110100",10866 => "01011110",10867 => "10100101",10868 => "00000011",10869 => "00001001",10870 => "11011001",10871 => "01101101",10872 => "00001010",10873 => "00110111",10874 => "00110110",10875 => "10101011",10876 => "01111000",10877 => "10000010",10878 => "01100011",10879 => "11110010",10880 => "01000110",10881 => "01000111",10882 => "10000010",10883 => "11111101",10884 => "00100010",10885 => "11111110",10886 => "10100000",10887 => "01011011",10888 => "00100101",10889 => "01011110",10890 => "10000110",10891 => "01101010",10892 => "01100010",10893 => "11000101",10894 => "10111000",10895 => "10011101",10896 => "10110001",10897 => "10001110",10898 => "11111001",10899 => "11101001",10900 => "10111101",10901 => "00101011",10902 => "01100111",10903 => "01001100",10904 => "01010101",10905 => "00101000",10906 => "00100011",10907 => "01101101",10908 => "00111000",10909 => "10010100",10910 => "00101100",10911 => "00110110",10912 => "01010010",10913 => "00010011",10914 => "00101000",10915 => "00010001",10916 => "00111100",10917 => "00011110",10918 => "10110100",10919 => "11000011",10920 => "00100111",10921 => "01011110",10922 => "00000101",10923 => "10111011",10924 => "01101010",10925 => "00110000",10926 => "11001010",10927 => "10011100",10928 => "00010000",10929 => "00011011",10930 => "01110110",10931 => "10001101",10932 => "00110110",10933 => "10100111",10934 => "11101111",10935 => "00000000",10936 => "10011010",10937 => "01010011",10938 => "10100100",10939 => "00010101",10940 => "01110001",10941 => "11000101",10942 => "11000100",10943 => "01010001",10944 => "10100001",10945 => "00001011",10946 => "11101110",10947 => "10001000",10948 => "01110111",10949 => "10011100",10950 => "01111000",10951 => "01001000",10952 => "01111101",10953 => "00001010",10954 => "00001001",10955 => "00100011",10956 => "11110010",10957 => "11011001",10958 => "10011100",10959 => "00110110",10960 => "01001010",10961 => "00011001",10962 => "11110111",10963 => "00100100",10964 => "00001110",10965 => "00110011",10966 => "11110001",10967 => "00110010",10968 => "01001111",10969 => "10000111",10970 => "00000110",10971 => "00110010",10972 => "10000111",10973 => "11110110",10974 => "11100110",10975 => "11011110",10976 => "01101111",10977 => "10110010",10978 => "00100000",10979 => "00000010",10980 => "01111110",10981 => "00100010",10982 => "00100010",10983 => "11110000",10984 => "00101101",10985 => "10100101",10986 => "11111001",10987 => "00110111",10988 => "10011101",10989 => "11011110",10990 => "11001101",10991 => "10100010",10992 => "10001001",10993 => "11011100",10994 => "10101010",10995 => "00011011",10996 => "01011001",10997 => "10110011",10998 => "00011101",10999 => "10011100",11000 => "11110110",11001 => "11010000",11002 => "11111010",11003 => "00111111",11004 => "10101010",11005 => "10010111",11006 => "10110010",11007 => "10011110",11008 => "11110000",11009 => "11101001",11010 => "10011010",11011 => "10110010",11012 => "01011001",11013 => "11010000",11014 => "11010110",11015 => "11101011",11016 => "10110011",11017 => "00001100",11018 => "00101100",11019 => "00111100",11020 => "00111000",11021 => "00001111",11022 => "00000000",11023 => "01100100",11024 => "11110101",11025 => "00101000",11026 => "00000011",11027 => "01010101",11028 => "11010001",11029 => "01101101",11030 => "11011101",11031 => "01110111",11032 => "00111000",11033 => "10010001",11034 => "01101101",11035 => "01111011",11036 => "10001110",11037 => "01000111",11038 => "01010101",11039 => "00110011",11040 => "00000010",11041 => "11100000",11042 => "01011100",11043 => "11100100",11044 => "01011011",11045 => "00100010",11046 => "01000001",11047 => "11110101",11048 => "10001010",11049 => "00111000",11050 => "11110111",11051 => "01000100",11052 => "10001110",11053 => "00010110",11054 => "00100110",11055 => "01000001",11056 => "00111110",11057 => "10011000",11058 => "10010111",11059 => "01010011",11060 => "10110110",11061 => "10111110",11062 => "11110100",11063 => "01100010",11064 => "11010001",11065 => "01001101",11066 => "10010010",11067 => "01100000",11068 => "00010111",11069 => "11100011",11070 => "11010101",11071 => "01100000",11072 => "11011011",11073 => "10000111",11074 => "10000100",11075 => "11100000",11076 => "11011010",11077 => "11001100",11078 => "00010111",11079 => "10110001",11080 => "11001110",11081 => "10110011",11082 => "00000100",11083 => "10101100",11084 => "00111011",11085 => "01111001",11086 => "00000100",11087 => "01000001",11088 => "01101010",11089 => "01111100",11090 => "11101011",11091 => "00111001",11092 => "00111101",11093 => "01110000",11094 => "01111011",11095 => "00101010",11096 => "10101111",11097 => "10011000",11098 => "01010110",11099 => "11100101",11100 => "11010001",11101 => "10001011",11102 => "11000100",11103 => "10111001",11104 => "00100110",11105 => "01010101",11106 => "10011001",11107 => "11101111",11108 => "00101010",11109 => "10010001",11110 => "11011001",11111 => "11000110",11112 => "00011111",11113 => "10100001",11114 => "10100011",11115 => "01001111",11116 => "11010000",11117 => "00011001",11118 => "01010101",11119 => "01001000",11120 => "10100101",11121 => "00110001",11122 => "11111000",11123 => "10100100",11124 => "01110001",11125 => "11010011",11126 => "01010011",11127 => "01100000",11128 => "00100000",11129 => "10111001",11130 => "10000010",11131 => "00000001",11132 => "00011011",11133 => "10110001",11134 => "01011111",11135 => "00000111",11136 => "00100111",11137 => "10101110",11138 => "01011101",11139 => "01001101",11140 => "11101011",11141 => "10011101",11142 => "11010001",11143 => "11010111",11144 => "10011111",11145 => "00001010",11146 => "01011101",11147 => "10001010",11148 => "00110001",11149 => "11011000",11150 => "10000000",11151 => "11110101",11152 => "01101000",11153 => "01111101",11154 => "00001000",11155 => "11000101",11156 => "00111100",11157 => "10000001",11158 => "10100101",11159 => "01111010",11160 => "01110010",11161 => "00011010",11162 => "01000010",11163 => "11101101",11164 => "01110100",11165 => "00000011",11166 => "01101101",11167 => "01011000",11168 => "01111101",11169 => "00111101",11170 => "10101010",11171 => "00100010",11172 => "01110011",11173 => "10000000",11174 => "10110110",11175 => "01000011",11176 => "11100101",11177 => "10101111",11178 => "10110100",11179 => "01000100",11180 => "10101111",11181 => "00101101",11182 => "01101011",11183 => "01001001",11184 => "01010101",11185 => "10111000",11186 => "01000000",11187 => "00111100",11188 => "01010000",11189 => "11011111",11190 => "11011110",11191 => "01110110",11192 => "10110111",11193 => "11001001",11194 => "10010010",11195 => "01011001",11196 => "00111100",11197 => "01000001",11198 => "01001010",11199 => "10100000",11200 => "10111110",11201 => "00101111",11202 => "11010011",11203 => "11100111",11204 => "00101100",11205 => "11101010",11206 => "10101001",11207 => "00011010",11208 => "01111101",11209 => "11000101",11210 => "01011010",11211 => "11010110",11212 => "10100000",11213 => "10101001",11214 => "11000010",11215 => "00000001",11216 => "10000110",11217 => "00001100",11218 => "11011010",11219 => "01001110",11220 => "10100100",11221 => "01011111",11222 => "11010010",11223 => "11011101",11224 => "11100110",11225 => "01001110",11226 => "10111000",11227 => "00100101",11228 => "01101110",11229 => "11001000",11230 => "10011000",11231 => "01100110",11232 => "01110000",11233 => "11011101",11234 => "00101010",11235 => "00000001",11236 => "01101111",11237 => "00001110",11238 => "00110010",11239 => "00110001",11240 => "11101010",11241 => "01011010",11242 => "00111010",11243 => "10001010",11244 => "11100101",11245 => "10110010",11246 => "10011100",11247 => "00101011",11248 => "11001111",11249 => "01110010",11250 => "10000000",11251 => "11100101",11252 => "01100101",11253 => "01010000",11254 => "11000011",11255 => "00110000",11256 => "00001010",11257 => "11001001",11258 => "01011110",11259 => "10011110",11260 => "01000110",11261 => "11100110",11262 => "00111101",11263 => "10100001",11264 => "01001100",11265 => "01111111",11266 => "11001001",11267 => "00100000",11268 => "10001100",11269 => "01101110",11270 => "00001111",11271 => "00000111",11272 => "11110100",11273 => "11101100",11274 => "10110101",11275 => "00111010",11276 => "11100101",11277 => "01011110",11278 => "01101001",11279 => "11101010",11280 => "11110000",11281 => "11000010",11282 => "10011010",11283 => "01011001",11284 => "01101101",11285 => "11101110",11286 => "01000000",11287 => "11110001",11288 => "01000001",11289 => "10010110",11290 => "11011111",11291 => "01011010",11292 => "00101011",11293 => "01010100",11294 => "01000001",11295 => "00011010",11296 => "01110100",11297 => "00100011",11298 => "00111111",11299 => "11110101",11300 => "01100100",11301 => "10010110",11302 => "01010000",11303 => "11101111",11304 => "00100100",11305 => "10110101",11306 => "01101001",11307 => "11000000",11308 => "11011111",11309 => "10010010",11310 => "11001000",11311 => "11111010",11312 => "10001001",11313 => "01011000",11314 => "01010001",11315 => "00001011",11316 => "11011011",11317 => "01101111",11318 => "11010000",11319 => "10110010",11320 => "00101111",11321 => "11111011",11322 => "00011000",11323 => "11111101",11324 => "00001011",11325 => "01101111",11326 => "11000111",11327 => "10111111",11328 => "01001010",11329 => "10110111",11330 => "11010001",11331 => "00110010",11332 => "00100110",11333 => "10101010",11334 => "01000101",11335 => "11010011",11336 => "11100101",11337 => "01100101",11338 => "11101010",11339 => "10110100",11340 => "10110000",11341 => "11101010",11342 => "00101000",11343 => "01000011",11344 => "01010000",11345 => "11001001",11346 => "11011000",11347 => "10100001",11348 => "11000000",11349 => "01000011",11350 => "11011010",11351 => "00110011",11352 => "00000000",11353 => "00011101",11354 => "01010101",11355 => "00001111",11356 => "01110111",11357 => "01000110",11358 => "01010011",11359 => "01000000",11360 => "11111000",11361 => "00011010",11362 => "11101100",11363 => "11000100",11364 => "00011111",11365 => "01010111",11366 => "11100111",11367 => "11010010",11368 => "00000110",11369 => "11010011",11370 => "01000110",11371 => "10101101",11372 => "00000000",11373 => "11010010",11374 => "01001110",11375 => "00110101",11376 => "00001010",11377 => "00101011",11378 => "11101000",11379 => "10011000",11380 => "00100110",11381 => "11100100",11382 => "10000100",11383 => "01101000",11384 => "11111100",11385 => "00011100",11386 => "00011000",11387 => "10011111",11388 => "11101101",11389 => "10001010",11390 => "11100011",11391 => "11000011",11392 => "10001110",11393 => "01011110",11394 => "11001010",11395 => "00100110",11396 => "00111001",11397 => "11011100",11398 => "11110011",11399 => "01000110",11400 => "10010111",11401 => "11100001",11402 => "11101001",11403 => "01000100",11404 => "00101000",11405 => "10001010",11406 => "11001001",11407 => "11110100",11408 => "01101100",11409 => "00100001",11410 => "10100101",11411 => "01111101",11412 => "00111101",11413 => "11010111",11414 => "00000111",11415 => "10110110",11416 => "00010110",11417 => "10010101",11418 => "11011101",11419 => "01000101",11420 => "00110001",11421 => "01000111",11422 => "11111000",11423 => "10111001",11424 => "11100011",11425 => "01111100",11426 => "11000110",11427 => "00111001",11428 => "10011001",11429 => "01011100",11430 => "00100111",11431 => "11111111",11432 => "01001000",11433 => "11001000",11434 => "10111011",11435 => "11101101",11436 => "10101010",11437 => "11011101",11438 => "00101101",11439 => "11010111",11440 => "00011010",11441 => "10011110",11442 => "00011011",11443 => "10101011",11444 => "10100000",11445 => "00011100",11446 => "10110000",11447 => "11101110",11448 => "10101110",11449 => "10001110",11450 => "00011010",11451 => "10110000",11452 => "11000010",11453 => "00100000",11454 => "00100111",11455 => "01000001",11456 => "01110111",11457 => "10001010",11458 => "01110110",11459 => "01011000",11460 => "00010010",11461 => "11110000",11462 => "01100111",11463 => "00011001",11464 => "10100010",11465 => "10001001",11466 => "00111000",11467 => "11001101",11468 => "00100010",11469 => "11000101",11470 => "01011011",11471 => "11000011",11472 => "11000110",11473 => "01101110",11474 => "01101001",11475 => "00001011",11476 => "10001110",11477 => "10101110",11478 => "00011001",11479 => "10110111",11480 => "10010111",11481 => "11011010",11482 => "11011010",11483 => "01000010",11484 => "11111110",11485 => "10001100",11486 => "11100010",11487 => "00100110",11488 => "00100000",11489 => "11111010",11490 => "01111111",11491 => "00110110",11492 => "10001101",11493 => "01101011",11494 => "00111100",11495 => "01000100",11496 => "00100101",11497 => "01100100",11498 => "10000010",11499 => "11111100",11500 => "11110001",11501 => "11010101",11502 => "10000100",11503 => "00001111",11504 => "10100100",11505 => "00010001",11506 => "10111010",11507 => "10100101",11508 => "01111011",11509 => "11010001",11510 => "10000111",11511 => "11000010",11512 => "01000000",11513 => "11010110",11514 => "00010111",11515 => "10010011",11516 => "11010001",11517 => "10101011",11518 => "00001001",11519 => "01001101",11520 => "00111001",11521 => "01100100",11522 => "00010000",11523 => "00111000",11524 => "00100111",11525 => "01011001",11526 => "01100111",11527 => "11001100",11528 => "10110001",11529 => "11111001",11530 => "10101101",11531 => "01011000",11532 => "00100110",11533 => "00010001",11534 => "10110100",11535 => "11001010",11536 => "01100110",11537 => "01000110",11538 => "11000101",11539 => "11011111",11540 => "00111010",11541 => "00111001",11542 => "10111110",11543 => "00001010",11544 => "01011001",11545 => "10000111",11546 => "01111010",11547 => "10100001",11548 => "00111100",11549 => "01001101",11550 => "01000010",11551 => "11110010",11552 => "00000110",11553 => "11011111",11554 => "00111100",11555 => "00110010",11556 => "00110010",11557 => "11101010",11558 => "00111110",11559 => "00110011",11560 => "00111100",11561 => "10110110",11562 => "11100000",11563 => "00011101",11564 => "11010001",11565 => "00100011",11566 => "11111010",11567 => "01010101",11568 => "10001000",11569 => "01111110",11570 => "00110001",11571 => "01101111",11572 => "00111001",11573 => "00010010",11574 => "01010110",11575 => "01001001",11576 => "00110101",11577 => "00110010",11578 => "10010011",11579 => "00111110",11580 => "01110000",11581 => "00111110",11582 => "10000010",11583 => "10000010",11584 => "01010110",11585 => "01101100",11586 => "11001000",11587 => "11100000",11588 => "11110001",11589 => "01100110",11590 => "11000101",11591 => "10000011",11592 => "11100011",11593 => "10010110",11594 => "00101101",11595 => "10100010",11596 => "00111001",11597 => "11111100",11598 => "01111111",11599 => "01010110",11600 => "11100111",11601 => "11101111",11602 => "11011111",11603 => "01001101",11604 => "01010011",11605 => "11101110",11606 => "11110010",11607 => "11011011",11608 => "00111000",11609 => "10100010",11610 => "00000100",11611 => "10110101",11612 => "00010111",11613 => "11101100",11614 => "01001111",11615 => "11100111",11616 => "10111110",11617 => "01111000",11618 => "00011110",11619 => "00101000",11620 => "01111110",11621 => "00110110",11622 => "10001001",11623 => "00110100",11624 => "00011100",11625 => "01001001",11626 => "00111110",11627 => "11011110",11628 => "00100011",11629 => "11111110",11630 => "00000100",11631 => "10100101",11632 => "00010110",11633 => "01101101",11634 => "01111001",11635 => "00101011",11636 => "00100010",11637 => "11000010",11638 => "10011100",11639 => "11011010",11640 => "01110111",11641 => "11110001",11642 => "11110010",11643 => "11010000",11644 => "11101010",11645 => "00000000",11646 => "11100011",11647 => "10010000",11648 => "01110110",11649 => "10111010",11650 => "10010001",11651 => "10010000",11652 => "11110111",11653 => "10110110",11654 => "00011001",11655 => "01010010",11656 => "00000000",11657 => "00001101",11658 => "01100101",11659 => "01000111",11660 => "10110001",11661 => "10100100",11662 => "11110111",11663 => "00100111",11664 => "01100011",11665 => "00011100",11666 => "10101001",11667 => "11111100",11668 => "00101010",11669 => "00011111",11670 => "00101100",11671 => "11000111",11672 => "11010110",11673 => "01011110",11674 => "11000110",11675 => "11011110",11676 => "10110110",11677 => "01000010",11678 => "10000111",11679 => "01101011",11680 => "01100001",11681 => "10011101",11682 => "11111010",11683 => "01111000",11684 => "00110100",11685 => "11101110",11686 => "10110010",11687 => "01111010",11688 => "11011001",11689 => "11110100",11690 => "10101101",11691 => "00000001",11692 => "11011000",11693 => "11011101",11694 => "00100001",11695 => "01000000",11696 => "01000111",11697 => "00000101",11698 => "01101011",11699 => "11001010",11700 => "00010000",11701 => "11010001",11702 => "01100100",11703 => "11001101",11704 => "10101011",11705 => "10100001",11706 => "00111101",11707 => "10011101",11708 => "00010011",11709 => "10100101",11710 => "11111011",11711 => "01100111",11712 => "11010011",11713 => "11011000",11714 => "00010111",11715 => "01000100",11716 => "10011010",11717 => "00001100",11718 => "10010110",11719 => "10111110",11720 => "10111100",11721 => "01010111",11722 => "11011111",11723 => "11000010",11724 => "01010101",11725 => "11101001",11726 => "00101100",11727 => "00100111",11728 => "01100111",11729 => "11100001",11730 => "01110000",11731 => "00111011",11732 => "10101011",11733 => "00000000",11734 => "11100111",11735 => "11101111",11736 => "00000111",11737 => "11011001",11738 => "00000001",11739 => "11110111",11740 => "01100100",11741 => "00011010",11742 => "00000001",11743 => "10110000",11744 => "10110011",11745 => "10000111",11746 => "11010101",11747 => "10011101",11748 => "01000001",11749 => "01100101",11750 => "11110101",11751 => "11111000",11752 => "11011110",11753 => "11110110",11754 => "11011100",11755 => "11101010",11756 => "00100011",11757 => "01110000",11758 => "11001010",11759 => "00001101",11760 => "01111001",11761 => "11100000",11762 => "00110000",11763 => "11100111",11764 => "11111111",11765 => "11100100",11766 => "10010101",11767 => "01000001",11768 => "00001101",11769 => "00100000",11770 => "10101010",11771 => "01010101",11772 => "11110011",11773 => "10010101",11774 => "10101111",11775 => "11111001",11776 => "11011111",11777 => "01011110",11778 => "10001111",11779 => "01100111",11780 => "11000111",11781 => "01100011",11782 => "01111000",11783 => "01111101",11784 => "00001111",11785 => "10111011",11786 => "00110011",11787 => "01110100",11788 => "01101101",11789 => "10000011",11790 => "01100110",11791 => "01000101",11792 => "11001010",11793 => "01101110",11794 => "11011110",11795 => "10010000",11796 => "10110010",11797 => "10111110",11798 => "01001001",11799 => "00101011",11800 => "01101101",11801 => "11101100",11802 => "01000101",11803 => "11011111",11804 => "01101110",11805 => "11001100",11806 => "00010011",11807 => "11011101",11808 => "00011101",11809 => "00000100",11810 => "10101101",11811 => "11011100",11812 => "11001110",11813 => "10011100",11814 => "10001011",11815 => "10110111",11816 => "00111111",11817 => "01001011",11818 => "01111111",11819 => "11110000",11820 => "11110001",11821 => "11011110",11822 => "00110101",11823 => "01100010",11824 => "10001101",11825 => "10010010",11826 => "11011010",11827 => "11100011",11828 => "00011111",11829 => "10110011",11830 => "11000000",11831 => "01100001",11832 => "10000100",11833 => "11011011",11834 => "00000110",11835 => "10110111",11836 => "00010000",11837 => "10001101",11838 => "10000010",11839 => "10001000",11840 => "01011101",11841 => "01111001",11842 => "10010100",11843 => "11101000",11844 => "01010111",11845 => "01001010",11846 => "01000101",11847 => "10001110",11848 => "10000000",11849 => "00110001",11850 => "01011110",11851 => "01011100",11852 => "00011000",11853 => "00010011",11854 => "00111111",11855 => "11110001",11856 => "00001011",11857 => "00001010",11858 => "00001111",11859 => "01110101",11860 => "01010100",11861 => "11111100",11862 => "10001001",11863 => "00110110",11864 => "11111000",11865 => "11001101",11866 => "10110000",11867 => "00111101",11868 => "11111000",11869 => "01100111",11870 => "10010011",11871 => "01001001",11872 => "11011011",11873 => "00001011",11874 => "00111100",11875 => "10111001",11876 => "01000101",11877 => "00101010",11878 => "01010111",11879 => "01010110",11880 => "00000010",11881 => "01001000",11882 => "01100001",11883 => "10000000",11884 => "00011110",11885 => "10001001",11886 => "10000100",11887 => "00000100",11888 => "00100101",11889 => "01100111",11890 => "01001101",11891 => "11100000",11892 => "11101001",11893 => "00010101",11894 => "10000110",11895 => "01100101",11896 => "01011100",11897 => "00100000",11898 => "00110110",11899 => "10010011",11900 => "00101010",11901 => "10100000",11902 => "01000001",11903 => "11011101",11904 => "01010101",11905 => "11000001",11906 => "01110001",11907 => "01111110",11908 => "01010001",11909 => "10001000",11910 => "10101111",11911 => "01110000",11912 => "00100111",11913 => "10100010",11914 => "00100010",11915 => "01110100",11916 => "10110010",11917 => "01010000",11918 => "10011001",11919 => "00011011",11920 => "01000011",11921 => "10010111",11922 => "10010101",11923 => "01011101",11924 => "11101011",11925 => "10011101",11926 => "01110100",11927 => "00101110",11928 => "00000000",11929 => "10100001",11930 => "01110111",11931 => "01011011",11932 => "01111000",11933 => "00100110",11934 => "01011001",11935 => "01111110",11936 => "11111011",11937 => "11101001",11938 => "01100101",11939 => "11110001",11940 => "00011000",11941 => "10100110",11942 => "10101110",11943 => "00011111",11944 => "01110010",11945 => "11000110",11946 => "10001010",11947 => "11100011",11948 => "01010000",11949 => "01100010",11950 => "10001000",11951 => "11010100",11952 => "00010111",11953 => "11001111",11954 => "01100110",11955 => "00101110",11956 => "10101100",11957 => "00100000",11958 => "10110100",11959 => "00101000",11960 => "11001001",11961 => "00001000",11962 => "11101110",11963 => "10101101",11964 => "01010110",11965 => "00010101",11966 => "11100101",11967 => "00011000",11968 => "11110010",11969 => "01110000",11970 => "01011001",11971 => "00100010",11972 => "00011100",11973 => "11010010",11974 => "11111101",11975 => "01010001",11976 => "00110011",11977 => "00110000",11978 => "10000001",11979 => "01011011",11980 => "10011110",11981 => "10000011",11982 => "10010000",11983 => "11011000",11984 => "01011001",11985 => "10010101",11986 => "00110001",11987 => "11001010",11988 => "01000100",11989 => "01101101",11990 => "11010111",11991 => "11110010",11992 => "01111000",11993 => "01011011",11994 => "10011110",11995 => "10101001",11996 => "10110111",11997 => "11110110",11998 => "11011000",11999 => "10111100",12000 => "01101110",12001 => "01010111",12002 => "00010111",12003 => "00011100",12004 => "01001101",12005 => "11110111",12006 => "10001010",12007 => "01110101",12008 => "01110111",12009 => "00110011",12010 => "10110001",12011 => "00001111",12012 => "01010100",12013 => "01100011",12014 => "01100010",12015 => "11011101",12016 => "11010001",12017 => "01001110",12018 => "00110011",12019 => "10100101",12020 => "10001100",12021 => "10110110",12022 => "10110010",12023 => "01100100",12024 => "00001101",12025 => "01100010",12026 => "10010011",12027 => "11010010",12028 => "10011101",12029 => "11001000",12030 => "11111101",12031 => "10000010",12032 => "01010011",12033 => "00111000",12034 => "00101110",12035 => "00110000",12036 => "01101001",12037 => "10001000",12038 => "00001001",12039 => "10110110",12040 => "11010000",12041 => "10000001",12042 => "01001111",12043 => "10010100",12044 => "00101001",12045 => "11111111",12046 => "01010101",12047 => "11110000",12048 => "00000111",12049 => "01001100",12050 => "01001101",12051 => "00000000",12052 => "00001100",12053 => "01011110",12054 => "11001011",12055 => "00110010",12056 => "11101000",12057 => "11001111",12058 => "11110000",12059 => "10010101",12060 => "10011000",12061 => "01100011",12062 => "10000100",12063 => "11001010",12064 => "00101111",12065 => "00100111",12066 => "01011100",12067 => "11111101",12068 => "11111100",12069 => "10011110",12070 => "00111001",12071 => "00111100",12072 => "01011101",12073 => "11010000",12074 => "10101110",12075 => "11011100",12076 => "10110010",12077 => "00100110",12078 => "11011001",12079 => "10100001",12080 => "11110110",12081 => "00110000",12082 => "10000010",12083 => "00010011",12084 => "10101111",12085 => "01101001",12086 => "10110100",12087 => "00100110",12088 => "10010110",12089 => "00110000",12090 => "10111101",12091 => "10101110",12092 => "10101000",12093 => "10100001",12094 => "01000000",12095 => "11100011",12096 => "11000010",12097 => "01111000",12098 => "01101110",12099 => "11001000",12100 => "00100100",12101 => "10010101",12102 => "11001000",12103 => "00010101",12104 => "11011110",12105 => "10110111",12106 => "11011010",12107 => "10001100",12108 => "00000101",12109 => "01010000",12110 => "11110011",12111 => "10101010",12112 => "11001100",12113 => "01111010",12114 => "10010011",12115 => "10111001",12116 => "00000111",12117 => "00101111",12118 => "11011001",12119 => "10111111",12120 => "01011011",12121 => "01101010",12122 => "01001011",12123 => "01101011",12124 => "00000011",12125 => "01111000",12126 => "01001101",12127 => "01101001",12128 => "01000101",12129 => "10110111",12130 => "00011111",12131 => "10010010",12132 => "11111100",12133 => "10010000",12134 => "10100111",12135 => "10010111",12136 => "11100010",12137 => "00011101",12138 => "00101001",12139 => "00000001",12140 => "00101110",12141 => "00011110",12142 => "00111001",12143 => "10001101",12144 => "11010101",12145 => "00010000",12146 => "00111000",12147 => "00000110",12148 => "00111100",12149 => "11111001",12150 => "10111111",12151 => "01111000",12152 => "01010100",12153 => "01000000",12154 => "01010001",12155 => "10111000",12156 => "10001111",12157 => "10101011",12158 => "11100110",12159 => "01110111",12160 => "00000011",12161 => "00111101",12162 => "10001011",12163 => "11100101",12164 => "11101100",12165 => "01000111",12166 => "00000011",12167 => "01110000",12168 => "10100111",12169 => "10011110",12170 => "01110001",12171 => "11100110",12172 => "01110010",12173 => "00011011",12174 => "01110101",12175 => "01011110",12176 => "11001001",12177 => "01001011",12178 => "01101100",12179 => "11110010",12180 => "00110001",12181 => "11010010",12182 => "11110101",12183 => "01001011",12184 => "11011111",12185 => "01110010",12186 => "11100000",12187 => "01111011",12188 => "01110010",12189 => "01110001",12190 => "01011011",12191 => "00000111",12192 => "11001100",12193 => "00111000",12194 => "00001001",12195 => "11000011",12196 => "10000101",12197 => "00000100",12198 => "00010100",12199 => "10101010",12200 => "11111100",12201 => "11101101",12202 => "00111110",12203 => "10111101",12204 => "10000000",12205 => "11010110",12206 => "11000100",12207 => "10011110",12208 => "10010100",12209 => "11110001",12210 => "00111110",12211 => "01001011",12212 => "01101001",12213 => "01010111",12214 => "10101001",12215 => "00111010",12216 => "00110111",12217 => "11001101",12218 => "00110010",12219 => "01111111",12220 => "11001011",12221 => "01110111",12222 => "01011010",12223 => "01011100",12224 => "11011111",12225 => "11010010",12226 => "11001010",12227 => "10100010",12228 => "01011000",12229 => "01111010",12230 => "10101000",12231 => "01000110",12232 => "11000010",12233 => "01001101",12234 => "10001000",12235 => "10111110",12236 => "01011101",12237 => "11100011",12238 => "00110001",12239 => "01110110",12240 => "01001110",12241 => "11110001",12242 => "11111000",12243 => "01011111",12244 => "01000000",12245 => "00111001",12246 => "00010001",12247 => "11001010",12248 => "11101100",12249 => "11011010",12250 => "00101000",12251 => "00001110",12252 => "00001111",12253 => "10010001",12254 => "10100010",12255 => "00001000",12256 => "01100111",12257 => "10011111",12258 => "01101111",12259 => "01001100",12260 => "10110110",12261 => "01010110",12262 => "10010010",12263 => "11100011",12264 => "01010111",12265 => "01100010",12266 => "00100100",12267 => "11001010",12268 => "00110011",12269 => "01110110",12270 => "01000000",12271 => "11011001",12272 => "11010101",12273 => "11011100",12274 => "01101110",12275 => "10000000",12276 => "00110110",12277 => "00011110",12278 => "10100001",12279 => "10000101",12280 => "10110011",12281 => "01101111",12282 => "11001001",12283 => "11001100",12284 => "01111010",12285 => "11001101",12286 => "00000010",12287 => "11011001",12288 => "10101000",12289 => "11001101",12290 => "10100000",12291 => "01001001",12292 => "00011110",12293 => "10100111",12294 => "11011100",12295 => "00100010",12296 => "01001111",12297 => "10000111",12298 => "00111000",12299 => "01000000",12300 => "11010010",12301 => "11100101",12302 => "10000100",12303 => "01110101",12304 => "10001010",12305 => "00100100",12306 => "11000110",12307 => "00010110",12308 => "00110111",12309 => "01101001",12310 => "11001100",12311 => "10010000",12312 => "01001000",12313 => "10101101",12314 => "10110101",12315 => "10010111",12316 => "10110100",12317 => "00100101",12318 => "11000011",12319 => "01101000",12320 => "01110100",12321 => "11100111",12322 => "00110000",12323 => "01101011",12324 => "01011100",12325 => "00000100",12326 => "10000100",12327 => "00111100",12328 => "11110011",12329 => "10000011",12330 => "01110111",12331 => "11011000",12332 => "10110110",12333 => "11101110",12334 => "01001011",12335 => "11101011",12336 => "01111110",12337 => "10011111",12338 => "00000010",12339 => "00001010",12340 => "10001101",12341 => "11100100",12342 => "10011111",12343 => "01110110",12344 => "00100110",12345 => "00001010",12346 => "10101010",12347 => "00101111",12348 => "11100101",12349 => "00000100",12350 => "11001110",12351 => "01000001",12352 => "11001011",12353 => "00101000",12354 => "11001111",12355 => "11100001",12356 => "01001110",12357 => "00001000",12358 => "00001001",12359 => "00010101",12360 => "01100001",12361 => "11111010",12362 => "11100110",12363 => "00011101",12364 => "10000100",12365 => "00101101",12366 => "00001000",12367 => "01010010",12368 => "01001010",12369 => "01001011",12370 => "11010110",12371 => "10001101",12372 => "00010100",12373 => "01100011",12374 => "01111111",12375 => "10101100",12376 => "10011101",12377 => "01110100",12378 => "01111111",12379 => "11001101",12380 => "00101101",12381 => "11111010",12382 => "00101000",12383 => "01001011",12384 => "10000011",12385 => "11110001",12386 => "11101100",12387 => "10100110",12388 => "11010101",12389 => "11101110",12390 => "01000100",12391 => "00000000",12392 => "11010101",12393 => "11011011",12394 => "01001111",12395 => "10111001",12396 => "10101110",12397 => "11101110",12398 => "11100101",12399 => "11101000",12400 => "11010011",12401 => "01010010",12402 => "00011100",12403 => "00101010",12404 => "00011100",12405 => "10000001",12406 => "10010101",12407 => "00101110",12408 => "00001101",12409 => "11111011",12410 => "00101000",12411 => "10101010",12412 => "00000110",12413 => "10111001",12414 => "01110101",12415 => "11011101",12416 => "11111001",12417 => "11010101",12418 => "11100110",12419 => "11001100",12420 => "11000101",12421 => "11110111",12422 => "00101110",12423 => "00101101",12424 => "11011000",12425 => "11011001",12426 => "11100010",12427 => "00001010",12428 => "10001101",12429 => "11101011",12430 => "10100010",12431 => "11001001",12432 => "00101011",12433 => "11001111",12434 => "11101000",12435 => "01100110",12436 => "01100111",12437 => "11011110",12438 => "00000000",12439 => "01000010",12440 => "00101101",12441 => "11101010",12442 => "11101110",12443 => "10111111",12444 => "00000110",12445 => "00110011",12446 => "11001000",12447 => "10110110",12448 => "11101000",12449 => "00011101",12450 => "01100110",12451 => "10011001",12452 => "00011001",12453 => "10110000",12454 => "00111011",12455 => "00110001",12456 => "10110101",12457 => "00011100",12458 => "11101010",12459 => "00000011",12460 => "11111111",12461 => "01001001",12462 => "01100100",12463 => "11101110",12464 => "01110100",12465 => "00011011",12466 => "01011011",12467 => "10000000",12468 => "10100001",12469 => "00101110",12470 => "10101100",12471 => "01001110",12472 => "11000000",12473 => "01011000",12474 => "10101001",12475 => "11001011",12476 => "01110110",12477 => "01110001",12478 => "00000011",12479 => "01001101",12480 => "00110101",12481 => "11111011",12482 => "10010001",12483 => "01011110",12484 => "01010100",12485 => "11100000",12486 => "00110100",12487 => "10110100",12488 => "11001000",12489 => "10011110",12490 => "11001101",12491 => "01100101",12492 => "10010111",12493 => "11100110",12494 => "11010100",12495 => "00110011",12496 => "11100011",12497 => "10111000",12498 => "00101000",12499 => "00010010",12500 => "11010001",12501 => "00101101",12502 => "00100000",12503 => "01111001",12504 => "00011100",12505 => "11011000",12506 => "00111101",12507 => "10101100",12508 => "01001001",12509 => "10100010",12510 => "00100111",12511 => "00111000",12512 => "11000010",12513 => "01010010",12514 => "01010100",12515 => "01111001",12516 => "00001111",12517 => "11010110",12518 => "00101011",12519 => "11100010",12520 => "01100100",12521 => "01010110",12522 => "11011000",12523 => "00010100",12524 => "00001000",12525 => "00011111",12526 => "00011101",12527 => "10010110",12528 => "01011011",12529 => "11110011",12530 => "11111001",12531 => "01101101",12532 => "10001100",12533 => "11000001",12534 => "01010000",12535 => "00001001",12536 => "00111110",12537 => "01001000",12538 => "10011101",12539 => "01100101",12540 => "11111010",12541 => "01011101",12542 => "00110101",12543 => "11101000",12544 => "00111010",12545 => "00001111",12546 => "00111010",12547 => "00001011",12548 => "00100110",12549 => "10011101",12550 => "00010010",12551 => "01000100",12552 => "00001010",12553 => "00011100",12554 => "10001100",12555 => "11011001",12556 => "11011000",12557 => "00100101",12558 => "00010001",12559 => "00010101",12560 => "00000001",12561 => "10011011",12562 => "01101011",12563 => "01111011",12564 => "11101100",12565 => "10010011",12566 => "01011011",12567 => "10010111",12568 => "00100111",12569 => "00110100",12570 => "00011011",12571 => "10101010",12572 => "11111110",12573 => "11110001",12574 => "00010000",12575 => "01001110",12576 => "00110111",12577 => "00110111",12578 => "01000001",12579 => "01000000",12580 => "10000000",12581 => "00101010",12582 => "10001100",12583 => "10110100",12584 => "10100100",12585 => "01001001",12586 => "00010001",12587 => "01011011",12588 => "01110100",12589 => "10001000",12590 => "01101110",12591 => "10101100",12592 => "10010100",12593 => "10100000",12594 => "00010001",12595 => "00100111",12596 => "11011001",12597 => "11101000",12598 => "10100010",12599 => "11001000",12600 => "10110110",12601 => "00110110",12602 => "01101001",12603 => "01001101",12604 => "11100000",12605 => "00001010",12606 => "00010101",12607 => "10101110",12608 => "00101011",12609 => "10110110",12610 => "00000111",12611 => "11111110",12612 => "00000001",12613 => "10110110",12614 => "01111100",12615 => "01111101",12616 => "10111011",12617 => "01000001",12618 => "00011011",12619 => "00010100",12620 => "01100110",12621 => "01101011",12622 => "00110000",12623 => "00100101",12624 => "00000110",12625 => "00010010",12626 => "00001000",12627 => "10111000",12628 => "11000110",12629 => "10101100",12630 => "10101011",12631 => "10110100",12632 => "00111011",12633 => "01110100",12634 => "00100101",12635 => "01010101",12636 => "00010110",12637 => "01011101",12638 => "10111100",12639 => "00110001",12640 => "00001110",12641 => "01010110",12642 => "01100010",12643 => "00101101",12644 => "10000111",12645 => "11110100",12646 => "01111001",12647 => "10110000",12648 => "10010011",12649 => "00101110",12650 => "00010100",12651 => "10001111",12652 => "10001100",12653 => "00000010",12654 => "10100110",12655 => "00010110",12656 => "00000001",12657 => "00100001",12658 => "11001001",12659 => "01100101",12660 => "01101011",12661 => "01111111",12662 => "00110010",12663 => "01001010",12664 => "10110000",12665 => "11011001",12666 => "00101100",12667 => "11000010",12668 => "10011110",12669 => "10101001",12670 => "11000110",12671 => "10111101",12672 => "01101110",12673 => "01101111",12674 => "10110110",12675 => "01111010",12676 => "10010000",12677 => "10100100",12678 => "01010111",12679 => "00110010",12680 => "11001101",12681 => "11001100",12682 => "10010010",12683 => "10111100",12684 => "00110111",12685 => "01110111",12686 => "11111101",12687 => "01001101",12688 => "01101100",12689 => "10010010",12690 => "11111001",12691 => "00100000",12692 => "00110010",12693 => "11100000",12694 => "00111101",12695 => "00111010",12696 => "00100001",12697 => "00011110",12698 => "11011111",12699 => "01101100",12700 => "10101111",12701 => "01000101",12702 => "00001011",12703 => "00000010",12704 => "11000011",12705 => "10100100",12706 => "01011111",12707 => "01011110",12708 => "11110001",12709 => "10100010",12710 => "10000101",12711 => "00001001",12712 => "10111001",12713 => "11111101",12714 => "10000011",12715 => "11111100",12716 => "11011011",12717 => "10011100",12718 => "10011101",12719 => "10111100",12720 => "11010010",12721 => "01011110",12722 => "01010110",12723 => "10010000",12724 => "10101110",12725 => "01000100",12726 => "10010001",12727 => "11111111",12728 => "11010011",12729 => "10010001",12730 => "00100010",12731 => "10010011",12732 => "11001111",12733 => "11000011",12734 => "01101111",12735 => "01101001",12736 => "11000011",12737 => "00111010",12738 => "10001001",12739 => "00110110",12740 => "00000111",12741 => "10101000",12742 => "11001100",12743 => "11000001",12744 => "01010101",12745 => "10000011",12746 => "10111111",12747 => "01110000",12748 => "10000010",12749 => "11101001",12750 => "00011110",12751 => "10101101",12752 => "10001010",12753 => "00111000",12754 => "11101101",12755 => "01010111",12756 => "10110110",12757 => "11100001",12758 => "01111001",12759 => "01010000",12760 => "00111011",12761 => "11110111",12762 => "10101011",12763 => "01100001",12764 => "01111110",12765 => "11100111",12766 => "11101001",12767 => "00001000",12768 => "10000110",12769 => "10111110",12770 => "01110011",12771 => "00110101",12772 => "11100000",12773 => "11011010",12774 => "11011100",12775 => "00101011",12776 => "10000110",12777 => "10111101",12778 => "10000110",12779 => "11001101",12780 => "00000001",12781 => "01110101",12782 => "01110000",12783 => "11111101",12784 => "11001111",12785 => "11011111",12786 => "10101001",12787 => "00010101",12788 => "11111010",12789 => "11101101",12790 => "00010101",12791 => "01000001",12792 => "11010100",12793 => "11001101",12794 => "11010110",12795 => "00001110",12796 => "00001101",12797 => "00001011",12798 => "01110000",12799 => "00110010",12800 => "01010100",12801 => "11110000",12802 => "00111111",12803 => "10101111",12804 => "11001100",12805 => "10001111",12806 => "00100100",12807 => "10000111",12808 => "11010111",12809 => "10010000",12810 => "00101111",12811 => "11100100",12812 => "10111100",12813 => "10010010",12814 => "00001101",12815 => "10011010",12816 => "10111111",12817 => "10010000",12818 => "11100011",12819 => "00010101",12820 => "11100111",12821 => "10011101",12822 => "10001000",12823 => "10111011",12824 => "11111101",12825 => "01010000",12826 => "11100100",12827 => "00011011",12828 => "11100100",12829 => "00011111",12830 => "11010010",12831 => "00000101",12832 => "10010011",12833 => "00011110",12834 => "10110010",12835 => "10100101",12836 => "00110011",12837 => "10110001",12838 => "11010011",12839 => "01110010",12840 => "01000011",12841 => "01111111",12842 => "00000000",12843 => "01100010",12844 => "00001110",12845 => "11111011",12846 => "00001001",12847 => "01110000",12848 => "10100100",12849 => "11110111",12850 => "01000110",12851 => "10010000",12852 => "01110100",12853 => "00110011",12854 => "00010010",12855 => "10010101",12856 => "10000010",12857 => "01100011",12858 => "10001111",12859 => "01000000",12860 => "11111101",12861 => "01100101",12862 => "01111000",12863 => "00010110",12864 => "10001011",12865 => "01011101",12866 => "10010101",12867 => "01011011",12868 => "00010101",12869 => "10011111",12870 => "10101101",12871 => "00001010",12872 => "00100000",12873 => "00011100",12874 => "01000010",12875 => "00001010",12876 => "11100000",12877 => "11010011",12878 => "10110111",12879 => "01000000",12880 => "10000110",12881 => "00100110",12882 => "10111011",12883 => "11100111",12884 => "10110011",12885 => "10011110",12886 => "10111101",12887 => "10011100",12888 => "00110000",12889 => "01100001",12890 => "01011010",12891 => "10010000",12892 => "01111111",12893 => "11011010",12894 => "10011100",12895 => "10010011",12896 => "10110101",12897 => "10000101",12898 => "01101101",12899 => "10101000",12900 => "00000111",12901 => "01000111",12902 => "10000010",12903 => "01110011",12904 => "01000011",12905 => "01001000",12906 => "10010110",12907 => "01100111",12908 => "11101110",12909 => "10100010",12910 => "11101101",12911 => "11100110",12912 => "01110100",12913 => "00010110",12914 => "01101100",12915 => "10111110",12916 => "01000011",12917 => "01110100",12918 => "00101101",12919 => "11000000",12920 => "10001101",12921 => "11111000",12922 => "11111101",12923 => "01100011",12924 => "11001000",12925 => "01011100",12926 => "00010000",12927 => "11110010",12928 => "10111101",12929 => "11111011",12930 => "11110110",12931 => "10111110",12932 => "00000110",12933 => "01100100",12934 => "01001010",12935 => "01110101",12936 => "11011010",12937 => "10001001",12938 => "01101011",12939 => "10101101",12940 => "11000000",12941 => "11001111",12942 => "01111101",12943 => "11001010",12944 => "00000100",12945 => "10101001",12946 => "10001110",12947 => "11001101",12948 => "11010011",12949 => "00111110",12950 => "10100111",12951 => "10111100",12952 => "00010100",12953 => "00000001",12954 => "00011001",12955 => "00010100",12956 => "00001010",12957 => "00000100",12958 => "01010110",12959 => "00100000",12960 => "00011001",12961 => "10111110",12962 => "01100001",12963 => "11010100",12964 => "00011000",12965 => "11111010",12966 => "01011101",12967 => "00110101",12968 => "00001100",12969 => "10000111",12970 => "00110010",12971 => "11000101",12972 => "01000110",12973 => "00111101",12974 => "01111100",12975 => "10111101",12976 => "01101111",12977 => "01100001",12978 => "10000000",12979 => "10111100",12980 => "01101011",12981 => "01101000",12982 => "11001110",12983 => "00011000",12984 => "01000011",12985 => "10100100",12986 => "10100101",12987 => "00011010",12988 => "00010000",12989 => "00001000",12990 => "11101010",12991 => "01001111",12992 => "01100010",12993 => "00101000",12994 => "10110111",12995 => "00000100",12996 => "11100110",12997 => "10000100",12998 => "11110011",12999 => "00111001",13000 => "11101011",13001 => "10101000",13002 => "01010100",13003 => "11100100",13004 => "10101110",13005 => "01111001",13006 => "00100001",13007 => "10100110",13008 => "01100000",13009 => "10001000",13010 => "10110111",13011 => "10001100",13012 => "01110011",13013 => "00001010",13014 => "10000010",13015 => "11011110",13016 => "11101010",13017 => "10111001",13018 => "00011100",13019 => "11010010",13020 => "00001110",13021 => "10000101",13022 => "11000111",13023 => "10011101",13024 => "00111111",13025 => "10111100",13026 => "01000110",13027 => "11010001",13028 => "00010111",13029 => "01100111",13030 => "00001011",13031 => "01110010",13032 => "10001010",13033 => "11010010",13034 => "01011000",13035 => "01011000",13036 => "10011011",13037 => "11011010",13038 => "00101001",13039 => "10001001",13040 => "10110010",13041 => "10000101",13042 => "10110111",13043 => "00000000",13044 => "01100001",13045 => "01110001",13046 => "11000101",13047 => "11101011",13048 => "10101010",13049 => "01100000",13050 => "11110111",13051 => "00101101",13052 => "00111011",13053 => "00011110",13054 => "00010101",13055 => "00111000",13056 => "00001010",13057 => "01100001",13058 => "10011111",13059 => "00110110",13060 => "01011000",13061 => "00111111",13062 => "11000011",13063 => "01110011",13064 => "00110101",13065 => "11111010",13066 => "00100011",13067 => "11101010",13068 => "01101101",13069 => "00110010",13070 => "11110000",13071 => "00101100",13072 => "01000110",13073 => "00100101",13074 => "01000111",13075 => "10100000",13076 => "11101100",13077 => "01011111",13078 => "10011001",13079 => "11111011",13080 => "00100100",13081 => "11101010",13082 => "01101000",13083 => "00101001",13084 => "00011010",13085 => "00101001",13086 => "01010011",13087 => "01011100",13088 => "00010010",13089 => "11100010",13090 => "10010101",13091 => "01001100",13092 => "00110101",13093 => "10110001",13094 => "01111100",13095 => "10001010",13096 => "00000000",13097 => "01001111",13098 => "00000100",13099 => "11010111",13100 => "11110100",13101 => "00010101",13102 => "11111001",13103 => "10000011",13104 => "10001110",13105 => "00001001",13106 => "10100110",13107 => "11111001",13108 => "00110110",13109 => "01110001",13110 => "11000010",13111 => "10000111",13112 => "10111100",13113 => "00011010",13114 => "10000110",13115 => "11101110",13116 => "11111110",13117 => "00110111",13118 => "01110101",13119 => "00110010",13120 => "10110101",13121 => "01010010",13122 => "11000101",13123 => "01000011",13124 => "00101101",13125 => "01011111",13126 => "00000100",13127 => "10001010",13128 => "01100010",13129 => "01010001",13130 => "00011011",13131 => "00111000",13132 => "10010001",13133 => "11111111",13134 => "00010000",13135 => "01110110",13136 => "10101010",13137 => "00110100",13138 => "10011011",13139 => "10101111",13140 => "10101001",13141 => "01010101",13142 => "01110101",13143 => "01111100",13144 => "01001001",13145 => "10110110",13146 => "11000011",13147 => "01001100",13148 => "10000101",13149 => "10010101",13150 => "10111110",13151 => "01001111",13152 => "11010011",13153 => "10000010",13154 => "01001110",13155 => "10101110",13156 => "11000010",13157 => "11101001",13158 => "01000111",13159 => "00111001",13160 => "00110010",13161 => "00100001",13162 => "01010000",13163 => "11001110",13164 => "01000010",13165 => "01101000",13166 => "00100000",13167 => "01011000",13168 => "10111010",13169 => "11001100",13170 => "11001110",13171 => "01000111",13172 => "11100110",13173 => "01111110",13174 => "00010110",13175 => "11001010",13176 => "01001000",13177 => "11011110",13178 => "11110111",13179 => "01001111",13180 => "00110001",13181 => "00000010",13182 => "10001011",13183 => "01010011",13184 => "00100000",13185 => "10101000",13186 => "10111010",13187 => "10111010",13188 => "00110010",13189 => "11001000",13190 => "01100001",13191 => "01111100",13192 => "01111000",13193 => "10000101",13194 => "00100111",13195 => "00101011",13196 => "00000001",13197 => "11111000",13198 => "00011011",13199 => "11011100",13200 => "11111001",13201 => "01000110",13202 => "01100000",13203 => "10111000",13204 => "10111011",13205 => "00011000",13206 => "11010011",13207 => "01110110",13208 => "10101100",13209 => "10010110",13210 => "11100111",13211 => "01101000",13212 => "01110011",13213 => "00001010",13214 => "10001101",13215 => "10110111",13216 => "00001111",13217 => "11011100",13218 => "10101000",13219 => "01000100",13220 => "01110001",13221 => "10110001",13222 => "11001010",13223 => "01010010",13224 => "10111101",13225 => "10111011",13226 => "10100100",13227 => "01001111",13228 => "01100011",13229 => "01111110",13230 => "10011111",13231 => "01000110",13232 => "00001111",13233 => "11010100",13234 => "01001110",13235 => "01001000",13236 => "11000110",13237 => "01000100",13238 => "01011110",13239 => "11110010",13240 => "00000101",13241 => "00000001",13242 => "00101000",13243 => "11110101",13244 => "01111010",13245 => "10000111",13246 => "01000110",13247 => "11000001",13248 => "01000101",13249 => "11000111",13250 => "10100000",13251 => "11101110",13252 => "10110101",13253 => "00001011",13254 => "00011110",13255 => "10011010",13256 => "10000001",13257 => "10000010",13258 => "11000110",13259 => "01100100",13260 => "00011001",13261 => "10000011",13262 => "10001010",13263 => "11001111",13264 => "01110011",13265 => "10000001",13266 => "10010010",13267 => "00001010",13268 => "10111110",13269 => "01100111",13270 => "10000111",13271 => "01110111",13272 => "10011100",13273 => "01001101",13274 => "01110110",13275 => "00010000",13276 => "10111100",13277 => "10100000",13278 => "01101010",13279 => "01100101",13280 => "00001000",13281 => "11010111",13282 => "00111011",13283 => "11111001",13284 => "11001001",13285 => "01010110",13286 => "11101111",13287 => "11010000",13288 => "11010011",13289 => "00000001",13290 => "01001101",13291 => "00100100",13292 => "11010000",13293 => "00111010",13294 => "10000000",13295 => "11010111",13296 => "00100001",13297 => "11101000",13298 => "11000110",13299 => "10011111",13300 => "00111011",13301 => "10101000",13302 => "00101010",13303 => "01101101",13304 => "00000000",13305 => "10001011",13306 => "01110011",13307 => "01011001",13308 => "10010100",13309 => "00110110",13310 => "10010010",13311 => "00110101",13312 => "11100110",13313 => "10110001",13314 => "11001111",13315 => "10011001",13316 => "00011000",13317 => "01110000",13318 => "01010011",13319 => "01001111",13320 => "10010111",13321 => "01010010",13322 => "11011101",13323 => "00011100",13324 => "01100000",13325 => "10000111",13326 => "01111000",13327 => "00100111",13328 => "11001111",13329 => "10100111",13330 => "10110011",13331 => "10000000",13332 => "11010000",13333 => "10001000",13334 => "10001010",13335 => "10100100",13336 => "01011001",13337 => "11100101",13338 => "00011101",13339 => "01110010",13340 => "11100101",13341 => "01100100",13342 => "11010101",13343 => "11011001",13344 => "11111101",13345 => "10101111",13346 => "11111101",13347 => "00010101",13348 => "11001110",13349 => "00011101",13350 => "11000101",13351 => "11111000",13352 => "01001111",13353 => "11000110",13354 => "00100100",13355 => "00101000",13356 => "10100000",13357 => "00011101",13358 => "11010001",13359 => "11000110",13360 => "00110011",13361 => "10010111",13362 => "11010101",13363 => "10101001",13364 => "10111111",13365 => "10100010",13366 => "01100111",13367 => "01111000",13368 => "10000111",13369 => "00011010",13370 => "00111101",13371 => "00111110",13372 => "10010000",13373 => "01111001",13374 => "00100000",13375 => "00100000",13376 => "11011011",13377 => "00000110",13378 => "11100100",13379 => "11110011",13380 => "11111101",13381 => "00110000",13382 => "11111000",13383 => "10111001",13384 => "10100101",13385 => "10001010",13386 => "11100000",13387 => "11110011",13388 => "11110111",13389 => "11011111",13390 => "01001000",13391 => "01011000",13392 => "01000010",13393 => "01010000",13394 => "00001001",13395 => "10110111",13396 => "01001100",13397 => "00111101",13398 => "10100001",13399 => "11100100",13400 => "01000011",13401 => "00111111",13402 => "00111101",13403 => "01011110",13404 => "10000000",13405 => "01100010",13406 => "10100100",13407 => "00110011",13408 => "01111010",13409 => "01000110",13410 => "00011101",13411 => "10000000",13412 => "01000100",13413 => "11010101",13414 => "11010110",13415 => "00110100",13416 => "11101110",13417 => "01000001",13418 => "11101011",13419 => "11111100",13420 => "11100000",13421 => "01000110",13422 => "01000010",13423 => "11000011",13424 => "11010111",13425 => "01011100",13426 => "01110101",13427 => "00000011",13428 => "01000000",13429 => "10001011",13430 => "11111011",13431 => "11100100",13432 => "10001111",13433 => "11010111",13434 => "10101100",13435 => "00001110",13436 => "11101110",13437 => "00110010",13438 => "00011000",13439 => "00110011",13440 => "00010011",13441 => "01111101",13442 => "11000000",13443 => "10110010",13444 => "11011001",13445 => "10010000",13446 => "10110001",13447 => "01011011",13448 => "10100000",13449 => "01100000",13450 => "01001001",13451 => "00000001",13452 => "11000001",13453 => "00101100",13454 => "01001010",13455 => "11100100",13456 => "00110100",13457 => "01111011",13458 => "11010011",13459 => "11001111",13460 => "00001010",13461 => "11101100",13462 => "11111011",13463 => "10101000",13464 => "11001111",13465 => "11011110",13466 => "10110111",13467 => "11110110",13468 => "11101110",13469 => "00100000",13470 => "00110011",13471 => "11111100",13472 => "11100000",13473 => "01101011",13474 => "00100000",13475 => "01000000",13476 => "01101000",13477 => "10101101",13478 => "11110110",13479 => "11001001",13480 => "01010010",13481 => "01001010",13482 => "10100010",13483 => "00101001",13484 => "10010000",13485 => "01111111",13486 => "10100010",13487 => "01110111",13488 => "11000000",13489 => "10100011",13490 => "10000001",13491 => "11110011",13492 => "01011101",13493 => "10011100",13494 => "00010001",13495 => "01100111",13496 => "11011011",13497 => "00000010",13498 => "11111101",13499 => "11101111",13500 => "10100100",13501 => "10101111",13502 => "00110110",13503 => "01010101",13504 => "01010011",13505 => "00101010",13506 => "11101100",13507 => "01000011",13508 => "10111001",13509 => "00011100",13510 => "00100100",13511 => "10011000",13512 => "01110101",13513 => "01011110",13514 => "00000100",13515 => "11111001",13516 => "10001011",13517 => "01001110",13518 => "11000110",13519 => "01111111",13520 => "10011000",13521 => "01110111",13522 => "11110101",13523 => "10011010",13524 => "10010000",13525 => "11001111",13526 => "11000011",13527 => "01110101",13528 => "10111010",13529 => "01011010",13530 => "10111000",13531 => "01101101",13532 => "01100000",13533 => "01011011",13534 => "11000001",13535 => "11110011",13536 => "11000000",13537 => "01100000",13538 => "11110101",13539 => "00110011",13540 => "11110110",13541 => "00001101",13542 => "10001010",13543 => "11100001",13544 => "01110110",13545 => "10100111",13546 => "01110101",13547 => "01111111",13548 => "11101011",13549 => "01000011",13550 => "01110100",13551 => "11100110",13552 => "01111100",13553 => "01001110",13554 => "11000000",13555 => "00101000",13556 => "00110001",13557 => "00001100",13558 => "11111110",13559 => "11100110",13560 => "11001100",13561 => "10000000",13562 => "00100000",13563 => "11111011",13564 => "01011011",13565 => "00011110",13566 => "01101010",13567 => "10100010",13568 => "01101001",13569 => "10111011",13570 => "11111110",13571 => "11111110",13572 => "10110001",13573 => "10001000",13574 => "10001101",13575 => "11001010",13576 => "10101011",13577 => "01001001",13578 => "10001110",13579 => "11100010",13580 => "01000011",13581 => "10101010",13582 => "00100100",13583 => "10000110",13584 => "00101101",13585 => "11111110",13586 => "00100101",13587 => "10110111",13588 => "11110111",13589 => "01000100",13590 => "10111001",13591 => "00011001",13592 => "10000101",13593 => "00001000",13594 => "11101001",13595 => "10000000",13596 => "11100100",13597 => "10110000",13598 => "10000010",13599 => "11001101",13600 => "10111101",13601 => "11001111",13602 => "00001010",13603 => "00110011",13604 => "11101100",13605 => "00101110",13606 => "10011101",13607 => "11001000",13608 => "01001010",13609 => "10010011",13610 => "10010101",13611 => "10011111",13612 => "01110110",13613 => "00110100",13614 => "01011100",13615 => "11111110",13616 => "01110000",13617 => "11011111",13618 => "11100000",13619 => "01011010",13620 => "10111111",13621 => "01000100",13622 => "10000000",13623 => "00011001",13624 => "00010101",13625 => "01011100",13626 => "00011000",13627 => "01100100",13628 => "01001000",13629 => "00111000",13630 => "00110001",13631 => "00101111",13632 => "01000100",13633 => "10011000",13634 => "00010111",13635 => "10010101",13636 => "00100101",13637 => "00110000",13638 => "11100111",13639 => "11111110",13640 => "01101110",13641 => "10001110",13642 => "01110100",13643 => "10010010",13644 => "11001000",13645 => "00100111",13646 => "01010111",13647 => "11100111",13648 => "10110111",13649 => "00111101",13650 => "10001101",13651 => "00101100",13652 => "00011111",13653 => "01110011",13654 => "11100011",13655 => "01011110",13656 => "01110000",13657 => "00001010",13658 => "00100100",13659 => "11101011",13660 => "10011101",13661 => "11011001",13662 => "10110100",13663 => "10111100",13664 => "11000100",13665 => "10001111",13666 => "11100010",13667 => "10100000",13668 => "11111101",13669 => "11011111",13670 => "10100000",13671 => "10000000",13672 => "10100100",13673 => "10000101",13674 => "01001110",13675 => "01011001",13676 => "00100011",13677 => "10100100",13678 => "00111010",13679 => "10011110",13680 => "01010101",13681 => "00101100",13682 => "01001111",13683 => "10111000",13684 => "00011110",13685 => "01001111",13686 => "01100001",13687 => "01101100",13688 => "01010101",13689 => "01111110",13690 => "01010011",13691 => "11111100",13692 => "11110011",13693 => "10100101",13694 => "10011101",13695 => "10011100",13696 => "01001110",13697 => "11101001",13698 => "01000111",13699 => "10001110",13700 => "11110100",13701 => "00011110",13702 => "11110111",13703 => "00100111",13704 => "11001011",13705 => "00101110",13706 => "00011100",13707 => "00001010",13708 => "00101110",13709 => "01110111",13710 => "11100001",13711 => "10110110",13712 => "10010101",13713 => "00100011",13714 => "10010110",13715 => "00100001",13716 => "01001101",13717 => "01000100",13718 => "00110001",13719 => "11101101",13720 => "11100000",13721 => "11101001",13722 => "00100110",13723 => "00110101",13724 => "11000110",13725 => "00010000",13726 => "10001001",13727 => "10111100",13728 => "01011001",13729 => "01000001",13730 => "11100111",13731 => "01101010",13732 => "11000001",13733 => "10110101",13734 => "10110110",13735 => "00000000",13736 => "00110100",13737 => "10000001",13738 => "11000111",13739 => "11100011",13740 => "00011001",13741 => "10101010",13742 => "11001100",13743 => "10001101",13744 => "01010110",13745 => "10000100",13746 => "01010010",13747 => "01011101",13748 => "01001011",13749 => "01101101",13750 => "01101010",13751 => "10101001",13752 => "11001111",13753 => "01110101",13754 => "10000010",13755 => "01010000",13756 => "01000010",13757 => "11010001",13758 => "00011010",13759 => "10000001",13760 => "00101101",13761 => "01101110",13762 => "10010110",13763 => "10011000",13764 => "01110111",13765 => "00110110",13766 => "10000010",13767 => "01101001",13768 => "01110101",13769 => "00101101",13770 => "01000111",13771 => "00101110",13772 => "10111101",13773 => "00001101",13774 => "01000001",13775 => "11101011",13776 => "11111110",13777 => "10110111",13778 => "10110001",13779 => "11011001",13780 => "00101011",13781 => "10010011",13782 => "00010011",13783 => "00001111",13784 => "11001101",13785 => "10000001",13786 => "11101010",13787 => "01100010",13788 => "01011100",13789 => "00001010",13790 => "00111010",13791 => "01000100",13792 => "01000001",13793 => "10001101",13794 => "10110000",13795 => "00100101",13796 => "01011100",13797 => "01111111",13798 => "01100000",13799 => "01011001",13800 => "11101001",13801 => "11001111",13802 => "00011001",13803 => "11010011",13804 => "01001100",13805 => "11111100",13806 => "10101011",13807 => "11010011",13808 => "10011100",13809 => "01111111",13810 => "10100100",13811 => "01000110",13812 => "01000110",13813 => "10010011",13814 => "11100011",13815 => "00010100",13816 => "00100101",13817 => "01011101",13818 => "11011001",13819 => "01110000",13820 => "10001100",13821 => "00110001",13822 => "01011101",13823 => "11000110",13824 => "10100000",13825 => "10001100",13826 => "11111100",13827 => "10010010",13828 => "01010110",13829 => "01110000",13830 => "10001001",13831 => "01100000",13832 => "01011110",13833 => "00000100",13834 => "00000011",13835 => "01111110",13836 => "01110011",13837 => "11001010",13838 => "10100110",13839 => "01010010",13840 => "01010001",13841 => "10111110",13842 => "01111110",13843 => "10101000",13844 => "01110001",13845 => "01000011",13846 => "11000011",13847 => "00101011",13848 => "10100101",13849 => "11000110",13850 => "11011011",13851 => "10111100",13852 => "10101010",13853 => "10010010",13854 => "00100010",13855 => "11010010",13856 => "01100010",13857 => "10001001",13858 => "11001101",13859 => "10100011",13860 => "01001001",13861 => "11100010",13862 => "01111100",13863 => "11001110",13864 => "00100111",13865 => "00100100",13866 => "11010101",13867 => "00110011",13868 => "11110011",13869 => "00000011",13870 => "11001001",13871 => "01100101",13872 => "01110110",13873 => "00000000",13874 => "00000000",13875 => "01011100",13876 => "10111001",13877 => "01100000",13878 => "00000111",13879 => "01000010",13880 => "11101010",13881 => "00000011",13882 => "10010000",13883 => "10001100",13884 => "01011110",13885 => "00101100",13886 => "01000001",13887 => "10101000",13888 => "11111000",13889 => "00100010",13890 => "01001111",13891 => "11101100",13892 => "11111110",13893 => "11100100",13894 => "00010010",13895 => "01111100",13896 => "00101110",13897 => "01000010",13898 => "10101011",13899 => "00000011",13900 => "11010000",13901 => "11100011",13902 => "10111101",13903 => "10111100",13904 => "01010101",13905 => "11100110",13906 => "01001100",13907 => "00011010",13908 => "11101000",13909 => "11010010",13910 => "01111000",13911 => "00110110",13912 => "10001101",13913 => "11100001",13914 => "10111111",13915 => "00110010",13916 => "10111101",13917 => "10011010",13918 => "10011010",13919 => "10011111",13920 => "00011000",13921 => "10100111",13922 => "01100000",13923 => "01110000",13924 => "10000000",13925 => "00110011",13926 => "11000110",13927 => "10100000",13928 => "00001000",13929 => "10101001",13930 => "10001100",13931 => "00111011",13932 => "10010111",13933 => "11101010",13934 => "10001000",13935 => "00101110",13936 => "10100101",13937 => "01111000",13938 => "00000001",13939 => "01011111",13940 => "10010010",13941 => "01011110",13942 => "10100100",13943 => "11000101",13944 => "01000000",13945 => "00011000",13946 => "01111000",13947 => "01110100",13948 => "01010001",13949 => "10110101",13950 => "01011011",13951 => "11111100",13952 => "00001010",13953 => "01001001",13954 => "01110101",13955 => "10110000",13956 => "10111100",13957 => "11011010",13958 => "01111001",13959 => "10011000",13960 => "10011111",13961 => "11111110",13962 => "11101001",13963 => "00001011",13964 => "01100111",13965 => "00101110",13966 => "11000011",13967 => "10010111",13968 => "01011100",13969 => "11010011",13970 => "11111000",13971 => "10111100",13972 => "01110011",13973 => "11100011",13974 => "01111000",13975 => "10001011",13976 => "01000110",13977 => "01000111",13978 => "01100001",13979 => "00000111",13980 => "10000011",13981 => "01011000",13982 => "00000100",13983 => "00111110",13984 => "01110111",13985 => "00001011",13986 => "11011101",13987 => "11101110",13988 => "01111101",13989 => "10001100",13990 => "00000111",13991 => "00001010",13992 => "11100000",13993 => "11000000",13994 => "01001011",13995 => "01101000",13996 => "01001111",13997 => "00000000",13998 => "00000100",13999 => "11110001",14000 => "10110011",14001 => "11111111",14002 => "10010000",14003 => "10001000",14004 => "01000111",14005 => "01000100",14006 => "10000001",14007 => "00110101",14008 => "00011011",14009 => "10101000",14010 => "00010110",14011 => "00011101",14012 => "01000000",14013 => "00111000",14014 => "01101000",14015 => "00101111",14016 => "10011011",14017 => "00100101",14018 => "00001011",14019 => "01011000",14020 => "10000100",14021 => "01000000",14022 => "00000100",14023 => "11111110",14024 => "00110001",14025 => "10010111",14026 => "00010001",14027 => "11110110",14028 => "10010110",14029 => "10001101",14030 => "11010011",14031 => "10010010",14032 => "00100111",14033 => "10000000",14034 => "10010001",14035 => "11011111",14036 => "10011100",14037 => "10110010",14038 => "10011110",14039 => "11001100",14040 => "11010100",14041 => "10011111",14042 => "00101010",14043 => "01110000",14044 => "00111011",14045 => "01011001",14046 => "11100001",14047 => "10111101",14048 => "10000110",14049 => "10010111",14050 => "01110001",14051 => "11011100",14052 => "01111111",14053 => "00010011",14054 => "00110010",14055 => "00110101",14056 => "01001110",14057 => "11110101",14058 => "11001111",14059 => "10001001",14060 => "01000011",14061 => "10100011",14062 => "00100110",14063 => "10111010",14064 => "01001101",14065 => "10111010",14066 => "00100000",14067 => "01010010",14068 => "11111111",14069 => "01111100",14070 => "01010011",14071 => "00111000",14072 => "00110000",14073 => "11111100",14074 => "01000001",14075 => "00000011",14076 => "01101011",14077 => "01100001",14078 => "00100001",14079 => "00101010",14080 => "10110000",14081 => "10110000",14082 => "10100111",14083 => "10011010",14084 => "10100010",14085 => "11101011",14086 => "00101111",14087 => "00001111",14088 => "11000100",14089 => "10000110",14090 => "00010010",14091 => "00001001",14092 => "11101010",14093 => "01110111",14094 => "11101100",14095 => "01011010",14096 => "11000001",14097 => "00100100",14098 => "10011111",14099 => "11001010",14100 => "11011110",14101 => "00101110",14102 => "10100010",14103 => "10001000",14104 => "11110110",14105 => "10011011",14106 => "11100100",14107 => "01111001",14108 => "10110011",14109 => "01100111",14110 => "11100001",14111 => "00101110",14112 => "10010100",14113 => "10100100",14114 => "10110101",14115 => "10001010",14116 => "00011011",14117 => "11110010",14118 => "11000010",14119 => "01011101",14120 => "11011110",14121 => "10000010",14122 => "11001111",14123 => "11011010",14124 => "01101001",14125 => "01000100",14126 => "11001000",14127 => "01000111",14128 => "00101100",14129 => "11010010",14130 => "11010011",14131 => "10100111",14132 => "00101010",14133 => "00101100",14134 => "01000000",14135 => "01000100",14136 => "01000011",14137 => "10010001",14138 => "11111001",14139 => "11100111",14140 => "11110001",14141 => "10111001",14142 => "11000110",14143 => "10110001",14144 => "10101010",14145 => "01101001",14146 => "10001100",14147 => "01110001",14148 => "00010100",14149 => "10101111",14150 => "11010011",14151 => "10011101",14152 => "11000100",14153 => "01010110",14154 => "11011100",14155 => "11101100",14156 => "11010011",14157 => "01010000",14158 => "10000110",14159 => "10111000",14160 => "11101100",14161 => "01100110",14162 => "00001110",14163 => "11111001",14164 => "10100101",14165 => "10100000",14166 => "00010010",14167 => "10001000",14168 => "00110111",14169 => "11101101",14170 => "11100000",14171 => "10000110",14172 => "10011011",14173 => "10100101",14174 => "00111110",14175 => "01111100",14176 => "00111100",14177 => "11010001",14178 => "11110001",14179 => "00000101",14180 => "11111001",14181 => "01100110",14182 => "10000111",14183 => "00101100",14184 => "11011111",14185 => "00010011",14186 => "11011100",14187 => "01100101",14188 => "00001001",14189 => "00010100",14190 => "00101100",14191 => "10010100",14192 => "01100010",14193 => "01001011",14194 => "10100110",14195 => "11110000",14196 => "11011101",14197 => "10111001",14198 => "11100111",14199 => "11000000",14200 => "10111111",14201 => "10011110",14202 => "01100001",14203 => "10110100",14204 => "11110101",14205 => "00011010",14206 => "00011100",14207 => "11000100",14208 => "01110101",14209 => "11001000",14210 => "11001011",14211 => "11010001",14212 => "10011110",14213 => "00111010",14214 => "01011100",14215 => "11000000",14216 => "00111011",14217 => "10011011",14218 => "01101100",14219 => "00001001",14220 => "00100100",14221 => "01111010",14222 => "00111110",14223 => "10101000",14224 => "01110101",14225 => "10010101",14226 => "10111111",14227 => "10100010",14228 => "00110001",14229 => "01111011",14230 => "00111110",14231 => "00100110",14232 => "01110100",14233 => "00001011",14234 => "01111000",14235 => "10000000",14236 => "00100100",14237 => "00000001",14238 => "01011001",14239 => "01111111",14240 => "11010001",14241 => "11111111",14242 => "10001000",14243 => "00110101",14244 => "10000110",14245 => "10101100",14246 => "10110011",14247 => "11010100",14248 => "01110110",14249 => "01101000",14250 => "01000010",14251 => "11101000",14252 => "01011001",14253 => "01011010",14254 => "10000110",14255 => "11111001",14256 => "00011110",14257 => "10001100",14258 => "11001100",14259 => "11111100",14260 => "11111000",14261 => "10010110",14262 => "11011010",14263 => "00011000",14264 => "01000101",14265 => "10011110",14266 => "01010101",14267 => "11110011",14268 => "01110001",14269 => "10101000",14270 => "00010101",14271 => "00001000",14272 => "00000101",14273 => "10100010",14274 => "00000100",14275 => "00010100",14276 => "01000000",14277 => "01001110",14278 => "10000100",14279 => "11000000",14280 => "11011100",14281 => "11001011",14282 => "11110001",14283 => "01100111",14284 => "01001000",14285 => "01100110",14286 => "10110000",14287 => "11011011",14288 => "10010000",14289 => "10010011",14290 => "01011101",14291 => "11100000",14292 => "01101010",14293 => "10000110",14294 => "01001100",14295 => "01111000",14296 => "10001011",14297 => "10010001",14298 => "00001011",14299 => "11000100",14300 => "11100011",14301 => "01001111",14302 => "00111101",14303 => "10110010",14304 => "10100001",14305 => "10000100",14306 => "10111011",14307 => "11010000",14308 => "00110110",14309 => "01100011",14310 => "11110111",14311 => "01101100",14312 => "01010001",14313 => "00100001",14314 => "00000101",14315 => "10001101",14316 => "01000111",14317 => "11011110",14318 => "11101110",14319 => "10000010",14320 => "01110000",14321 => "11100000",14322 => "11011100",14323 => "01101101",14324 => "10011110",14325 => "01110100",14326 => "01110001",14327 => "00100010",14328 => "00010001",14329 => "00100100",14330 => "01101011",14331 => "00000011",14332 => "01110011",14333 => "10011001",14334 => "01010000",14335 => "00011100",14336 => "10111000",14337 => "01000110",14338 => "00001110",14339 => "00110110",14340 => "10111010",14341 => "11011100",14342 => "01100111",14343 => "10101001",14344 => "00110001",14345 => "00011001",14346 => "01110000",14347 => "10100001",14348 => "01000000",14349 => "01111001",14350 => "00111011",14351 => "11101110",14352 => "01011000",14353 => "00101001",14354 => "00110001",14355 => "10101111",14356 => "10100111",14357 => "00000010",14358 => "11001111",14359 => "01011000",14360 => "00010100",14361 => "00001010",14362 => "01101011",14363 => "00000010",14364 => "01011100",14365 => "10110001",14366 => "00011101",14367 => "11100111",14368 => "01011100",14369 => "10000001",14370 => "00110011",14371 => "01101101",14372 => "01101010",14373 => "11011111",14374 => "10011110",14375 => "01001011",14376 => "01101110",14377 => "10011111",14378 => "11000000",14379 => "10000100",14380 => "01110000",14381 => "11100001",14382 => "11110101",14383 => "01110010",14384 => "00111101",14385 => "00101101",14386 => "11101011",14387 => "01011010",14388 => "01100010",14389 => "00111101",14390 => "00011011",14391 => "10110100",14392 => "01100101",14393 => "01001011",14394 => "01110110",14395 => "10000100",14396 => "00011110",14397 => "01101100",14398 => "10111000",14399 => "01000111",14400 => "11010001",14401 => "01001001",14402 => "00011101",14403 => "11010110",14404 => "11010001",14405 => "10111100",14406 => "11101110",14407 => "00010010",14408 => "11100010",14409 => "01000111",14410 => "00000000",14411 => "01001000",14412 => "01001011",14413 => "11010000",14414 => "11011011",14415 => "10001000",14416 => "00000000",14417 => "11101010",14418 => "10111101",14419 => "00001101",14420 => "11001010",14421 => "00000110",14422 => "10011100",14423 => "01011111",14424 => "11010011",14425 => "10100010",14426 => "01000101",14427 => "10110110",14428 => "01011111",14429 => "11110100",14430 => "01110001",14431 => "00111011",14432 => "11110110",14433 => "00001011",14434 => "00111010",14435 => "00010010",14436 => "10001110",14437 => "00001110",14438 => "10010101",14439 => "01101111",14440 => "01010100",14441 => "00010000",14442 => "11000010",14443 => "00111100",14444 => "11101110",14445 => "00001000",14446 => "10011111",14447 => "11000111",14448 => "00010101",14449 => "00100110",14450 => "11000100",14451 => "01001110",14452 => "10111010",14453 => "01110110",14454 => "11101001",14455 => "10100111",14456 => "10000100",14457 => "10110001",14458 => "10011111",14459 => "01001100",14460 => "01000001",14461 => "00100110",14462 => "00010010",14463 => "11110110",14464 => "10001010",14465 => "10100011",14466 => "10110010",14467 => "00001100",14468 => "00011110",14469 => "10011100",14470 => "00101010",14471 => "11100011",14472 => "01101100",14473 => "10100000",14474 => "11100011",14475 => "10110111",14476 => "10100111",14477 => "01010101",14478 => "00000101",14479 => "10011011",14480 => "11110100",14481 => "10010111",14482 => "10100001",14483 => "01011001",14484 => "00010111",14485 => "10101111",14486 => "00001010",14487 => "11000000",14488 => "00110101",14489 => "01110010",14490 => "00111001",14491 => "00010100",14492 => "11010111",14493 => "01010101",14494 => "01111000",14495 => "11110010",14496 => "10011001",14497 => "00010010",14498 => "00101010",14499 => "00111010",14500 => "10001111",14501 => "00111101",14502 => "10110100",14503 => "00011001",14504 => "01000001",14505 => "00101111",14506 => "10110010",14507 => "10111010",14508 => "11000111",14509 => "01101110",14510 => "11001000",14511 => "10111100",14512 => "10111100",14513 => "00101100",14514 => "10100010",14515 => "11011101",14516 => "10110000",14517 => "10101011",14518 => "10111101",14519 => "01111100",14520 => "10110010",14521 => "00000001",14522 => "10101111",14523 => "00001100",14524 => "01110101",14525 => "00110011",14526 => "11011111",14527 => "10111000",14528 => "10100000",14529 => "01111001",14530 => "01001101",14531 => "11100111",14532 => "10011111",14533 => "10011111",14534 => "00110111",14535 => "01111100",14536 => "10100111",14537 => "10111101",14538 => "11100000",14539 => "10100000",14540 => "00010010",14541 => "00011010",14542 => "11100101",14543 => "01001101",14544 => "00100001",14545 => "01110110",14546 => "01110111",14547 => "11110101",14548 => "11110000",14549 => "00010001",14550 => "01111000",14551 => "10101111",14552 => "11101000",14553 => "01001111",14554 => "11000110",14555 => "11101000",14556 => "01001100",14557 => "11110011",14558 => "00111011",14559 => "10000001",14560 => "11010110",14561 => "11111110",14562 => "00110111",14563 => "01011111",14564 => "00101110",14565 => "01110010",14566 => "00111101",14567 => "11101110",14568 => "01110101",14569 => "11100101",14570 => "10100011",14571 => "01011101",14572 => "00111001",14573 => "01110001",14574 => "10001010",14575 => "10000100",14576 => "00000111",14577 => "01101100",14578 => "00111000",14579 => "10111001",14580 => "01110000",14581 => "00111110",14582 => "11101110",14583 => "11100101",14584 => "00100111",14585 => "01110001",14586 => "10111001",14587 => "10001100",14588 => "11110011",14589 => "01010111",14590 => "10111000",14591 => "11011100",14592 => "11101011",14593 => "01100001",14594 => "01011011",14595 => "10101010",14596 => "11000111",14597 => "01100010",14598 => "00110111",14599 => "11111111",14600 => "10101111",14601 => "11011010",14602 => "01011001",14603 => "01111111",14604 => "00110011",14605 => "00010001",14606 => "01101100",14607 => "11010011",14608 => "00111111",14609 => "11011100",14610 => "11111110",14611 => "00011100",14612 => "01101101",14613 => "00111001",14614 => "10011001",14615 => "01001000",14616 => "01111001",14617 => "11000110",14618 => "00101100",14619 => "00100111",14620 => "10001111",14621 => "01110110",14622 => "01110010",14623 => "10110101",14624 => "00101000",14625 => "11001001",14626 => "01011001",14627 => "01000010",14628 => "01000100",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00111001" report "FAIL high bits" severity failure;
assert RAM(0) = "00100100" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
