 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "11011101",3 => "10011001",4 => "01111101",5 => "01000001",6 => "11101111",7 => "11110010",8 => "11001001",9 => "01111001",10 => "00010110",11 => "00001010",12 => "11011000",13 => "01000101",14 => "10001111",15 => "00111000",16 => "11011010",17 => "10010111",18 => "01000100",19 => "00100111",20 => "11110101",21 => "10010100",22 => "10111011",23 => "01100000",24 => "10111101",25 => "01101100",26 => "01100010",27 => "11001111",28 => "01100001",29 => "01011010",30 => "11100011",31 => "00111000",32 => "11110000",33 => "01010111",34 => "10011110",35 => "11100001",36 => "10001111",37 => "10111001",38 => "11101011",39 => "01101111",40 => "00000001",41 => "00111000",42 => "00111111",43 => "00001110",44 => "10110110",45 => "00000011",46 => "10110110",47 => "01010010",48 => "10010001",49 => "01100010",50 => "10010100",51 => "11011101",52 => "10011110",53 => "11100101",54 => "00100000",55 => "00100111",56 => "11011011",57 => "11111100",58 => "00111100",59 => "11111001",60 => "11100000",61 => "10000110",62 => "01010001",63 => "11100010",64 => "10010111",65 => "00100011",66 => "00110100",67 => "10000101",68 => "11011001",69 => "00000000",70 => "10110000",71 => "01010011",72 => "00001000",73 => "00100101",74 => "11000101",75 => "11100100",76 => "10111011",77 => "01111011",78 => "00111110",79 => "00111011",80 => "01101111",81 => "10010010",82 => "11001101",83 => "01111111",84 => "01100011",85 => "01001101",86 => "01000011",87 => "11111101",88 => "00001111",89 => "11000010",90 => "01100100",91 => "00011111",92 => "10010101",93 => "11100001",94 => "00111010",95 => "10011001",96 => "10110000",97 => "11111010",98 => "00100001",99 => "00110011",100 => "10111110",101 => "10100001",102 => "10000011",103 => "00101011",104 => "01111000",105 => "11101101",106 => "10010101",107 => "01010110",108 => "10101010",109 => "11010011",110 => "11101010",111 => "11111000",112 => "00101010",113 => "10110001",114 => "10100100",115 => "11110101",116 => "11011000",117 => "00100101",118 => "11000101",119 => "01101010",120 => "01111101",121 => "00111001",122 => "00101001",123 => "00100010",124 => "01001011",125 => "01001001",126 => "11011001",127 => "10111001",128 => "11110000",129 => "00111100",130 => "11001111",131 => "00100000",132 => "00001011",133 => "01101110",134 => "10111111",135 => "01111010",136 => "11000110",137 => "01111111",138 => "10110010",139 => "11010001",140 => "01101010",141 => "10100101",142 => "11000010",143 => "10000000",144 => "11110011",145 => "10011100",146 => "11001010",147 => "01101001",148 => "11010011",149 => "11001101",150 => "11110001",151 => "10011000",152 => "10110010",153 => "11111100",154 => "10101111",155 => "01101111",156 => "01010101",157 => "11111010",158 => "01001100",159 => "10110011",160 => "11110001",161 => "00101000",162 => "00101111",163 => "01000001",164 => "10010011",165 => "01100100",166 => "11101001",167 => "11111100",168 => "00000001",169 => "00000111",170 => "01000011",171 => "00110010",172 => "10011111",173 => "10000101",174 => "00001100",175 => "01011010",176 => "11011111",177 => "10000000",178 => "01111100",179 => "11001010",180 => "01100010",181 => "11010010",182 => "11101100",183 => "11001010",184 => "10100000",185 => "00111000",186 => "01111100",187 => "01000100",188 => "00001010",189 => "01000010",190 => "00010111",191 => "00000100",192 => "10001000",193 => "00111110",194 => "10001000",195 => "10010011",196 => "11111011",197 => "11100000",198 => "00000010",199 => "10001101",200 => "11101110",201 => "10110000",202 => "10101011",203 => "11000011",204 => "10000101",205 => "10110011",206 => "10001100",207 => "10111001",208 => "11001010",209 => "11011111",210 => "11001000",211 => "11001001",212 => "00111000",213 => "00101011",214 => "00111000",215 => "00010001",216 => "01001010",217 => "01001110",218 => "00001000",219 => "00101110",220 => "11110010",221 => "10100111",222 => "10111111",223 => "00100101",224 => "10101010",225 => "10101110",226 => "10100100",227 => "00011111",228 => "00001111",229 => "10010000",230 => "11000000",231 => "11000010",232 => "11101011",233 => "10111111",234 => "00011001",235 => "11100011",236 => "11010110",237 => "10111101",238 => "10001100",239 => "10101110",240 => "10001010",241 => "01110010",242 => "00011110",243 => "00011010",244 => "00010001",245 => "00001001",246 => "00111001",247 => "10010010",248 => "10101010",249 => "00111000",250 => "00010010",251 => "00011101",252 => "01011110",253 => "01100100",254 => "11101001",255 => "10101011",256 => "11110101",257 => "10001110",258 => "11101101",259 => "10011111",260 => "01111010",261 => "10100000",262 => "01010100",263 => "10111100",264 => "01100111",265 => "01000111",266 => "01001010",267 => "00100001",268 => "00001110",269 => "11110101",270 => "00001101",271 => "00111000",272 => "00000001",273 => "00101100",274 => "10100010",275 => "11100110",276 => "01000110",277 => "01110001",278 => "01101011",279 => "11111101",280 => "00100101",281 => "01101000",282 => "01100010",283 => "00000001",284 => "01100110",285 => "11100000",286 => "01101110",287 => "11000100",288 => "01010000",289 => "10111111",290 => "10000000",291 => "10100010",292 => "00000100",293 => "10011110",294 => "11110110",295 => "11100100",296 => "00000001",297 => "00100111",298 => "10101011",299 => "01110111",300 => "00001111",301 => "00111111",302 => "10100110",303 => "01110010",304 => "11010100",305 => "11010101",306 => "01101011",307 => "01111011",308 => "01100000",309 => "00101100",310 => "01110111",311 => "01110011",312 => "10101001",313 => "00101101",314 => "10101010",315 => "00001001",316 => "10011100",317 => "00000101",318 => "10010111",319 => "11010001",320 => "10010100",321 => "01110000",322 => "10001010",323 => "00010110",324 => "10000111",325 => "00010101",326 => "01001111",327 => "10101101",328 => "01111110",329 => "00010000",330 => "10001001",331 => "10011101",332 => "00110001",333 => "00110000",334 => "01111010",335 => "10101001",336 => "11001010",337 => "01110110",338 => "11111111",339 => "01100011",340 => "11110001",341 => "10101001",342 => "11100101",343 => "01001101",344 => "00000101",345 => "00011110",346 => "10010000",347 => "11110101",348 => "00111110",349 => "01010101",350 => "10110111",351 => "01101111",352 => "01011100",353 => "00100111",354 => "01110010",355 => "11100001",356 => "11000110",357 => "10011010",358 => "01011101",359 => "01001000",360 => "00101001",361 => "00110110",362 => "00011111",363 => "01010101",364 => "00101110",365 => "10001101",366 => "11110001",367 => "11101010",368 => "01111000",369 => "11010100",370 => "10011111",371 => "10011101",372 => "10011110",373 => "01010110",374 => "11011101",375 => "01111101",376 => "11110110",377 => "10010111",378 => "10001101",379 => "01100010",380 => "10001010",381 => "11110010",382 => "01011101",383 => "11011100",384 => "00100100",385 => "01100011",386 => "00110110",387 => "01111010",388 => "00010101",389 => "00101101",390 => "00010100",391 => "01111000",392 => "10101000",393 => "01101111",394 => "10101111",395 => "11001110",396 => "11110001",397 => "10100100",398 => "00010011",399 => "10010000",400 => "00011011",401 => "00011001",402 => "01100101",403 => "10111111",404 => "11010001",405 => "10000101",406 => "11001010",407 => "00000001",408 => "11000010",409 => "10010110",410 => "10011100",411 => "11101100",412 => "01010100",413 => "01101010",414 => "01011101",415 => "10011010",416 => "00100101",417 => "10101100",418 => "11010101",419 => "01101101",420 => "11011110",421 => "00010110",422 => "01111001",423 => "01010101",424 => "10010110",425 => "11110001",426 => "01000001",427 => "01001010",428 => "01011010",429 => "01001111",430 => "00101010",431 => "01110001",432 => "00000100",433 => "11100100",434 => "00111101",435 => "01111010",436 => "00101000",437 => "10100011",438 => "00101001",439 => "10000010",440 => "11000101",441 => "01001101",442 => "11011011",443 => "11011000",444 => "11110100",445 => "10100000",446 => "01000101",447 => "01110100",448 => "11110110",449 => "01111110",450 => "00011111",451 => "00100010",452 => "00001011",453 => "00111100",454 => "11110111",455 => "01111111",456 => "10001001",457 => "00110101",458 => "10000011",459 => "00010011",460 => "11101100",461 => "10111110",462 => "10100001",463 => "11111101",464 => "10110000",465 => "11010000",466 => "10000111",467 => "11110101",468 => "01000011",469 => "01111001",470 => "11010110",471 => "01111000",472 => "10101110",473 => "11101100",474 => "11101100",475 => "11001010",476 => "00001110",477 => "11110101",478 => "10110000",479 => "10000100",480 => "10001111",481 => "00101001",482 => "10110110",483 => "00111101",484 => "11110100",485 => "01110011",486 => "10111011",487 => "00000011",488 => "01111000",489 => "11101111",490 => "10010101",491 => "10001100",492 => "10111001",493 => "01000101",494 => "11101101",495 => "01101010",496 => "00000110",497 => "01101010",498 => "10111110",499 => "10010000",500 => "10101010",501 => "10010010",502 => "10110110",503 => "10001110",504 => "10111001",505 => "01011100",506 => "00000010",507 => "00110110",508 => "00101110",509 => "00001001",510 => "11000100",511 => "11101010",512 => "11010010",513 => "00100111",514 => "10010000",515 => "11111100",516 => "11100001",517 => "11101101",518 => "00001101",519 => "11110100",520 => "01000101",521 => "10111000",522 => "00111010",523 => "11100100",524 => "11110110",525 => "11000101",526 => "01001010",527 => "11011110",528 => "10011110",529 => "11111001",530 => "00000000",531 => "11111111",532 => "00110010",533 => "11100010",534 => "10000010",535 => "11101011",536 => "10001001",537 => "00100010",538 => "01111111",539 => "10001111",540 => "10100100",541 => "11000010",542 => "11111110",543 => "10110110",544 => "11111011",545 => "01100111",546 => "01010111",547 => "11100011",548 => "11000010",549 => "00000011",550 => "10010100",551 => "01111011",552 => "01001000",553 => "01101001",554 => "00110010",555 => "00010001",556 => "11000111",557 => "11001110",558 => "10111000",559 => "00100001",560 => "11111100",561 => "00100000",562 => "01000001",563 => "00010100",564 => "10100111",565 => "00110010",566 => "00101111",567 => "00010110",568 => "00100110",569 => "00101101",570 => "01001110",571 => "00011011",572 => "01101111",573 => "11111011",574 => "11011100",575 => "01101101",576 => "10110111",577 => "00011000",578 => "10110101",579 => "11000111",580 => "00100010",581 => "10001100",582 => "10000110",583 => "01100111",584 => "01101100",585 => "11100101",586 => "01100000",587 => "01100011",588 => "10000100",589 => "00101010",590 => "00001011",591 => "01010011",592 => "00000010",593 => "00110110",594 => "00101010",595 => "01000000",596 => "11010000",597 => "10111001",598 => "00111010",599 => "10001011",600 => "11111011",601 => "01100101",602 => "11111111",603 => "10011100",604 => "11101100",605 => "01011001",606 => "00111010",607 => "10010001",608 => "11001000",609 => "10000000",610 => "01010010",611 => "01000101",612 => "01111101",613 => "00100010",614 => "01000100",615 => "11111001",616 => "10011001",617 => "00100000",618 => "01001011",619 => "00010111",620 => "00010110",621 => "01001011",622 => "01000100",623 => "00111001",624 => "01001010",625 => "01101000",626 => "10001011",627 => "11100001",628 => "01010001",629 => "11100110",630 => "11101010",631 => "10000100",632 => "00001000",633 => "01100000",634 => "01101010",635 => "01011001",636 => "10010010",637 => "01001000",638 => "11100010",639 => "10110111",640 => "11100101",641 => "11100111",642 => "01000111",643 => "00110110",644 => "11100000",645 => "01101001",646 => "01100110",647 => "10101110",648 => "10100010",649 => "10100100",650 => "00001110",651 => "00100011",652 => "11101010",653 => "10000010",654 => "10000011",655 => "00011010",656 => "11110110",657 => "01111100",658 => "10000110",659 => "01010011",660 => "01110001",661 => "00110110",662 => "11011011",663 => "00110111",664 => "01110000",665 => "00001000",666 => "00100011",667 => "01010001",668 => "10110110",669 => "11011001",670 => "11000001",671 => "00100010",672 => "10001000",673 => "10100000",674 => "11010100",675 => "10110110",676 => "00111010",677 => "01100111",678 => "10000001",679 => "11100011",680 => "10101011",681 => "00011011",682 => "00011011",683 => "10100111",684 => "11001000",685 => "11011000",686 => "11110010",687 => "01001011",688 => "10110110",689 => "01101100",690 => "10100110",691 => "11000000",692 => "00110100",693 => "00010111",694 => "10010100",695 => "10110010",696 => "11001001",697 => "11110011",698 => "11011110",699 => "00010111",700 => "11001111",701 => "00111000",702 => "01111000",703 => "11101010",704 => "10101010",705 => "01111000",706 => "01100111",707 => "11110100",708 => "01101011",709 => "10001001",710 => "10100011",711 => "00000110",712 => "11011110",713 => "00101110",714 => "00110000",715 => "01111001",716 => "01011001",717 => "10100001",718 => "10110100",719 => "11011010",720 => "11101100",721 => "11001101",722 => "00101101",723 => "01101000",724 => "00011011",725 => "00000001",726 => "00111110",727 => "10011011",728 => "11100010",729 => "11010001",730 => "10011000",731 => "10011010",732 => "01111000",733 => "10010110",734 => "00010000",735 => "00000111",736 => "10111101",737 => "10111001",738 => "10110001",739 => "00001001",740 => "00000110",741 => "10110000",742 => "00011111",743 => "00000111",744 => "11010001",745 => "11100010",746 => "00001110",747 => "00000001",748 => "01011100",749 => "10000101",750 => "00110010",751 => "11111110",752 => "11011010",753 => "00000000",754 => "01100100",755 => "00101111",756 => "00011001",757 => "01110111",758 => "01101101",759 => "10011111",760 => "00100101",761 => "10011111",762 => "11101011",763 => "10100100",764 => "00010111",765 => "01110100",766 => "01101110",767 => "11001010",768 => "11100101",769 => "01110000",770 => "00010000",771 => "10010001",772 => "00010101",773 => "01101110",774 => "01101010",775 => "01101000",776 => "10111100",777 => "00000110",778 => "00100011",779 => "01110001",780 => "10011011",781 => "10100110",782 => "10110001",783 => "00010110",784 => "10011101",785 => "10101001",786 => "11101000",787 => "00110110",788 => "11111101",789 => "00101101",790 => "11111110",791 => "10101111",792 => "01010111",793 => "11000101",794 => "11100101",795 => "00001100",796 => "10011110",797 => "11111001",798 => "01010001",799 => "01000011",800 => "11110100",801 => "10000111",802 => "01011000",803 => "01100100",804 => "11110100",805 => "10101111",806 => "10010101",807 => "11000011",808 => "11010101",809 => "00010100",810 => "00010011",811 => "00011010",812 => "00000001",813 => "10000100",814 => "01110101",815 => "01100100",816 => "00010010",817 => "01110001",818 => "11001010",819 => "10110001",820 => "10011101",821 => "00011111",822 => "00010001",823 => "01010110",824 => "00001001",825 => "11110000",826 => "10110011",827 => "10011001",828 => "01010011",829 => "10000101",830 => "00000010",831 => "11100001",832 => "01111011",833 => "01000000",834 => "00101101",835 => "10010010",836 => "00101100",837 => "00001000",838 => "10010001",839 => "01101101",840 => "01111001",841 => "11111111",842 => "10100010",843 => "01010101",844 => "00110000",845 => "00000100",846 => "11000110",847 => "01110101",848 => "00111010",849 => "00100010",850 => "00010110",851 => "01011100",852 => "10001010",853 => "10101100",854 => "11000101",855 => "10010000",856 => "10110111",857 => "10101000",858 => "11101101",859 => "01111111",860 => "10111001",861 => "01001110",862 => "01100100",863 => "11011010",864 => "00010111",865 => "00100011",866 => "00101111",867 => "10111001",868 => "11110001",869 => "01110110",870 => "10000000",871 => "00001110",872 => "01000000",873 => "11100001",874 => "01111001",875 => "11010101",876 => "01010110",877 => "11011100",878 => "10010000",879 => "01011111",880 => "01111100",881 => "00101010",882 => "11001010",883 => "11000000",884 => "11011011",885 => "10000000",886 => "11100000",887 => "01110000",888 => "11010010",889 => "00000001",890 => "10001101",891 => "00100111",892 => "10010110",893 => "00110101",894 => "00010110",895 => "00100001",896 => "01010011",897 => "11001011",898 => "01111110",899 => "11101100",900 => "10100010",901 => "00110001",902 => "11111010",903 => "10001001",904 => "01010110",905 => "11001110",906 => "00110010",907 => "00111100",908 => "01100010",909 => "11000110",910 => "00100110",911 => "10001011",912 => "10000101",913 => "11100111",914 => "00101011",915 => "11000111",916 => "11100000",917 => "01001111",918 => "11010010",919 => "10011011",920 => "00100000",921 => "10101100",922 => "01101110",923 => "00101110",924 => "01111101",925 => "10000100",926 => "10001101",927 => "10011010",928 => "10000011",929 => "01110000",930 => "01101011",931 => "00010101",932 => "10100110",933 => "01011110",934 => "11001111",935 => "00011011",936 => "10101110",937 => "11111010",938 => "11000011",939 => "01000011",940 => "01110110",941 => "00001100",942 => "01001001",943 => "01100111",944 => "11001001",945 => "00111010",946 => "00110000",947 => "10101101",948 => "00110010",949 => "11101100",950 => "11000111",951 => "00110000",952 => "11111011",953 => "00100000",954 => "00110110",955 => "10000111",956 => "00111001",957 => "11110101",958 => "00001001",959 => "11110111",960 => "11001010",961 => "10001000",962 => "11011111",963 => "01000000",964 => "01010111",965 => "10100000",966 => "10111101",967 => "11111000",968 => "11000010",969 => "10101010",970 => "10011000",971 => "00100110",972 => "00111010",973 => "10100000",974 => "11101001",975 => "10111011",976 => "00110100",977 => "10010001",978 => "00010101",979 => "11000100",980 => "01011110",981 => "10111011",982 => "11010110",983 => "01100011",984 => "01111001",985 => "11111000",986 => "11001011",987 => "11111000",988 => "10111111",989 => "10001101",990 => "00100011",991 => "00000111",992 => "01011000",993 => "10101111",994 => "00001001",995 => "10010100",996 => "10010101",997 => "11111010",998 => "00001010",999 => "01110011",1000 => "01101010",1001 => "01010010",1002 => "01100110",1003 => "10011111",1004 => "11011111",1005 => "10111101",1006 => "10111100",1007 => "10110011",1008 => "01001111",1009 => "00100011",1010 => "11010110",1011 => "10001100",1012 => "01010100",1013 => "00011110",1014 => "10100110",1015 => "10111100",1016 => "01011000",1017 => "00100011",1018 => "11101010",1019 => "01010111",1020 => "11101111",1021 => "00010100",1022 => "11011100",1023 => "10011111",1024 => "11011101",1025 => "10111101",1026 => "01001000",1027 => "10110101",1028 => "00101110",1029 => "11001111",1030 => "11011111",1031 => "10101001",1032 => "10110111",1033 => "01010001",1034 => "11101100",1035 => "11001001",1036 => "11111001",1037 => "11011101",1038 => "01010110",1039 => "01101010",1040 => "00101000",1041 => "01101000",1042 => "10000011",1043 => "01110000",1044 => "10110011",1045 => "00110111",1046 => "11100011",1047 => "10010100",1048 => "01011101",1049 => "11010100",1050 => "00111001",1051 => "10010111",1052 => "01111101",1053 => "11011010",1054 => "00000010",1055 => "01101010",1056 => "01111100",1057 => "10100111",1058 => "01010010",1059 => "11110000",1060 => "11000001",1061 => "00011011",1062 => "10101110",1063 => "01100110",1064 => "00000101",1065 => "00111111",1066 => "11010000",1067 => "11010000",1068 => "11001111",1069 => "11011000",1070 => "00101111",1071 => "10110011",1072 => "10101000",1073 => "01000000",1074 => "01011110",1075 => "11100011",1076 => "00100011",1077 => "00111001",1078 => "11001000",1079 => "10010011",1080 => "11110110",1081 => "01010010",1082 => "10100101",1083 => "00111001",1084 => "00111111",1085 => "11001110",1086 => "00010100",1087 => "01110101",1088 => "10101110",1089 => "11001111",1090 => "01011101",1091 => "10001000",1092 => "10001111",1093 => "11111010",1094 => "01100010",1095 => "00101011",1096 => "10010000",1097 => "10111001",1098 => "10110000",1099 => "10000011",1100 => "11001111",1101 => "10101111",1102 => "01011001",1103 => "00011010",1104 => "11001101",1105 => "01100001",1106 => "11110100",1107 => "10001110",1108 => "00010111",1109 => "10110001",1110 => "01001001",1111 => "00100111",1112 => "10100101",1113 => "01010110",1114 => "10100101",1115 => "01101111",1116 => "00011100",1117 => "01011000",1118 => "01010001",1119 => "10000100",1120 => "01101000",1121 => "11111010",1122 => "11001000",1123 => "00111111",1124 => "11100100",1125 => "11111001",1126 => "11000001",1127 => "11011011",1128 => "01111011",1129 => "01011000",1130 => "01101010",1131 => "01110001",1132 => "00110010",1133 => "10100011",1134 => "11011010",1135 => "00110100",1136 => "00110010",1137 => "00010011",1138 => "00000000",1139 => "10110111",1140 => "11011010",1141 => "00111111",1142 => "01101110",1143 => "00111100",1144 => "10001001",1145 => "10010001",1146 => "01111010",1147 => "00001011",1148 => "10111011",1149 => "01010011",1150 => "01100100",1151 => "01001100",1152 => "01101011",1153 => "01110101",1154 => "10001101",1155 => "00010010",1156 => "10010000",1157 => "00000101",1158 => "01000101",1159 => "11000101",1160 => "00110100",1161 => "01001011",1162 => "11010100",1163 => "11111011",1164 => "10111111",1165 => "00110110",1166 => "11110001",1167 => "10110111",1168 => "11000001",1169 => "10101110",1170 => "01000001",1171 => "01110100",1172 => "01000010",1173 => "01000100",1174 => "00010010",1175 => "10011100",1176 => "10100101",1177 => "11001101",1178 => "01000000",1179 => "00110111",1180 => "00101010",1181 => "10110110",1182 => "10001011",1183 => "00001010",1184 => "10001010",1185 => "00101011",1186 => "11110100",1187 => "10111010",1188 => "01100101",1189 => "10001110",1190 => "01010001",1191 => "11111000",1192 => "10100100",1193 => "10001110",1194 => "11110101",1195 => "10110101",1196 => "10010011",1197 => "00111111",1198 => "01010110",1199 => "11000111",1200 => "10001111",1201 => "10111011",1202 => "01111101",1203 => "11000101",1204 => "10101010",1205 => "11001001",1206 => "01110001",1207 => "00110010",1208 => "11101000",1209 => "11111110",1210 => "00100010",1211 => "00000101",1212 => "00111101",1213 => "11000001",1214 => "10111001",1215 => "10011111",1216 => "11100111",1217 => "00000110",1218 => "11110101",1219 => "11000010",1220 => "10011101",1221 => "00000110",1222 => "01110111",1223 => "10110101",1224 => "11011001",1225 => "10100110",1226 => "00010101",1227 => "10001101",1228 => "01100010",1229 => "01100000",1230 => "10000001",1231 => "11100011",1232 => "10110111",1233 => "10011100",1234 => "01111110",1235 => "01101101",1236 => "01010100",1237 => "10101101",1238 => "11101000",1239 => "10110000",1240 => "00010110",1241 => "00000110",1242 => "00000110",1243 => "10001110",1244 => "10110101",1245 => "01100010",1246 => "00011101",1247 => "10000111",1248 => "10011110",1249 => "01111101",1250 => "00000101",1251 => "10000100",1252 => "10011110",1253 => "01110110",1254 => "01100011",1255 => "01111011",1256 => "11110100",1257 => "11111011",1258 => "01101010",1259 => "11110010",1260 => "01101100",1261 => "01111001",1262 => "00111010",1263 => "11111011",1264 => "01110010",1265 => "00010101",1266 => "10010000",1267 => "00101100",1268 => "11010101",1269 => "00110001",1270 => "00111001",1271 => "00000010",1272 => "01111000",1273 => "01011101",1274 => "01001000",1275 => "10111000",1276 => "00111100",1277 => "01000001",1278 => "11001110",1279 => "00000000",1280 => "10100100",1281 => "11101010",1282 => "01011000",1283 => "11111000",1284 => "11001111",1285 => "11000000",1286 => "11000111",1287 => "11101010",1288 => "00101011",1289 => "11010011",1290 => "00100110",1291 => "01101111",1292 => "10001100",1293 => "11011111",1294 => "11111100",1295 => "00010101",1296 => "10001000",1297 => "10011110",1298 => "01100001",1299 => "01000110",1300 => "10011110",1301 => "10000110",1302 => "00010010",1303 => "00010011",1304 => "10011001",1305 => "00100100",1306 => "11010011",1307 => "00100001",1308 => "00010100",1309 => "10010110",1310 => "10011101",1311 => "10111100",1312 => "10111101",1313 => "01000010",1314 => "11110001",1315 => "11111101",1316 => "00010001",1317 => "10110101",1318 => "00111111",1319 => "11010100",1320 => "01111111",1321 => "01010111",1322 => "01110101",1323 => "10101011",1324 => "01100001",1325 => "10110101",1326 => "00111000",1327 => "10100011",1328 => "10000110",1329 => "00010010",1330 => "10110111",1331 => "11010010",1332 => "01000010",1333 => "01011001",1334 => "10111000",1335 => "00111111",1336 => "10001001",1337 => "01100101",1338 => "10010101",1339 => "01101000",1340 => "01000010",1341 => "11000011",1342 => "01100001",1343 => "10001101",1344 => "01111101",1345 => "10011100",1346 => "01000011",1347 => "00110001",1348 => "11100100",1349 => "01101000",1350 => "11011011",1351 => "11000110",1352 => "10110000",1353 => "11001010",1354 => "01101001",1355 => "01010010",1356 => "01010111",1357 => "00100010",1358 => "01111111",1359 => "00001100",1360 => "11001111",1361 => "00111100",1362 => "01100001",1363 => "01110100",1364 => "10010000",1365 => "10000000",1366 => "10010110",1367 => "10000111",1368 => "11101101",1369 => "01111000",1370 => "00000001",1371 => "11011110",1372 => "11010010",1373 => "11011001",1374 => "00000101",1375 => "00000010",1376 => "00010111",1377 => "10001111",1378 => "00111010",1379 => "10011101",1380 => "11001010",1381 => "11001100",1382 => "01110111",1383 => "00011111",1384 => "01010101",1385 => "11011011",1386 => "11000001",1387 => "00001110",1388 => "00000100",1389 => "01110110",1390 => "00001111",1391 => "11111111",1392 => "00110101",1393 => "00101011",1394 => "00001101",1395 => "01110000",1396 => "00010011",1397 => "10110010",1398 => "01100010",1399 => "11101110",1400 => "01110110",1401 => "10001010",1402 => "10100111",1403 => "00000100",1404 => "00101001",1405 => "00000110",1406 => "10000110",1407 => "11111111",1408 => "01111111",1409 => "10100111",1410 => "10110001",1411 => "01111001",1412 => "01111000",1413 => "10010010",1414 => "01110110",1415 => "10000111",1416 => "10101011",1417 => "11011010",1418 => "01101111",1419 => "11001111",1420 => "10001010",1421 => "10001011",1422 => "01011011",1423 => "10101111",1424 => "11100011",1425 => "10001000",1426 => "01010101",1427 => "11011011",1428 => "00101110",1429 => "10110101",1430 => "00010000",1431 => "00011000",1432 => "01011100",1433 => "10111101",1434 => "11100000",1435 => "01110100",1436 => "11110010",1437 => "00000010",1438 => "01110101",1439 => "11111000",1440 => "00011110",1441 => "10010111",1442 => "01010111",1443 => "11010011",1444 => "01001111",1445 => "11001100",1446 => "10110101",1447 => "00000101",1448 => "11001110",1449 => "10110001",1450 => "01000000",1451 => "01011011",1452 => "11100010",1453 => "01010110",1454 => "11111110",1455 => "10100011",1456 => "00001111",1457 => "11100111",1458 => "01100000",1459 => "11100101",1460 => "01010011",1461 => "10100101",1462 => "11101100",1463 => "10110010",1464 => "11000110",1465 => "01101111",1466 => "00011111",1467 => "11110111",1468 => "11101011",1469 => "01111111",1470 => "11010000",1471 => "11111000",1472 => "00100111",1473 => "11010010",1474 => "00001000",1475 => "11001000",1476 => "10110100",1477 => "11100110",1478 => "11100001",1479 => "10101111",1480 => "11010000",1481 => "10001010",1482 => "11110110",1483 => "00011101",1484 => "10111111",1485 => "00010110",1486 => "00000011",1487 => "01000110",1488 => "11000100",1489 => "00001100",1490 => "10001101",1491 => "11111111",1492 => "11010101",1493 => "11010011",1494 => "00100110",1495 => "00100001",1496 => "00111110",1497 => "10110001",1498 => "01011011",1499 => "11011001",1500 => "00011101",1501 => "10001101",1502 => "00011100",1503 => "00101000",1504 => "11111010",1505 => "11101011",1506 => "11000011",1507 => "11010000",1508 => "00111011",1509 => "11010000",1510 => "10000000",1511 => "00011000",1512 => "11001011",1513 => "01100101",1514 => "00111000",1515 => "00111001",1516 => "10100100",1517 => "00001010",1518 => "01010001",1519 => "11100010",1520 => "11100101",1521 => "01010010",1522 => "00000100",1523 => "11110110",1524 => "10111011",1525 => "10001011",1526 => "01011001",1527 => "10000100",1528 => "11101110",1529 => "01111010",1530 => "10000000",1531 => "00000011",1532 => "10010100",1533 => "11011011",1534 => "10100010",1535 => "11110001",1536 => "00001001",1537 => "01010110",1538 => "11010111",1539 => "10110001",1540 => "00110101",1541 => "11100000",1542 => "01001100",1543 => "10100110",1544 => "11111010",1545 => "11000111",1546 => "11110111",1547 => "01110110",1548 => "00011100",1549 => "11011001",1550 => "01110111",1551 => "01001001",1552 => "10000101",1553 => "10010011",1554 => "00110101",1555 => "01011011",1556 => "11100001",1557 => "11111000",1558 => "10000100",1559 => "00101111",1560 => "01110010",1561 => "11111111",1562 => "01000110",1563 => "11111010",1564 => "11101000",1565 => "11011111",1566 => "11100111",1567 => "01011110",1568 => "10010101",1569 => "10110111",1570 => "01000010",1571 => "10110100",1572 => "10101011",1573 => "01000001",1574 => "01101001",1575 => "00110100",1576 => "00011100",1577 => "10010110",1578 => "00010111",1579 => "11010001",1580 => "10001101",1581 => "01000001",1582 => "10111011",1583 => "00111001",1584 => "01111010",1585 => "10100101",1586 => "01000011",1587 => "10000010",1588 => "00100011",1589 => "10111111",1590 => "10111100",1591 => "00111101",1592 => "11011010",1593 => "10101100",1594 => "11000000",1595 => "10000000",1596 => "01011110",1597 => "01001010",1598 => "01000101",1599 => "11000110",1600 => "00101111",1601 => "00000100",1602 => "01011011",1603 => "10110111",1604 => "01011011",1605 => "10011001",1606 => "10001101",1607 => "00101000",1608 => "00101000",1609 => "01001101",1610 => "00101101",1611 => "10001110",1612 => "11011010",1613 => "10100000",1614 => "11010101",1615 => "00000010",1616 => "01010111",1617 => "01110001",1618 => "11000000",1619 => "10110000",1620 => "01100001",1621 => "01101111",1622 => "10001101",1623 => "00100011",1624 => "00101110",1625 => "00000010",1626 => "11011110",1627 => "00000010",1628 => "01001011",1629 => "00110000",1630 => "10001101",1631 => "10010101",1632 => "11011110",1633 => "11100110",1634 => "01111011",1635 => "00001101",1636 => "11111101",1637 => "00111010",1638 => "01000011",1639 => "00101010",1640 => "10101110",1641 => "11101011",1642 => "00110100",1643 => "01011010",1644 => "01101010",1645 => "00100101",1646 => "01111110",1647 => "01101111",1648 => "00000101",1649 => "01001100",1650 => "10100000",1651 => "00010111",1652 => "01110101",1653 => "10110110",1654 => "10000100",1655 => "11001010",1656 => "10110010",1657 => "01001110",1658 => "11110001",1659 => "10100000",1660 => "01100100",1661 => "11101101",1662 => "11110011",1663 => "00011110",1664 => "10111111",1665 => "10100010",1666 => "01111111",1667 => "01100010",1668 => "10100001",1669 => "10011000",1670 => "10011101",1671 => "11111111",1672 => "00010011",1673 => "00001010",1674 => "00100001",1675 => "10111010",1676 => "01100101",1677 => "11011101",1678 => "00000101",1679 => "01111001",1680 => "01001000",1681 => "11001010",1682 => "11001010",1683 => "01000001",1684 => "10010111",1685 => "11111000",1686 => "10111011",1687 => "11111010",1688 => "10011001",1689 => "01000101",1690 => "10101111",1691 => "11000010",1692 => "11000110",1693 => "11101001",1694 => "00101100",1695 => "11101101",1696 => "11111110",1697 => "11100101",1698 => "11001101",1699 => "01111110",1700 => "10110101",1701 => "01101010",1702 => "11000100",1703 => "00100010",1704 => "01000011",1705 => "11001001",1706 => "01111111",1707 => "10000100",1708 => "11010111",1709 => "11100111",1710 => "11110000",1711 => "00110100",1712 => "10101111",1713 => "01111011",1714 => "00110010",1715 => "11000100",1716 => "11011001",1717 => "01000001",1718 => "11101100",1719 => "00001010",1720 => "00101111",1721 => "10111101",1722 => "10110100",1723 => "01010110",1724 => "11000001",1725 => "00010001",1726 => "00001100",1727 => "01010100",1728 => "10001010",1729 => "10111101",1730 => "01100110",1731 => "00000111",1732 => "00111000",1733 => "11000110",1734 => "01010111",1735 => "11101110",1736 => "00000110",1737 => "11001111",1738 => "10010011",1739 => "10011110",1740 => "10011000",1741 => "01001100",1742 => "00010010",1743 => "00101101",1744 => "00101101",1745 => "00100000",1746 => "01101011",1747 => "10010001",1748 => "01011000",1749 => "11010001",1750 => "00010110",1751 => "01011110",1752 => "00011011",1753 => "01110100",1754 => "00111101",1755 => "10101101",1756 => "11011011",1757 => "00101011",1758 => "11011001",1759 => "11011100",1760 => "00000110",1761 => "01000101",1762 => "00010000",1763 => "10000011",1764 => "00011000",1765 => "01001001",1766 => "10110000",1767 => "01000010",1768 => "11100101",1769 => "10101011",1770 => "11100100",1771 => "00011111",1772 => "01000011",1773 => "10101001",1774 => "01011100",1775 => "00010011",1776 => "10000011",1777 => "11101100",1778 => "10111110",1779 => "00100011",1780 => "10011000",1781 => "00000010",1782 => "00010011",1783 => "11011101",1784 => "10011010",1785 => "10001110",1786 => "11010010",1787 => "01001111",1788 => "10010010",1789 => "11111011",1790 => "01110100",1791 => "01001100",1792 => "01000111",1793 => "10100001",1794 => "01010010",1795 => "11100100",1796 => "00011101",1797 => "01100010",1798 => "10000010",1799 => "00000010",1800 => "10110001",1801 => "01000010",1802 => "10001010",1803 => "10100010",1804 => "00111101",1805 => "00011000",1806 => "01000001",1807 => "10000010",1808 => "11010101",1809 => "11111101",1810 => "00011101",1811 => "11111001",1812 => "11010110",1813 => "01010111",1814 => "00010001",1815 => "11001010",1816 => "11011010",1817 => "01101100",1818 => "01001101",1819 => "11010100",1820 => "01011111",1821 => "11100110",1822 => "00100010",1823 => "01101001",1824 => "00010011",1825 => "01101011",1826 => "01011101",1827 => "10100101",1828 => "10000111",1829 => "10000100",1830 => "10000110",1831 => "10111011",1832 => "11011000",1833 => "10111110",1834 => "11010110",1835 => "00010101",1836 => "10011010",1837 => "01001011",1838 => "11101101",1839 => "10100000",1840 => "11111110",1841 => "00000001",1842 => "10111011",1843 => "00010011",1844 => "11100100",1845 => "10011111",1846 => "10010001",1847 => "00110110",1848 => "10110000",1849 => "00111000",1850 => "11101010",1851 => "01110001",1852 => "10010011",1853 => "10001010",1854 => "10001001",1855 => "01110000",1856 => "11010001",1857 => "00011011",1858 => "00110101",1859 => "01001001",1860 => "01101110",1861 => "01100001",1862 => "01101100",1863 => "10111111",1864 => "00101001",1865 => "11100010",1866 => "00100111",1867 => "10100001",1868 => "11110001",1869 => "10001000",1870 => "11010001",1871 => "10111101",1872 => "11001101",1873 => "10111001",1874 => "00100101",1875 => "10000111",1876 => "10011000",1877 => "01110000",1878 => "01011110",1879 => "10010000",1880 => "11100000",1881 => "01101110",1882 => "00110011",1883 => "11001000",1884 => "11100011",1885 => "00000000",1886 => "11111110",1887 => "01000010",1888 => "10110000",1889 => "11100000",1890 => "00111010",1891 => "10110100",1892 => "01111001",1893 => "00001001",1894 => "01100000",1895 => "10110000",1896 => "00010001",1897 => "01110111",1898 => "01001111",1899 => "11000110",1900 => "10101000",1901 => "11000101",1902 => "00011110",1903 => "11111111",1904 => "11001110",1905 => "01100100",1906 => "10101110",1907 => "00011001",1908 => "11010100",1909 => "11101011",1910 => "10101001",1911 => "00000110",1912 => "00110100",1913 => "01000101",1914 => "00010101",1915 => "01110110",1916 => "01110101",1917 => "10100110",1918 => "00010000",1919 => "11001100",1920 => "00010101",1921 => "11011111",1922 => "00111101",1923 => "11111001",1924 => "00000110",1925 => "01101100",1926 => "00101110",1927 => "11010111",1928 => "00100110",1929 => "00000011",1930 => "01100001",1931 => "10111111",1932 => "00010000",1933 => "10111100",1934 => "10100111",1935 => "00011101",1936 => "10010100",1937 => "10001111",1938 => "11000010",1939 => "00000101",1940 => "10101100",1941 => "10100100",1942 => "10001110",1943 => "00101000",1944 => "00000000",1945 => "00111100",1946 => "01111000",1947 => "10001110",1948 => "10101100",1949 => "01001000",1950 => "10101111",1951 => "11100110",1952 => "00001011",1953 => "11110001",1954 => "00111001",1955 => "10101011",1956 => "11101000",1957 => "11000100",1958 => "01100001",1959 => "00110110",1960 => "10101010",1961 => "10000000",1962 => "00111101",1963 => "00011000",1964 => "00010101",1965 => "10110011",1966 => "11100000",1967 => "01110100",1968 => "00101100",1969 => "11100101",1970 => "01011111",1971 => "00101100",1972 => "11110001",1973 => "10110011",1974 => "01101110",1975 => "10100000",1976 => "01100110",1977 => "00001001",1978 => "10011000",1979 => "00010100",1980 => "00001001",1981 => "00001100",1982 => "10110000",1983 => "00111111",1984 => "11010110",1985 => "00010111",1986 => "10101110",1987 => "00100010",1988 => "00101101",1989 => "10010111",1990 => "11111001",1991 => "10100001",1992 => "01100101",1993 => "01110001",1994 => "00110000",1995 => "00111100",1996 => "10011110",1997 => "00010100",1998 => "01111010",1999 => "01000000",2000 => "10100000",2001 => "11111011",2002 => "01101110",2003 => "00011110",2004 => "11001011",2005 => "01010101",2006 => "11001110",2007 => "01101001",2008 => "00100101",2009 => "01100010",2010 => "00011101",2011 => "00111011",2012 => "11100100",2013 => "11100100",2014 => "01110001",2015 => "00110100",2016 => "11111110",2017 => "11101101",2018 => "11100001",2019 => "11000101",2020 => "00001110",2021 => "00010001",2022 => "00000011",2023 => "10111100",2024 => "00011100",2025 => "11010011",2026 => "01011110",2027 => "11010000",2028 => "10110011",2029 => "00000111",2030 => "01100110",2031 => "10010010",2032 => "00011000",2033 => "00101011",2034 => "01110111",2035 => "01011110",2036 => "11100111",2037 => "10010100",2038 => "00010101",2039 => "11110100",2040 => "01111000",2041 => "10000100",2042 => "11110100",2043 => "11101001",2044 => "11100000",2045 => "00100101",2046 => "00100001",2047 => "11101010",2048 => "01000101",2049 => "11111101",2050 => "00101110",2051 => "00111111",2052 => "11111100",2053 => "01101111",2054 => "00011100",2055 => "01011010",2056 => "00000100",2057 => "11110011",2058 => "10000101",2059 => "01000111",2060 => "11110010",2061 => "00000110",2062 => "11110001",2063 => "01101000",2064 => "00000101",2065 => "10111110",2066 => "01110010",2067 => "10101110",2068 => "11000101",2069 => "11100101",2070 => "10010011",2071 => "01100110",2072 => "11001110",2073 => "00000010",2074 => "10000100",2075 => "11101111",2076 => "11001101",2077 => "10001101",2078 => "00000100",2079 => "11000000",2080 => "00000110",2081 => "01110011",2082 => "10011101",2083 => "11110110",2084 => "01101000",2085 => "01000101",2086 => "01010011",2087 => "00100000",2088 => "01000101",2089 => "01101111",2090 => "00000101",2091 => "00000101",2092 => "11101100",2093 => "10101111",2094 => "00100101",2095 => "01100110",2096 => "01110001",2097 => "01110010",2098 => "10011101",2099 => "01011011",2100 => "11110101",2101 => "01011010",2102 => "01011111",2103 => "10110100",2104 => "01101011",2105 => "01011010",2106 => "11100001",2107 => "11101110",2108 => "11100110",2109 => "00111011",2110 => "00001111",2111 => "11111100",2112 => "10100010",2113 => "10010101",2114 => "11101011",2115 => "11101011",2116 => "01010100",2117 => "11001111",2118 => "01001110",2119 => "11110110",2120 => "10110110",2121 => "01000111",2122 => "11010111",2123 => "10101011",2124 => "10011001",2125 => "01110000",2126 => "01000101",2127 => "10111110",2128 => "10110101",2129 => "00010110",2130 => "10100101",2131 => "00110100",2132 => "11010010",2133 => "01001101",2134 => "00101000",2135 => "10001011",2136 => "01111111",2137 => "01101101",2138 => "00101100",2139 => "00100010",2140 => "00101111",2141 => "10110011",2142 => "10111001",2143 => "10100100",2144 => "00010011",2145 => "01101101",2146 => "11101010",2147 => "10000100",2148 => "01010101",2149 => "10000000",2150 => "11010010",2151 => "11010110",2152 => "00001100",2153 => "11011000",2154 => "10101100",2155 => "00011110",2156 => "10010100",2157 => "00100001",2158 => "01001011",2159 => "11111111",2160 => "01100111",2161 => "11010000",2162 => "00011000",2163 => "10110101",2164 => "10111111",2165 => "01000110",2166 => "11111010",2167 => "00100110",2168 => "10001101",2169 => "10100000",2170 => "00001111",2171 => "10111000",2172 => "00011010",2173 => "11001110",2174 => "00110110",2175 => "11011110",2176 => "01001110",2177 => "10100101",2178 => "01000010",2179 => "10011100",2180 => "10001111",2181 => "01110011",2182 => "10100110",2183 => "00010101",2184 => "10000010",2185 => "11000010",2186 => "01011000",2187 => "11010011",2188 => "11010010",2189 => "01001101",2190 => "11111111",2191 => "01001101",2192 => "01010010",2193 => "00110101",2194 => "00010001",2195 => "01110111",2196 => "11111111",2197 => "11100110",2198 => "11000011",2199 => "01110100",2200 => "10010101",2201 => "11011101",2202 => "00100110",2203 => "11011011",2204 => "10110010",2205 => "00110100",2206 => "01111010",2207 => "10000000",2208 => "11111110",2209 => "00100011",2210 => "01111101",2211 => "01100010",2212 => "10110110",2213 => "11001010",2214 => "10011010",2215 => "10011111",2216 => "10010000",2217 => "11100001",2218 => "00111001",2219 => "10100110",2220 => "00010000",2221 => "00001000",2222 => "01000111",2223 => "00111011",2224 => "10011011",2225 => "11001110",2226 => "01001101",2227 => "10110010",2228 => "10111111",2229 => "11001101",2230 => "00101010",2231 => "11001001",2232 => "11011111",2233 => "00101000",2234 => "11111000",2235 => "11110100",2236 => "01111101",2237 => "00110010",2238 => "11110101",2239 => "00001001",2240 => "10110000",2241 => "01111001",2242 => "01100000",2243 => "10101101",2244 => "11101101",2245 => "00011111",2246 => "01011010",2247 => "00100010",2248 => "10101100",2249 => "10001011",2250 => "01110100",2251 => "10110001",2252 => "11001000",2253 => "10110010",2254 => "01100001",2255 => "11001110",2256 => "00110110",2257 => "01110110",2258 => "00110000",2259 => "11110101",2260 => "10001000",2261 => "01100001",2262 => "01101101",2263 => "11010001",2264 => "00011110",2265 => "01110001",2266 => "00000000",2267 => "10000111",2268 => "01000100",2269 => "00011010",2270 => "01111000",2271 => "01111011",2272 => "00110100",2273 => "11001000",2274 => "11000101",2275 => "10011001",2276 => "10100101",2277 => "01100000",2278 => "01001010",2279 => "11110111",2280 => "10010110",2281 => "10101110",2282 => "01010000",2283 => "10111000",2284 => "10100100",2285 => "10111000",2286 => "00001111",2287 => "10010100",2288 => "00010010",2289 => "01100111",2290 => "11001111",2291 => "11011100",2292 => "00011011",2293 => "10011001",2294 => "00110001",2295 => "01010100",2296 => "11100001",2297 => "00001100",2298 => "10010011",2299 => "00000011",2300 => "11101010",2301 => "10010110",2302 => "10011011",2303 => "01100110",2304 => "01010010",2305 => "10000111",2306 => "10000010",2307 => "01110010",2308 => "00001100",2309 => "10110011",2310 => "01111101",2311 => "01111101",2312 => "10011110",2313 => "10011000",2314 => "00001011",2315 => "11100001",2316 => "01110010",2317 => "10010000",2318 => "11110110",2319 => "10000000",2320 => "11001010",2321 => "10111101",2322 => "01000011",2323 => "01001000",2324 => "10101111",2325 => "10010110",2326 => "01001010",2327 => "10011101",2328 => "11001000",2329 => "00011001",2330 => "11111101",2331 => "00000001",2332 => "00111001",2333 => "00101010",2334 => "00101010",2335 => "01000111",2336 => "10011010",2337 => "10111011",2338 => "11111101",2339 => "01110010",2340 => "11100101",2341 => "11101011",2342 => "00010010",2343 => "00101010",2344 => "01111100",2345 => "10000110",2346 => "00011000",2347 => "11110110",2348 => "00010111",2349 => "10001011",2350 => "00111110",2351 => "11010101",2352 => "01010101",2353 => "00110100",2354 => "10100111",2355 => "10011000",2356 => "11000111",2357 => "01010011",2358 => "01000101",2359 => "11011010",2360 => "11010000",2361 => "01101100",2362 => "11101001",2363 => "00110111",2364 => "00001100",2365 => "11110100",2366 => "10100011",2367 => "11001111",2368 => "01001100",2369 => "01011110",2370 => "10101101",2371 => "11001000",2372 => "01000110",2373 => "10000001",2374 => "10000000",2375 => "00100010",2376 => "01101101",2377 => "01111000",2378 => "00101001",2379 => "00110101",2380 => "10100101",2381 => "00010101",2382 => "01110100",2383 => "01100010",2384 => "10111111",2385 => "00011000",2386 => "11011100",2387 => "01011000",2388 => "01100100",2389 => "01001000",2390 => "00101000",2391 => "10000001",2392 => "10010100",2393 => "00100101",2394 => "11000101",2395 => "01110011",2396 => "10111000",2397 => "01100000",2398 => "11101011",2399 => "11011001",2400 => "01000011",2401 => "11110001",2402 => "10011000",2403 => "00011111",2404 => "11010100",2405 => "00111000",2406 => "11011011",2407 => "01011101",2408 => "10101011",2409 => "01010001",2410 => "00111110",2411 => "01110010",2412 => "10001001",2413 => "01110111",2414 => "10011000",2415 => "01110110",2416 => "00000101",2417 => "11100100",2418 => "11011011",2419 => "10011010",2420 => "00001000",2421 => "10000001",2422 => "10011111",2423 => "01011010",2424 => "11111001",2425 => "00001011",2426 => "10000010",2427 => "10111101",2428 => "11011101",2429 => "00011101",2430 => "11001101",2431 => "10001011",2432 => "01111100",2433 => "01010010",2434 => "01100100",2435 => "01001101",2436 => "01001110",2437 => "11101000",2438 => "11001001",2439 => "00100001",2440 => "01111100",2441 => "11101111",2442 => "11111011",2443 => "00000011",2444 => "10101101",2445 => "10100110",2446 => "11101100",2447 => "11001111",2448 => "00101100",2449 => "10010001",2450 => "01101100",2451 => "11100100",2452 => "01010111",2453 => "00001111",2454 => "01010101",2455 => "01100011",2456 => "10001100",2457 => "00100100",2458 => "11100011",2459 => "10110100",2460 => "11001000",2461 => "11101011",2462 => "00110001",2463 => "00100000",2464 => "11111110",2465 => "00110001",2466 => "11101110",2467 => "00100110",2468 => "10101001",2469 => "11011101",2470 => "11010001",2471 => "11110100",2472 => "01111100",2473 => "10010111",2474 => "00010010",2475 => "10000010",2476 => "10011110",2477 => "11001110",2478 => "01110100",2479 => "11101001",2480 => "00001000",2481 => "11000110",2482 => "00101100",2483 => "00010100",2484 => "10101001",2485 => "00011100",2486 => "00110001",2487 => "01001010",2488 => "01010111",2489 => "00011000",2490 => "01001100",2491 => "01111001",2492 => "11110110",2493 => "01101010",2494 => "01110000",2495 => "01100111",2496 => "10001111",2497 => "11101111",2498 => "01010100",2499 => "10110110",2500 => "11110111",2501 => "10010111",2502 => "00011011",2503 => "11000101",2504 => "01000000",2505 => "00000010",2506 => "10010110",2507 => "10100000",2508 => "01010101",2509 => "10101110",2510 => "10010101",2511 => "00111110",2512 => "10011011",2513 => "11010011",2514 => "10011111",2515 => "11001001",2516 => "01011000",2517 => "00000011",2518 => "00001100",2519 => "10111111",2520 => "10101100",2521 => "01101001",2522 => "01000110",2523 => "00100001",2524 => "10011000",2525 => "11001010",2526 => "10111010",2527 => "01110010",2528 => "01001010",2529 => "10111101",2530 => "01001110",2531 => "01011111",2532 => "00001110",2533 => "11100110",2534 => "00011101",2535 => "00001110",2536 => "11101110",2537 => "00000010",2538 => "00000000",2539 => "10111101",2540 => "11101000",2541 => "10011110",2542 => "01111111",2543 => "01000100",2544 => "00101001",2545 => "10001011",2546 => "00010001",2547 => "00111000",2548 => "10011100",2549 => "01001110",2550 => "10011010",2551 => "11011101",2552 => "10111010",2553 => "01001011",2554 => "00011110",2555 => "11101100",2556 => "01110110",2557 => "10011000",2558 => "10000110",2559 => "00010010",2560 => "11111111",2561 => "01000110",2562 => "11001100",2563 => "00011101",2564 => "10100110",2565 => "01101010",2566 => "10001100",2567 => "00001111",2568 => "11100001",2569 => "11010011",2570 => "10010111",2571 => "01110110",2572 => "01001010",2573 => "11110101",2574 => "10100100",2575 => "01000010",2576 => "00010110",2577 => "01111010",2578 => "10001010",2579 => "01101001",2580 => "10100100",2581 => "10001111",2582 => "11000111",2583 => "00100110",2584 => "00101001",2585 => "10001110",2586 => "00111010",2587 => "00110101",2588 => "00100011",2589 => "01110010",2590 => "01110111",2591 => "01111011",2592 => "11010111",2593 => "10111001",2594 => "10100000",2595 => "10111100",2596 => "11000111",2597 => "01010111",2598 => "01001010",2599 => "10100101",2600 => "11010001",2601 => "01000010",2602 => "01001000",2603 => "10101010",2604 => "11101100",2605 => "11001001",2606 => "10101100",2607 => "10000011",2608 => "10101100",2609 => "00000101",2610 => "01001100",2611 => "00111111",2612 => "11001101",2613 => "10011111",2614 => "10100001",2615 => "00100111",2616 => "11110110",2617 => "00001101",2618 => "10110000",2619 => "01111110",2620 => "10011100",2621 => "11001111",2622 => "11011101",2623 => "00001100",2624 => "11100000",2625 => "11110110",2626 => "01000010",2627 => "00001110",2628 => "01001010",2629 => "01000101",2630 => "10010100",2631 => "00011000",2632 => "11000100",2633 => "11100111",2634 => "00001000",2635 => "11101011",2636 => "01011101",2637 => "01111011",2638 => "11110111",2639 => "01001100",2640 => "01001111",2641 => "01000110",2642 => "10101101",2643 => "11000110",2644 => "11100001",2645 => "11011011",2646 => "01000101",2647 => "00110100",2648 => "10000100",2649 => "10110000",2650 => "01110011",2651 => "10101101",2652 => "00010110",2653 => "00110111",2654 => "10100101",2655 => "10001011",2656 => "11011010",2657 => "01011011",2658 => "11001110",2659 => "01000000",2660 => "00111100",2661 => "11111010",2662 => "11110110",2663 => "10111111",2664 => "10100000",2665 => "01100111",2666 => "11011111",2667 => "01111011",2668 => "11110000",2669 => "11011011",2670 => "00101011",2671 => "00110101",2672 => "00111111",2673 => "00100001",2674 => "01010110",2675 => "01100100",2676 => "01101001",2677 => "00111001",2678 => "01010110",2679 => "11011111",2680 => "11111100",2681 => "11110110",2682 => "10011111",2683 => "00010000",2684 => "01011110",2685 => "00100001",2686 => "01001010",2687 => "00100101",2688 => "00100010",2689 => "10101111",2690 => "00101101",2691 => "10110111",2692 => "10111000",2693 => "01010000",2694 => "01000111",2695 => "01110000",2696 => "10100101",2697 => "00111110",2698 => "01111111",2699 => "00110000",2700 => "00100110",2701 => "10111000",2702 => "00110010",2703 => "10100110",2704 => "01010011",2705 => "01101001",2706 => "01010110",2707 => "10110100",2708 => "11101011",2709 => "11011000",2710 => "00000000",2711 => "01101011",2712 => "10010101",2713 => "11101010",2714 => "01001100",2715 => "01000111",2716 => "10000101",2717 => "11111100",2718 => "01010011",2719 => "11101000",2720 => "11111111",2721 => "01000011",2722 => "00100000",2723 => "01110010",2724 => "10001000",2725 => "01001011",2726 => "11011001",2727 => "01101001",2728 => "11010101",2729 => "11010111",2730 => "01101111",2731 => "01110111",2732 => "10110011",2733 => "10101010",2734 => "11011001",2735 => "01010101",2736 => "00101000",2737 => "10010110",2738 => "10001101",2739 => "11001100",2740 => "11001011",2741 => "00110001",2742 => "01100100",2743 => "01001001",2744 => "11100000",2745 => "10111001",2746 => "11000010",2747 => "01010010",2748 => "11110100",2749 => "00100101",2750 => "00111101",2751 => "11011001",2752 => "01001010",2753 => "11111101",2754 => "01010010",2755 => "01101010",2756 => "11001001",2757 => "10011100",2758 => "11111110",2759 => "10000000",2760 => "11001100",2761 => "00111100",2762 => "00100101",2763 => "11111001",2764 => "10001001",2765 => "01111000",2766 => "10101100",2767 => "00001001",2768 => "00001100",2769 => "01010010",2770 => "00111001",2771 => "01010111",2772 => "01000110",2773 => "00111001",2774 => "10000111",2775 => "00110011",2776 => "00100011",2777 => "11101110",2778 => "00100110",2779 => "10110011",2780 => "10101100",2781 => "11011001",2782 => "00001010",2783 => "00110110",2784 => "01001001",2785 => "00010010",2786 => "11011111",2787 => "10010000",2788 => "10010110",2789 => "00101100",2790 => "01100010",2791 => "10110010",2792 => "01100001",2793 => "00001100",2794 => "11101101",2795 => "11101011",2796 => "00010011",2797 => "11010001",2798 => "10010111",2799 => "01011011",2800 => "01000101",2801 => "01110111",2802 => "01101101",2803 => "00110111",2804 => "01110010",2805 => "00100010",2806 => "11011110",2807 => "01101011",2808 => "11100100",2809 => "00001010",2810 => "10110100",2811 => "01010001",2812 => "11000000",2813 => "10010110",2814 => "01100011",2815 => "00000100",2816 => "11101110",2817 => "00110101",2818 => "10110100",2819 => "00001111",2820 => "00110011",2821 => "10010001",2822 => "01100011",2823 => "00000011",2824 => "11111000",2825 => "11010110",2826 => "10010010",2827 => "11010001",2828 => "00000000",2829 => "11010001",2830 => "11011111",2831 => "01100111",2832 => "11010001",2833 => "10110100",2834 => "00101111",2835 => "01111100",2836 => "01100010",2837 => "01000101",2838 => "11101011",2839 => "01110100",2840 => "10101101",2841 => "11010000",2842 => "10110111",2843 => "10011111",2844 => "00001100",2845 => "11011001",2846 => "11101011",2847 => "11101100",2848 => "10011101",2849 => "10100001",2850 => "01010101",2851 => "00111101",2852 => "00010101",2853 => "10101000",2854 => "10100000",2855 => "00011011",2856 => "10011110",2857 => "10111001",2858 => "01101000",2859 => "10101110",2860 => "11001010",2861 => "10101001",2862 => "01010000",2863 => "11001111",2864 => "00011010",2865 => "11111101",2866 => "10110011",2867 => "01011000",2868 => "01101011",2869 => "01111010",2870 => "10111001",2871 => "00000100",2872 => "00111000",2873 => "10011110",2874 => "11101010",2875 => "00001000",2876 => "00110000",2877 => "01101111",2878 => "11111011",2879 => "11111111",2880 => "10110100",2881 => "10010101",2882 => "11001011",2883 => "01000011",2884 => "10010101",2885 => "00010110",2886 => "11101101",2887 => "01100100",2888 => "00110000",2889 => "00000001",2890 => "11101001",2891 => "11101101",2892 => "11010101",2893 => "01000000",2894 => "01111110",2895 => "00111000",2896 => "01111100",2897 => "01010101",2898 => "01110000",2899 => "10110010",2900 => "00110111",2901 => "10010101",2902 => "11100110",2903 => "00010100",2904 => "10000011",2905 => "10011011",2906 => "10110101",2907 => "10100001",2908 => "00000010",2909 => "01000011",2910 => "00010100",2911 => "01001010",2912 => "11011010",2913 => "10111010",2914 => "11000010",2915 => "11010101",2916 => "00100011",2917 => "01110111",2918 => "01101110",2919 => "10110110",2920 => "01110111",2921 => "10001001",2922 => "11000010",2923 => "01101010",2924 => "11110100",2925 => "10011000",2926 => "10011010",2927 => "01101111",2928 => "01011100",2929 => "10011011",2930 => "01011000",2931 => "01101101",2932 => "01010111",2933 => "10100001",2934 => "11001001",2935 => "00000001",2936 => "00010110",2937 => "11001110",2938 => "00101000",2939 => "00100001",2940 => "11111010",2941 => "00100011",2942 => "11000011",2943 => "00011100",2944 => "11100100",2945 => "00100000",2946 => "01101000",2947 => "10100101",2948 => "10111011",2949 => "11100100",2950 => "00000010",2951 => "10010010",2952 => "11000000",2953 => "10010000",2954 => "10001100",2955 => "00000010",2956 => "11011100",2957 => "10011111",2958 => "10001011",2959 => "00001000",2960 => "00111000",2961 => "01100001",2962 => "11011111",2963 => "00010101",2964 => "00100110",2965 => "11101001",2966 => "01100011",2967 => "10010101",2968 => "00100100",2969 => "11101100",2970 => "01101110",2971 => "01100000",2972 => "11001111",2973 => "01111001",2974 => "01001001",2975 => "01110110",2976 => "00101101",2977 => "10100010",2978 => "11111000",2979 => "11000001",2980 => "01100111",2981 => "10010010",2982 => "01100100",2983 => "10110010",2984 => "11011110",2985 => "10110111",2986 => "11111111",2987 => "01101011",2988 => "01101110",2989 => "11010011",2990 => "11010010",2991 => "11011010",2992 => "11111110",2993 => "01111001",2994 => "10101100",2995 => "00010111",2996 => "11010001",2997 => "11010011",2998 => "11001010",2999 => "01000100",3000 => "11111110",3001 => "01000111",3002 => "10011111",3003 => "11101111",3004 => "01111010",3005 => "00001110",3006 => "01100100",3007 => "11110111",3008 => "01001000",3009 => "01110011",3010 => "11100011",3011 => "11000000",3012 => "10000111",3013 => "10000100",3014 => "00111011",3015 => "11101011",3016 => "00000011",3017 => "11111110",3018 => "11101111",3019 => "11011101",3020 => "11000101",3021 => "00100010",3022 => "01111111",3023 => "00010010",3024 => "01100001",3025 => "10110001",3026 => "11100100",3027 => "00101000",3028 => "11111111",3029 => "00100011",3030 => "10011001",3031 => "11101110",3032 => "01000001",3033 => "00111111",3034 => "01101001",3035 => "01101000",3036 => "10111000",3037 => "10000000",3038 => "11010000",3039 => "11101000",3040 => "01100010",3041 => "00011010",3042 => "01010100",3043 => "10010000",3044 => "00001111",3045 => "00101110",3046 => "01101100",3047 => "01010000",3048 => "01101110",3049 => "11110100",3050 => "11100100",3051 => "10011011",3052 => "10000100",3053 => "01011100",3054 => "01001011",3055 => "10111000",3056 => "11111010",3057 => "00111001",3058 => "00000100",3059 => "10000001",3060 => "00001011",3061 => "11011110",3062 => "10101000",3063 => "01000000",3064 => "11110110",3065 => "01101011",3066 => "00100100",3067 => "11001001",3068 => "00100100",3069 => "00100011",3070 => "00100011",3071 => "01001110",3072 => "01100010",3073 => "00010001",3074 => "11101101",3075 => "11001100",3076 => "10000010",3077 => "11000100",3078 => "11001010",3079 => "10011100",3080 => "11101000",3081 => "11100010",3082 => "11010011",3083 => "11100010",3084 => "10111110",3085 => "00111001",3086 => "11100101",3087 => "00001011",3088 => "00111111",3089 => "01111100",3090 => "11111100",3091 => "10011100",3092 => "01101111",3093 => "00111011",3094 => "00001000",3095 => "10001011",3096 => "10011011",3097 => "01100010",3098 => "10111010",3099 => "00110101",3100 => "10000010",3101 => "00001101",3102 => "00011101",3103 => "11100010",3104 => "10111011",3105 => "11101111",3106 => "01111001",3107 => "11011011",3108 => "01101111",3109 => "11110011",3110 => "00001001",3111 => "10001110",3112 => "01011000",3113 => "01110001",3114 => "00010111",3115 => "10100001",3116 => "10110001",3117 => "11001000",3118 => "01100100",3119 => "11001011",3120 => "11100011",3121 => "00110010",3122 => "11010011",3123 => "01001111",3124 => "00000101",3125 => "10100011",3126 => "10111000",3127 => "00010110",3128 => "10001011",3129 => "00110010",3130 => "01111100",3131 => "10111011",3132 => "11100010",3133 => "00101011",3134 => "10010011",3135 => "01111101",3136 => "11010011",3137 => "10001001",3138 => "11110100",3139 => "10010101",3140 => "10000110",3141 => "01110111",3142 => "01101010",3143 => "11010100",3144 => "00010111",3145 => "10100000",3146 => "01101001",3147 => "10100111",3148 => "10000000",3149 => "01000110",3150 => "11000000",3151 => "00001110",3152 => "00011100",3153 => "00000000",3154 => "11101100",3155 => "00011101",3156 => "11111100",3157 => "01100101",3158 => "10110000",3159 => "11110101",3160 => "00111000",3161 => "00000010",3162 => "00111011",3163 => "00100101",3164 => "10101101",3165 => "11001111",3166 => "11011000",3167 => "10011100",3168 => "10110010",3169 => "11001010",3170 => "01011101",3171 => "01100010",3172 => "01111101",3173 => "11110110",3174 => "11011110",3175 => "01100111",3176 => "10001000",3177 => "10010100",3178 => "11010001",3179 => "10111001",3180 => "00011000",3181 => "00111111",3182 => "11010010",3183 => "01111110",3184 => "00000000",3185 => "00001011",3186 => "11010010",3187 => "10011000",3188 => "11000111",3189 => "00101111",3190 => "01011001",3191 => "10001110",3192 => "01010000",3193 => "00011111",3194 => "11100101",3195 => "10010100",3196 => "10001100",3197 => "01100100",3198 => "10101001",3199 => "11010011",3200 => "10000111",3201 => "01011000",3202 => "01000101",3203 => "00100111",3204 => "00001010",3205 => "00010010",3206 => "10110100",3207 => "00101111",3208 => "11011011",3209 => "00111001",3210 => "01010100",3211 => "01011110",3212 => "11000101",3213 => "10000110",3214 => "01011110",3215 => "10000001",3216 => "11011110",3217 => "11010101",3218 => "01010100",3219 => "11110110",3220 => "00100001",3221 => "11100110",3222 => "10100111",3223 => "00100101",3224 => "01100011",3225 => "11111111",3226 => "00010101",3227 => "01000111",3228 => "00000100",3229 => "11110111",3230 => "11001010",3231 => "00111000",3232 => "01100110",3233 => "10111001",3234 => "11101010",3235 => "00111010",3236 => "11100100",3237 => "01110101",3238 => "11011011",3239 => "10000010",3240 => "01110110",3241 => "11001101",3242 => "11000111",3243 => "00101011",3244 => "01011001",3245 => "01100111",3246 => "00011110",3247 => "10101101",3248 => "11101110",3249 => "11110111",3250 => "00010111",3251 => "01001101",3252 => "00011000",3253 => "01100001",3254 => "00101100",3255 => "01110001",3256 => "01100111",3257 => "01011010",3258 => "11000101",3259 => "11101111",3260 => "01111110",3261 => "10110101",3262 => "10001010",3263 => "01111001",3264 => "00011111",3265 => "00111110",3266 => "00010101",3267 => "11001000",3268 => "00111011",3269 => "11010000",3270 => "01001001",3271 => "10111100",3272 => "10100001",3273 => "11001010",3274 => "10101011",3275 => "10001001",3276 => "00101111",3277 => "01111111",3278 => "10011101",3279 => "00010100",3280 => "01001011",3281 => "11100111",3282 => "11010001",3283 => "00011110",3284 => "11111100",3285 => "10001011",3286 => "00011100",3287 => "10101110",3288 => "11010111",3289 => "10000110",3290 => "00110110",3291 => "01000001",3292 => "00110110",3293 => "11001111",3294 => "00110000",3295 => "00001001",3296 => "01111100",3297 => "01011000",3298 => "10111100",3299 => "00010011",3300 => "11010110",3301 => "10010000",3302 => "10000101",3303 => "00000101",3304 => "10001101",3305 => "10010010",3306 => "10010011",3307 => "10100001",3308 => "00100100",3309 => "11000010",3310 => "00101101",3311 => "00000111",3312 => "01111000",3313 => "11100011",3314 => "01110000",3315 => "01101110",3316 => "01001110",3317 => "11110000",3318 => "01101001",3319 => "11000011",3320 => "01011000",3321 => "01111011",3322 => "01100000",3323 => "00001110",3324 => "01000001",3325 => "01011101",3326 => "11010010",3327 => "11100010",3328 => "01100010",3329 => "01010111",3330 => "01101011",3331 => "01110100",3332 => "11010000",3333 => "11110001",3334 => "00100100",3335 => "10000001",3336 => "01111110",3337 => "10110001",3338 => "10011101",3339 => "01000111",3340 => "10111001",3341 => "01111011",3342 => "01110000",3343 => "01001010",3344 => "11000110",3345 => "10101100",3346 => "00001100",3347 => "00011000",3348 => "11110100",3349 => "00100101",3350 => "11110000",3351 => "00111000",3352 => "11101110",3353 => "11111110",3354 => "00111011",3355 => "11000011",3356 => "01111000",3357 => "01001101",3358 => "10101000",3359 => "00101110",3360 => "00011111",3361 => "00110101",3362 => "10110111",3363 => "01101110",3364 => "10110001",3365 => "00100011",3366 => "10111001",3367 => "10100110",3368 => "10110001",3369 => "11100011",3370 => "11100101",3371 => "00000000",3372 => "00111101",3373 => "10101100",3374 => "00101101",3375 => "11101110",3376 => "01110111",3377 => "11101110",3378 => "10001001",3379 => "10101110",3380 => "10001110",3381 => "01011111",3382 => "10100100",3383 => "00100011",3384 => "10100101",3385 => "00010110",3386 => "10100011",3387 => "10011101",3388 => "10100011",3389 => "11100111",3390 => "00101010",3391 => "11111000",3392 => "11101000",3393 => "00111110",3394 => "11110011",3395 => "11000000",3396 => "11000011",3397 => "11001000",3398 => "01111100",3399 => "10011111",3400 => "11011010",3401 => "11100110",3402 => "00001011",3403 => "01000101",3404 => "10101001",3405 => "11101000",3406 => "11100110",3407 => "11001110",3408 => "10001001",3409 => "10111101",3410 => "01011010",3411 => "11011110",3412 => "11001100",3413 => "11110010",3414 => "10110100",3415 => "10111010",3416 => "11000011",3417 => "10110111",3418 => "01011010",3419 => "00001001",3420 => "00001000",3421 => "11000011",3422 => "00011011",3423 => "10111110",3424 => "01100111",3425 => "00001000",3426 => "11101101",3427 => "01111111",3428 => "11011000",3429 => "00111101",3430 => "11001001",3431 => "11011001",3432 => "11000000",3433 => "11010100",3434 => "10111111",3435 => "11011110",3436 => "00011011",3437 => "10111110",3438 => "10101111",3439 => "01110000",3440 => "00011001",3441 => "11000111",3442 => "11101110",3443 => "11101010",3444 => "10011000",3445 => "01101110",3446 => "00011101",3447 => "10010100",3448 => "01110010",3449 => "01011101",3450 => "10100110",3451 => "01111000",3452 => "10011100",3453 => "01001001",3454 => "01011010",3455 => "01000000",3456 => "01011011",3457 => "10100000",3458 => "01111110",3459 => "01010010",3460 => "10001100",3461 => "00011100",3462 => "01010011",3463 => "11111001",3464 => "10010000",3465 => "10110100",3466 => "10000110",3467 => "00011101",3468 => "11100110",3469 => "10111100",3470 => "10001001",3471 => "01001101",3472 => "11000101",3473 => "11000001",3474 => "11111000",3475 => "10100010",3476 => "10110101",3477 => "10001100",3478 => "00101100",3479 => "01101100",3480 => "00101100",3481 => "11011100",3482 => "00010000",3483 => "00000100",3484 => "11100000",3485 => "10111101",3486 => "01000010",3487 => "11000100",3488 => "00111000",3489 => "01010010",3490 => "10011011",3491 => "10100110",3492 => "11110110",3493 => "11001100",3494 => "11100011",3495 => "10001100",3496 => "10100001",3497 => "00011100",3498 => "10001110",3499 => "00110111",3500 => "10010101",3501 => "00100101",3502 => "11100101",3503 => "11111100",3504 => "11001100",3505 => "10100001",3506 => "11011010",3507 => "01010101",3508 => "00100100",3509 => "10001010",3510 => "11010101",3511 => "01000001",3512 => "01010111",3513 => "10101010",3514 => "00011110",3515 => "11001111",3516 => "00111001",3517 => "10101001",3518 => "00110111",3519 => "00000010",3520 => "11110111",3521 => "00011101",3522 => "11010001",3523 => "10010010",3524 => "10100100",3525 => "01110101",3526 => "00100000",3527 => "01110000",3528 => "10011100",3529 => "00101011",3530 => "01110000",3531 => "00111110",3532 => "01101110",3533 => "10101010",3534 => "10111000",3535 => "00011101",3536 => "11100011",3537 => "11111000",3538 => "01101010",3539 => "11011110",3540 => "00110110",3541 => "10011110",3542 => "10011100",3543 => "10011101",3544 => "01000000",3545 => "01010100",3546 => "00111101",3547 => "01110110",3548 => "10000011",3549 => "01001010",3550 => "11110010",3551 => "10000111",3552 => "00001111",3553 => "01000111",3554 => "01001110",3555 => "00010111",3556 => "01010110",3557 => "01101000",3558 => "11011100",3559 => "10010001",3560 => "10110011",3561 => "11011000",3562 => "01000011",3563 => "10101000",3564 => "00100100",3565 => "00111100",3566 => "00011000",3567 => "11010000",3568 => "00110101",3569 => "00111011",3570 => "01101010",3571 => "11000000",3572 => "01110011",3573 => "00001010",3574 => "10001001",3575 => "11100111",3576 => "10001111",3577 => "11011001",3578 => "10010011",3579 => "01111111",3580 => "01111101",3581 => "01010000",3582 => "01010011",3583 => "00011100",3584 => "01111011",3585 => "00101111",3586 => "01011111",3587 => "10100101",3588 => "00111000",3589 => "11001001",3590 => "10000001",3591 => "10011110",3592 => "11001010",3593 => "00100001",3594 => "01111001",3595 => "11001100",3596 => "10000011",3597 => "00100110",3598 => "11011001",3599 => "01010001",3600 => "11011010",3601 => "01111110",3602 => "01000110",3603 => "01001100",3604 => "00110000",3605 => "10110010",3606 => "00110101",3607 => "00011100",3608 => "00010000",3609 => "00100011",3610 => "00010111",3611 => "01100101",3612 => "10000001",3613 => "00111110",3614 => "01111111",3615 => "00110010",3616 => "10101101",3617 => "10010101",3618 => "10111001",3619 => "00001101",3620 => "01110100",3621 => "01001110",3622 => "10100111",3623 => "00101010",3624 => "00011001",3625 => "01101001",3626 => "11110011",3627 => "00010000",3628 => "11000000",3629 => "00110011",3630 => "11011111",3631 => "11001000",3632 => "11100000",3633 => "11101100",3634 => "01100010",3635 => "11111001",3636 => "01100111",3637 => "11011010",3638 => "10100111",3639 => "01001101",3640 => "00000100",3641 => "00101000",3642 => "11001110",3643 => "10010100",3644 => "01001001",3645 => "10101011",3646 => "01000011",3647 => "00100110",3648 => "10101110",3649 => "01101001",3650 => "00011111",3651 => "00111001",3652 => "10011011",3653 => "00010010",3654 => "01111010",3655 => "00010001",3656 => "11110111",3657 => "11100001",3658 => "00100001",3659 => "00100111",3660 => "01011001",3661 => "01101001",3662 => "00111110",3663 => "01101001",3664 => "00111110",3665 => "01001001",3666 => "00000110",3667 => "10100011",3668 => "01101101",3669 => "10101101",3670 => "10110010",3671 => "11010101",3672 => "10001000",3673 => "01000011",3674 => "00110011",3675 => "01111011",3676 => "11001111",3677 => "00011110",3678 => "10111011",3679 => "10100010",3680 => "01110101",3681 => "11101010",3682 => "11111100",3683 => "01000000",3684 => "00101001",3685 => "01100001",3686 => "00000010",3687 => "11100010",3688 => "11100011",3689 => "01100100",3690 => "11010001",3691 => "10111101",3692 => "00010011",3693 => "10111101",3694 => "10101000",3695 => "10101101",3696 => "01011011",3697 => "01111111",3698 => "01111010",3699 => "11001010",3700 => "10011000",3701 => "11010010",3702 => "01001110",3703 => "10000101",3704 => "00000010",3705 => "11111111",3706 => "10011111",3707 => "01010011",3708 => "01011011",3709 => "00001111",3710 => "10001111",3711 => "10010011",3712 => "10000101",3713 => "00111101",3714 => "10101000",3715 => "11011111",3716 => "00001010",3717 => "00001100",3718 => "10111101",3719 => "00010000",3720 => "01101101",3721 => "01000111",3722 => "01011010",3723 => "01101000",3724 => "01110100",3725 => "00100110",3726 => "00111000",3727 => "01000101",3728 => "10100001",3729 => "00101011",3730 => "10001101",3731 => "11110000",3732 => "01111111",3733 => "11110010",3734 => "11000000",3735 => "00011000",3736 => "00010110",3737 => "01100111",3738 => "11010100",3739 => "01100011",3740 => "10010100",3741 => "01010100",3742 => "00111100",3743 => "11001101",3744 => "10100110",3745 => "01110000",3746 => "10101000",3747 => "01100010",3748 => "10111110",3749 => "10011001",3750 => "11111111",3751 => "10111001",3752 => "10001010",3753 => "01111001",3754 => "01100101",3755 => "11010100",3756 => "11111000",3757 => "10011011",3758 => "10000110",3759 => "01001011",3760 => "10010000",3761 => "10110001",3762 => "01110000",3763 => "00101010",3764 => "10001001",3765 => "00011001",3766 => "00110110",3767 => "01011110",3768 => "10110001",3769 => "00001011",3770 => "01010000",3771 => "10010111",3772 => "10000001",3773 => "11111110",3774 => "11101101",3775 => "10101011",3776 => "00011010",3777 => "10110000",3778 => "10010001",3779 => "00100000",3780 => "00111000",3781 => "00000100",3782 => "10100010",3783 => "11000111",3784 => "11100100",3785 => "10000110",3786 => "10101110",3787 => "01111111",3788 => "00010011",3789 => "01111010",3790 => "10111010",3791 => "10101010",3792 => "00110100",3793 => "01101010",3794 => "00010111",3795 => "00000101",3796 => "10001101",3797 => "11000100",3798 => "11111001",3799 => "01011101",3800 => "11011010",3801 => "11001110",3802 => "00001100",3803 => "11000101",3804 => "01100111",3805 => "00000001",3806 => "00001001",3807 => "10000101",3808 => "01101011",3809 => "00110001",3810 => "01010000",3811 => "10101001",3812 => "11001011",3813 => "00000001",3814 => "01111001",3815 => "11101010",3816 => "01101010",3817 => "11001111",3818 => "11110111",3819 => "10110011",3820 => "11111011",3821 => "11110010",3822 => "10111100",3823 => "00010110",3824 => "01000111",3825 => "01010100",3826 => "10011011",3827 => "11001011",3828 => "10101001",3829 => "10001111",3830 => "11101110",3831 => "10000010",3832 => "10100000",3833 => "01000100",3834 => "01110001",3835 => "10011010",3836 => "00010101",3837 => "11100100",3838 => "01010100",3839 => "11000101",3840 => "10110100",3841 => "10011100",3842 => "01000000",3843 => "01001100",3844 => "10110011",3845 => "01011011",3846 => "01100100",3847 => "11001010",3848 => "11101011",3849 => "10001111",3850 => "01100001",3851 => "11110110",3852 => "10010001",3853 => "10010100",3854 => "01110010",3855 => "11111000",3856 => "10100100",3857 => "01011011",3858 => "00110111",3859 => "11101110",3860 => "00110111",3861 => "01000100",3862 => "11111010",3863 => "01001001",3864 => "10110100",3865 => "01011001",3866 => "11000110",3867 => "11000110",3868 => "01110101",3869 => "01010110",3870 => "10111011",3871 => "01011100",3872 => "00111110",3873 => "01001000",3874 => "10111011",3875 => "00010111",3876 => "11011011",3877 => "11001110",3878 => "00001010",3879 => "00100110",3880 => "01000100",3881 => "10000101",3882 => "11100110",3883 => "10010101",3884 => "11011010",3885 => "11101111",3886 => "11101100",3887 => "11001111",3888 => "10010101",3889 => "00011111",3890 => "10111011",3891 => "10011000",3892 => "01100101",3893 => "11010011",3894 => "10110110",3895 => "00010010",3896 => "01010010",3897 => "10111010",3898 => "01011100",3899 => "11010011",3900 => "10000111",3901 => "10111111",3902 => "11101111",3903 => "01000100",3904 => "01000100",3905 => "11100100",3906 => "01010000",3907 => "01110111",3908 => "01000011",3909 => "10111001",3910 => "11100101",3911 => "10101011",3912 => "10000011",3913 => "10101000",3914 => "10100110",3915 => "11000010",3916 => "01100101",3917 => "11111110",3918 => "00110101",3919 => "01100110",3920 => "00000110",3921 => "01110111",3922 => "01000111",3923 => "10010110",3924 => "01000001",3925 => "11001001",3926 => "01100000",3927 => "11011001",3928 => "00011001",3929 => "00000110",3930 => "01011011",3931 => "10110100",3932 => "00010011",3933 => "11010001",3934 => "00000011",3935 => "01011101",3936 => "00111010",3937 => "10111110",3938 => "10011011",3939 => "11111010",3940 => "10101010",3941 => "10101011",3942 => "01100111",3943 => "01111001",3944 => "11011011",3945 => "00100000",3946 => "11101001",3947 => "11001100",3948 => "10110101",3949 => "11100110",3950 => "00110010",3951 => "10011001",3952 => "00001000",3953 => "11100110",3954 => "00000011",3955 => "11011000",3956 => "01110111",3957 => "01110010",3958 => "00100001",3959 => "01101010",3960 => "10000110",3961 => "01101000",3962 => "10011001",3963 => "01010000",3964 => "01100001",3965 => "10010100",3966 => "01111001",3967 => "11101110",3968 => "01111010",3969 => "00001000",3970 => "11101011",3971 => "11000110",3972 => "01011010",3973 => "01010111",3974 => "01001010",3975 => "00110001",3976 => "00110010",3977 => "01011011",3978 => "11010101",3979 => "11011110",3980 => "00111011",3981 => "01110111",3982 => "01011100",3983 => "11011111",3984 => "11000001",3985 => "01010010",3986 => "11100110",3987 => "01011111",3988 => "01100011",3989 => "00010101",3990 => "00111010",3991 => "01000010",3992 => "01010010",3993 => "10010100",3994 => "01000101",3995 => "00011010",3996 => "10110111",3997 => "00111111",3998 => "01011010",3999 => "11110111",4000 => "00001010",4001 => "10100011",4002 => "11100101",4003 => "01001110",4004 => "01001011",4005 => "00010100",4006 => "01010001",4007 => "01011100",4008 => "10101010",4009 => "00010100",4010 => "01011101",4011 => "00110100",4012 => "11011111",4013 => "01001000",4014 => "00001010",4015 => "11001011",4016 => "00100110",4017 => "11001000",4018 => "01110000",4019 => "10101101",4020 => "00011001",4021 => "10110101",4022 => "10011010",4023 => "01010111",4024 => "10001101",4025 => "11010110",4026 => "00110100",4027 => "11010101",4028 => "10101101",4029 => "11011100",4030 => "10101111",4031 => "01110110",4032 => "11101010",4033 => "10001101",4034 => "01010010",4035 => "01000000",4036 => "11000111",4037 => "01010100",4038 => "10001110",4039 => "11111011",4040 => "00010100",4041 => "10011110",4042 => "11100101",4043 => "00100010",4044 => "01011000",4045 => "01011001",4046 => "00111011",4047 => "10010011",4048 => "01001110",4049 => "00110100",4050 => "11001101",4051 => "00001001",4052 => "11000011",4053 => "11100111",4054 => "10111101",4055 => "11110111",4056 => "10011101",4057 => "11001010",4058 => "11001100",4059 => "11101110",4060 => "10110110",4061 => "10000001",4062 => "00001011",4063 => "10011111",4064 => "10101001",4065 => "11110010",4066 => "11110011",4067 => "11101000",4068 => "00001010",4069 => "00101001",4070 => "00101100",4071 => "11110010",4072 => "10110010",4073 => "01000011",4074 => "00100000",4075 => "00110100",4076 => "01000000",4077 => "10001000",4078 => "00110001",4079 => "11001101",4080 => "01010010",4081 => "11011010",4082 => "10010111",4083 => "01011011",4084 => "10001100",4085 => "00011011",4086 => "00101110",4087 => "11100111",4088 => "11000010",4089 => "11100001",4090 => "01111011",4091 => "10101011",4092 => "00010011",4093 => "00100100",4094 => "01011110",4095 => "01011111",4096 => "01010110",4097 => "11111010",4098 => "01011001",4099 => "10001000",4100 => "00111001",4101 => "11100100",4102 => "01000111",4103 => "01011001",4104 => "10000001",4105 => "01001101",4106 => "00001100",4107 => "01101101",4108 => "10100001",4109 => "10101011",4110 => "11100100",4111 => "01110100",4112 => "01111000",4113 => "10000110",4114 => "11101001",4115 => "00111011",4116 => "01001011",4117 => "11100101",4118 => "00010000",4119 => "00100110",4120 => "10100010",4121 => "11101001",4122 => "10010111",4123 => "11001011",4124 => "01010110",4125 => "00011010",4126 => "01101010",4127 => "11100100",4128 => "11000001",4129 => "01101101",4130 => "00101101",4131 => "01101110",4132 => "00110110",4133 => "10011010",4134 => "10000100",4135 => "10111010",4136 => "10000010",4137 => "01111000",4138 => "10011010",4139 => "11011001",4140 => "01001110",4141 => "00011110",4142 => "11010000",4143 => "10001111",4144 => "11111010",4145 => "01101101",4146 => "00001001",4147 => "00010010",4148 => "10011010",4149 => "11010111",4150 => "11110011",4151 => "11101100",4152 => "00100011",4153 => "00010101",4154 => "00111001",4155 => "10111001",4156 => "00111010",4157 => "01010011",4158 => "01011111",4159 => "00011010",4160 => "00000011",4161 => "11011010",4162 => "10100010",4163 => "01101000",4164 => "01110111",4165 => "11110110",4166 => "00100011",4167 => "11001010",4168 => "10001110",4169 => "01001011",4170 => "01000001",4171 => "00111010",4172 => "10111000",4173 => "01011000",4174 => "11100111",4175 => "00001001",4176 => "01101110",4177 => "11111110",4178 => "10011010",4179 => "11100110",4180 => "00010111",4181 => "01011101",4182 => "00101000",4183 => "01110011",4184 => "00000011",4185 => "01111110",4186 => "11010001",4187 => "00001011",4188 => "11100011",4189 => "01110110",4190 => "01010111",4191 => "10110101",4192 => "00011000",4193 => "01001000",4194 => "00001111",4195 => "00011101",4196 => "11101100",4197 => "11110100",4198 => "00011010",4199 => "10000001",4200 => "10011011",4201 => "00010001",4202 => "10110000",4203 => "00011001",4204 => "11100010",4205 => "11011110",4206 => "01010101",4207 => "00001011",4208 => "00011111",4209 => "10101011",4210 => "00111101",4211 => "10101111",4212 => "01110001",4213 => "10101011",4214 => "10011100",4215 => "00011011",4216 => "01101100",4217 => "01110000",4218 => "00111000",4219 => "11111010",4220 => "00010110",4221 => "00111111",4222 => "10001110",4223 => "00111001",4224 => "11001110",4225 => "11101100",4226 => "11001000",4227 => "10101101",4228 => "01111101",4229 => "11110110",4230 => "11101011",4231 => "10111001",4232 => "00011111",4233 => "00101011",4234 => "10111110",4235 => "11110000",4236 => "00001010",4237 => "10001101",4238 => "11010011",4239 => "11101111",4240 => "11001110",4241 => "00001010",4242 => "11101001",4243 => "11011001",4244 => "00100011",4245 => "00010011",4246 => "10001110",4247 => "11111011",4248 => "11111010",4249 => "10011111",4250 => "10100000",4251 => "01011111",4252 => "00101011",4253 => "01111110",4254 => "10010000",4255 => "11100111",4256 => "10011111",4257 => "10010000",4258 => "10100110",4259 => "11001111",4260 => "00101101",4261 => "00110101",4262 => "10111000",4263 => "00101001",4264 => "01100011",4265 => "11101000",4266 => "00001011",4267 => "00010100",4268 => "11000010",4269 => "01110111",4270 => "01110101",4271 => "11000101",4272 => "10101001",4273 => "01011100",4274 => "00111100",4275 => "10001100",4276 => "11010110",4277 => "10101000",4278 => "11011100",4279 => "00111001",4280 => "10010011",4281 => "10000111",4282 => "11110100",4283 => "00000001",4284 => "11011000",4285 => "00001000",4286 => "11011100",4287 => "01100011",4288 => "11011010",4289 => "11011001",4290 => "01100000",4291 => "01000010",4292 => "10111001",4293 => "01110100",4294 => "11010011",4295 => "00111100",4296 => "01100000",4297 => "11011110",4298 => "11111111",4299 => "11001000",4300 => "11000011",4301 => "00101101",4302 => "10110100",4303 => "00001010",4304 => "01101011",4305 => "00000101",4306 => "11011001",4307 => "10011110",4308 => "01010110",4309 => "00100110",4310 => "10111100",4311 => "11011110",4312 => "00110001",4313 => "10110010",4314 => "11111100",4315 => "01110000",4316 => "00100110",4317 => "11111101",4318 => "10010110",4319 => "00100001",4320 => "11011101",4321 => "10000010",4322 => "00101101",4323 => "00111011",4324 => "00100101",4325 => "10011110",4326 => "10000100",4327 => "10000110",4328 => "10010000",4329 => "10001010",4330 => "01111110",4331 => "00101111",4332 => "11001011",4333 => "10110101",4334 => "10011110",4335 => "11111011",4336 => "00000110",4337 => "10111100",4338 => "00001101",4339 => "11100100",4340 => "01111000",4341 => "11011001",4342 => "00011000",4343 => "11001100",4344 => "01101101",4345 => "00010010",4346 => "00001011",4347 => "00011011",4348 => "00000010",4349 => "01100000",4350 => "10011101",4351 => "10100010",4352 => "00101100",4353 => "10111101",4354 => "00010000",4355 => "01100110",4356 => "01001011",4357 => "11100001",4358 => "10110000",4359 => "01100101",4360 => "10101000",4361 => "00100111",4362 => "00000000",4363 => "00100010",4364 => "11011111",4365 => "10101110",4366 => "00100000",4367 => "11010101",4368 => "01110110",4369 => "00011110",4370 => "11001010",4371 => "00101100",4372 => "11000001",4373 => "11011010",4374 => "00010010",4375 => "11111011",4376 => "00110000",4377 => "10110001",4378 => "00011000",4379 => "00010101",4380 => "11001101",4381 => "00011110",4382 => "10001101",4383 => "01101101",4384 => "01101110",4385 => "00100110",4386 => "10100100",4387 => "01011001",4388 => "10011110",4389 => "11011101",4390 => "10100001",4391 => "10111001",4392 => "11111110",4393 => "00110111",4394 => "11111101",4395 => "10011000",4396 => "01011100",4397 => "01010111",4398 => "01111010",4399 => "01011101",4400 => "00110010",4401 => "01101010",4402 => "10110111",4403 => "11011101",4404 => "00010110",4405 => "01011000",4406 => "00110110",4407 => "11110101",4408 => "01111000",4409 => "01101100",4410 => "00100110",4411 => "01000101",4412 => "10110010",4413 => "01100111",4414 => "10100101",4415 => "01011111",4416 => "11001011",4417 => "00100110",4418 => "01011001",4419 => "00000110",4420 => "10110001",4421 => "10011001",4422 => "10100010",4423 => "11010010",4424 => "01101011",4425 => "01111000",4426 => "10100110",4427 => "00000011",4428 => "10001000",4429 => "11010011",4430 => "00000111",4431 => "01110101",4432 => "01011100",4433 => "10101100",4434 => "10100000",4435 => "00010111",4436 => "00100010",4437 => "10110101",4438 => "11101011",4439 => "10110000",4440 => "00110110",4441 => "11000111",4442 => "10101111",4443 => "01110000",4444 => "10100010",4445 => "10001100",4446 => "00011101",4447 => "10110010",4448 => "00011111",4449 => "00010111",4450 => "10001110",4451 => "01001101",4452 => "01100101",4453 => "10110111",4454 => "11101001",4455 => "00101100",4456 => "10010110",4457 => "00000001",4458 => "01001100",4459 => "11000100",4460 => "10010010",4461 => "11111101",4462 => "00100111",4463 => "00011101",4464 => "01000101",4465 => "00001011",4466 => "00000010",4467 => "10100001",4468 => "01101111",4469 => "01111101",4470 => "11000111",4471 => "10010001",4472 => "11101111",4473 => "10101100",4474 => "01111010",4475 => "00010001",4476 => "01010111",4477 => "00111111",4478 => "11011011",4479 => "01001111",4480 => "10011110",4481 => "10100110",4482 => "11100101",4483 => "11010100",4484 => "01100111",4485 => "10000110",4486 => "01101001",4487 => "00000000",4488 => "01100011",4489 => "11110101",4490 => "10100000",4491 => "00111110",4492 => "01011001",4493 => "01010000",4494 => "10000110",4495 => "10011000",4496 => "00110100",4497 => "11100011",4498 => "00101101",4499 => "10110010",4500 => "10110001",4501 => "00011101",4502 => "01101011",4503 => "01011101",4504 => "10100011",4505 => "01000100",4506 => "11111011",4507 => "11101011",4508 => "10011001",4509 => "11100001",4510 => "11110011",4511 => "01100100",4512 => "01110010",4513 => "00111101",4514 => "00001010",4515 => "10000010",4516 => "11110100",4517 => "00111101",4518 => "11100010",4519 => "00110100",4520 => "00011011",4521 => "11110100",4522 => "00101001",4523 => "00100010",4524 => "10100101",4525 => "11001100",4526 => "01110111",4527 => "10000100",4528 => "01000111",4529 => "11010001",4530 => "10101100",4531 => "10010100",4532 => "01010000",4533 => "01011111",4534 => "11001110",4535 => "10000100",4536 => "01101110",4537 => "00011010",4538 => "01000100",4539 => "01000101",4540 => "01011000",4541 => "00100000",4542 => "11110010",4543 => "00010111",4544 => "10001100",4545 => "10101000",4546 => "01000000",4547 => "00111110",4548 => "01010011",4549 => "10000111",4550 => "10001101",4551 => "00101000",4552 => "00010011",4553 => "11000110",4554 => "11101100",4555 => "00000111",4556 => "01100001",4557 => "01001000",4558 => "11000101",4559 => "01001111",4560 => "00110101",4561 => "00001010",4562 => "01111001",4563 => "10000110",4564 => "01011001",4565 => "11000011",4566 => "11101101",4567 => "10000001",4568 => "10011100",4569 => "11111011",4570 => "01110000",4571 => "01101110",4572 => "01011001",4573 => "01000000",4574 => "11001000",4575 => "01000000",4576 => "00101001",4577 => "10100010",4578 => "10110111",4579 => "11111111",4580 => "00000101",4581 => "01011110",4582 => "00010010",4583 => "00110010",4584 => "10100010",4585 => "11111000",4586 => "11100101",4587 => "10110010",4588 => "11000010",4589 => "10100111",4590 => "00011111",4591 => "10111011",4592 => "01011101",4593 => "11101001",4594 => "10000100",4595 => "11101100",4596 => "11111000",4597 => "00010100",4598 => "01101100",4599 => "11110101",4600 => "11001110",4601 => "01001011",4602 => "00101000",4603 => "10100001",4604 => "11111010",4605 => "10011111",4606 => "10000101",4607 => "10111001",4608 => "10000010",4609 => "11101011",4610 => "00100001",4611 => "01101001",4612 => "01111110",4613 => "01010101",4614 => "01100100",4615 => "11011101",4616 => "00101110",4617 => "11110111",4618 => "10000000",4619 => "11001010",4620 => "11101011",4621 => "00110101",4622 => "01101101",4623 => "10010110",4624 => "01110111",4625 => "10010110",4626 => "10011100",4627 => "11010010",4628 => "10111100",4629 => "00011000",4630 => "00100100",4631 => "11101110",4632 => "11010110",4633 => "11011111",4634 => "10001110",4635 => "00000011",4636 => "11001101",4637 => "00100011",4638 => "01000011",4639 => "11010001",4640 => "00001001",4641 => "00000001",4642 => "10110111",4643 => "11010001",4644 => "00100100",4645 => "01010111",4646 => "11101101",4647 => "11100000",4648 => "11110110",4649 => "10100101",4650 => "01110000",4651 => "01001001",4652 => "10000100",4653 => "10000111",4654 => "10100000",4655 => "00000000",4656 => "10000001",4657 => "10100000",4658 => "10010110",4659 => "11010010",4660 => "01010010",4661 => "00001100",4662 => "11100001",4663 => "10001000",4664 => "10110110",4665 => "01111100",4666 => "11010100",4667 => "01101110",4668 => "01011010",4669 => "11110000",4670 => "10111000",4671 => "00110101",4672 => "00001100",4673 => "10001000",4674 => "11100011",4675 => "01011110",4676 => "00010101",4677 => "10000111",4678 => "00010110",4679 => "10110111",4680 => "10110001",4681 => "01111110",4682 => "00100100",4683 => "00011111",4684 => "00001001",4685 => "00011000",4686 => "00001101",4687 => "00111011",4688 => "01000011",4689 => "11010100",4690 => "01101001",4691 => "10011011",4692 => "01001110",4693 => "01100100",4694 => "00110110",4695 => "01011111",4696 => "10100100",4697 => "10111010",4698 => "00101000",4699 => "01001001",4700 => "11101101",4701 => "10011110",4702 => "01100111",4703 => "00011110",4704 => "10010110",4705 => "01101001",4706 => "01001011",4707 => "11010011",4708 => "10000101",4709 => "11101101",4710 => "11100100",4711 => "10010001",4712 => "00101101",4713 => "11110101",4714 => "00010110",4715 => "01001111",4716 => "00110011",4717 => "11011111",4718 => "00010110",4719 => "10111011",4720 => "11000110",4721 => "01010100",4722 => "01110111",4723 => "10111011",4724 => "11111010",4725 => "01001111",4726 => "00011010",4727 => "00000011",4728 => "01010010",4729 => "11001001",4730 => "10100110",4731 => "01010101",4732 => "00111101",4733 => "01010001",4734 => "11110010",4735 => "00011001",4736 => "11100100",4737 => "01111111",4738 => "00111001",4739 => "01011111",4740 => "10010100",4741 => "01011110",4742 => "00100111",4743 => "01000011",4744 => "01111100",4745 => "10110101",4746 => "11111010",4747 => "11111110",4748 => "01000001",4749 => "11111010",4750 => "11010110",4751 => "11101111",4752 => "10000110",4753 => "10010000",4754 => "00000001",4755 => "11100111",4756 => "00000010",4757 => "00101110",4758 => "11101011",4759 => "10110110",4760 => "01111101",4761 => "01000101",4762 => "11100011",4763 => "01110111",4764 => "10011011",4765 => "10001000",4766 => "11101101",4767 => "00101001",4768 => "01010000",4769 => "01011111",4770 => "10011100",4771 => "00011001",4772 => "10010010",4773 => "11100001",4774 => "10110010",4775 => "11011100",4776 => "11110111",4777 => "11111011",4778 => "00010011",4779 => "11111000",4780 => "00000110",4781 => "11111010",4782 => "11111001",4783 => "01101100",4784 => "11110010",4785 => "11101001",4786 => "10011000",4787 => "10100110",4788 => "00000101",4789 => "11011101",4790 => "11111011",4791 => "00010110",4792 => "00110011",4793 => "10100110",4794 => "11111001",4795 => "01011000",4796 => "10001000",4797 => "11011001",4798 => "01100111",4799 => "00001001",4800 => "00100100",4801 => "01010011",4802 => "00011001",4803 => "10111001",4804 => "01001100",4805 => "11001010",4806 => "11110011",4807 => "11100100",4808 => "01110110",4809 => "11011100",4810 => "10101011",4811 => "00000110",4812 => "11101011",4813 => "11001110",4814 => "00011111",4815 => "11110000",4816 => "01101101",4817 => "11000001",4818 => "11010100",4819 => "10111010",4820 => "11100010",4821 => "00111011",4822 => "11001001",4823 => "10100110",4824 => "11100100",4825 => "00110100",4826 => "00111010",4827 => "00101001",4828 => "10001000",4829 => "10111011",4830 => "01001010",4831 => "00111010",4832 => "01011111",4833 => "00010000",4834 => "01001001",4835 => "01010011",4836 => "00000110",4837 => "01111100",4838 => "00110010",4839 => "00000111",4840 => "11110001",4841 => "10000000",4842 => "11011100",4843 => "01111001",4844 => "11110110",4845 => "11000000",4846 => "01000111",4847 => "11111011",4848 => "10011000",4849 => "01110000",4850 => "11110010",4851 => "00001010",4852 => "11011101",4853 => "00110011",4854 => "10100100",4855 => "01011111",4856 => "01010100",4857 => "11101000",4858 => "01100000",4859 => "10000110",4860 => "10001000",4861 => "10110000",4862 => "00101001",4863 => "00101100",4864 => "11000111",4865 => "00011110",4866 => "01000010",4867 => "00001000",4868 => "11000111",4869 => "01001000",4870 => "00111110",4871 => "11111111",4872 => "01110001",4873 => "10111110",4874 => "00101101",4875 => "01000111",4876 => "11101001",4877 => "00010100",4878 => "01011110",4879 => "11000000",4880 => "01111001",4881 => "10111011",4882 => "01011010",4883 => "10100000",4884 => "11110110",4885 => "01110101",4886 => "01011101",4887 => "01110110",4888 => "00011011",4889 => "01101110",4890 => "00100010",4891 => "00011001",4892 => "11001010",4893 => "01011110",4894 => "10001011",4895 => "01011001",4896 => "00101000",4897 => "00010000",4898 => "01110000",4899 => "11011100",4900 => "11000000",4901 => "01111100",4902 => "11000000",4903 => "10000011",4904 => "00100111",4905 => "00010010",4906 => "10100001",4907 => "11111000",4908 => "01000010",4909 => "10101110",4910 => "11100110",4911 => "00011101",4912 => "00011000",4913 => "00010111",4914 => "10011101",4915 => "10000010",4916 => "11001110",4917 => "00000111",4918 => "10101000",4919 => "01100100",4920 => "11011100",4921 => "10100001",4922 => "10000110",4923 => "00111100",4924 => "01111101",4925 => "00111111",4926 => "00100001",4927 => "11101011",4928 => "11101111",4929 => "00000100",4930 => "00000100",4931 => "11000111",4932 => "00111101",4933 => "11011101",4934 => "00100001",4935 => "11101111",4936 => "11011000",4937 => "10001001",4938 => "00000001",4939 => "01110110",4940 => "00001001",4941 => "01001100",4942 => "10100011",4943 => "01000100",4944 => "11111001",4945 => "01110111",4946 => "00101100",4947 => "00001100",4948 => "10100000",4949 => "01010101",4950 => "10000001",4951 => "00101101",4952 => "11111010",4953 => "00011100",4954 => "10000100",4955 => "01000111",4956 => "01010001",4957 => "01101011",4958 => "11000011",4959 => "01111000",4960 => "11011101",4961 => "10000010",4962 => "01100101",4963 => "00010010",4964 => "01001001",4965 => "11011110",4966 => "11011101",4967 => "00001010",4968 => "10111001",4969 => "01111010",4970 => "01001010",4971 => "00001011",4972 => "00001111",4973 => "11110101",4974 => "11110110",4975 => "10101000",4976 => "00000110",4977 => "11111101",4978 => "00100000",4979 => "11100111",4980 => "11110110",4981 => "01100011",4982 => "00000110",4983 => "00101110",4984 => "11011111",4985 => "00111010",4986 => "10111100",4987 => "00101000",4988 => "01000001",4989 => "00011101",4990 => "01100010",4991 => "10110110",4992 => "11110100",4993 => "10111011",4994 => "00011111",4995 => "11001111",4996 => "01111011",4997 => "01100111",4998 => "00101110",4999 => "00100111",5000 => "00100111",5001 => "01100110",5002 => "00011110",5003 => "10011000",5004 => "00100010",5005 => "10010001",5006 => "11010001",5007 => "11101110",5008 => "10100101",5009 => "01101001",5010 => "00010111",5011 => "10101100",5012 => "00011000",5013 => "01111000",5014 => "01001110",5015 => "10010111",5016 => "10000010",5017 => "00100000",5018 => "01011010",5019 => "01101111",5020 => "00100100",5021 => "00010100",5022 => "00001111",5023 => "10110101",5024 => "10100110",5025 => "10000101",5026 => "11000100",5027 => "00010110",5028 => "00011111",5029 => "11010100",5030 => "10000000",5031 => "01011010",5032 => "01110010",5033 => "00110110",5034 => "01011011",5035 => "10010011",5036 => "10010100",5037 => "01101011",5038 => "01101111",5039 => "01010100",5040 => "11001101",5041 => "11011000",5042 => "10010111",5043 => "10111010",5044 => "10010111",5045 => "00111010",5046 => "11001111",5047 => "10011111",5048 => "01100101",5049 => "11000111",5050 => "10010001",5051 => "00001110",5052 => "00010001",5053 => "10000011",5054 => "10100010",5055 => "11100101",5056 => "11110001",5057 => "11000110",5058 => "10001010",5059 => "00100110",5060 => "01110110",5061 => "10110001",5062 => "11010110",5063 => "01100001",5064 => "11000011",5065 => "10001010",5066 => "10110100",5067 => "11011011",5068 => "11100100",5069 => "10111110",5070 => "01111000",5071 => "00000011",5072 => "00000000",5073 => "10000001",5074 => "11011101",5075 => "10011111",5076 => "11010011",5077 => "00010000",5078 => "00010010",5079 => "10010110",5080 => "11111010",5081 => "01110111",5082 => "01000110",5083 => "10111100",5084 => "01001111",5085 => "00011101",5086 => "10100100",5087 => "01101101",5088 => "10011110",5089 => "10000001",5090 => "11100010",5091 => "10100000",5092 => "00001001",5093 => "11111100",5094 => "10011001",5095 => "01001111",5096 => "11001100",5097 => "01101000",5098 => "11101011",5099 => "01110110",5100 => "00001010",5101 => "01010111",5102 => "10110011",5103 => "01001110",5104 => "11101001",5105 => "00101000",5106 => "10110110",5107 => "01100111",5108 => "11000111",5109 => "10011111",5110 => "01101001",5111 => "00000000",5112 => "11100010",5113 => "01000001",5114 => "11100001",5115 => "00001100",5116 => "01101000",5117 => "10101010",5118 => "11101000",5119 => "11101111",5120 => "10000011",5121 => "00111100",5122 => "11110100",5123 => "11110001",5124 => "01000101",5125 => "11100100",5126 => "00001000",5127 => "11010010",5128 => "01100101",5129 => "01110001",5130 => "10111001",5131 => "00001110",5132 => "01000000",5133 => "00100100",5134 => "00110011",5135 => "11001010",5136 => "11001110",5137 => "10010101",5138 => "00010100",5139 => "00011011",5140 => "00011100",5141 => "11000110",5142 => "00110101",5143 => "00011111",5144 => "00100111",5145 => "00100111",5146 => "10101010",5147 => "00010110",5148 => "10001001",5149 => "00000110",5150 => "00110000",5151 => "10100101",5152 => "11011010",5153 => "10001111",5154 => "10111101",5155 => "11110011",5156 => "11100001",5157 => "01010011",5158 => "11111010",5159 => "10001111",5160 => "01100010",5161 => "01001100",5162 => "11110110",5163 => "10111001",5164 => "01100100",5165 => "11110110",5166 => "00011000",5167 => "10111111",5168 => "01100001",5169 => "11111011",5170 => "10110000",5171 => "11110101",5172 => "10010100",5173 => "11111001",5174 => "00001111",5175 => "10001101",5176 => "01110100",5177 => "11000101",5178 => "10010110",5179 => "00110000",5180 => "00001010",5181 => "11110001",5182 => "00100011",5183 => "00011011",5184 => "00010010",5185 => "01011110",5186 => "00000011",5187 => "11101110",5188 => "00110000",5189 => "01101100",5190 => "11001110",5191 => "00000100",5192 => "11111100",5193 => "01011111",5194 => "11101100",5195 => "10010000",5196 => "10111111",5197 => "01010001",5198 => "00010000",5199 => "11101111",5200 => "11110100",5201 => "11111111",5202 => "11011011",5203 => "00011100",5204 => "10000111",5205 => "10010101",5206 => "01010111",5207 => "10000111",5208 => "11110101",5209 => "10110001",5210 => "11000111",5211 => "01011000",5212 => "11110010",5213 => "01100011",5214 => "11000000",5215 => "01001101",5216 => "10110100",5217 => "00111011",5218 => "01001001",5219 => "10101111",5220 => "11010011",5221 => "00000011",5222 => "01100101",5223 => "10110100",5224 => "00001001",5225 => "01110111",5226 => "10000010",5227 => "00100011",5228 => "01100111",5229 => "01010101",5230 => "00110111",5231 => "01101101",5232 => "10100000",5233 => "00110100",5234 => "01111101",5235 => "11001011",5236 => "01011100",5237 => "11000111",5238 => "10001111",5239 => "10100110",5240 => "10001101",5241 => "11100000",5242 => "11101011",5243 => "01101100",5244 => "00001110",5245 => "01011110",5246 => "11000001",5247 => "00111001",5248 => "10111011",5249 => "10010011",5250 => "01111100",5251 => "10110011",5252 => "00010100",5253 => "11111011",5254 => "01010101",5255 => "10010110",5256 => "01001001",5257 => "01101100",5258 => "10111010",5259 => "10100001",5260 => "11001000",5261 => "00011100",5262 => "10101010",5263 => "11010001",5264 => "01001100",5265 => "10100001",5266 => "10010110",5267 => "11110000",5268 => "00110111",5269 => "00010011",5270 => "10011100",5271 => "00000001",5272 => "11000101",5273 => "11000111",5274 => "11000111",5275 => "10011111",5276 => "10010101",5277 => "00011110",5278 => "10110010",5279 => "10100000",5280 => "11001000",5281 => "11010111",5282 => "10111111",5283 => "10111111",5284 => "11010000",5285 => "11010100",5286 => "10011011",5287 => "01001110",5288 => "00010111",5289 => "10101100",5290 => "10011010",5291 => "00000110",5292 => "01101110",5293 => "01011010",5294 => "01001100",5295 => "00011111",5296 => "00101100",5297 => "01001001",5298 => "11100000",5299 => "10100000",5300 => "00000001",5301 => "11101111",5302 => "11111111",5303 => "10001001",5304 => "11010001",5305 => "01110011",5306 => "00011011",5307 => "01110100",5308 => "01001110",5309 => "00101110",5310 => "01011111",5311 => "11101010",5312 => "01010000",5313 => "11111111",5314 => "10110101",5315 => "11111110",5316 => "01101101",5317 => "00001011",5318 => "01010010",5319 => "10101100",5320 => "00101010",5321 => "11001010",5322 => "11100011",5323 => "00111001",5324 => "01000010",5325 => "01101001",5326 => "01010001",5327 => "11100000",5328 => "01100010",5329 => "01010000",5330 => "11100001",5331 => "10011110",5332 => "11111001",5333 => "10110000",5334 => "00100101",5335 => "01010010",5336 => "01101110",5337 => "00110011",5338 => "01101111",5339 => "11111101",5340 => "10000110",5341 => "00100010",5342 => "00000010",5343 => "10110001",5344 => "10001010",5345 => "11000111",5346 => "11110110",5347 => "01101010",5348 => "01101010",5349 => "00000110",5350 => "10101100",5351 => "01100011",5352 => "00101011",5353 => "00101100",5354 => "10111010",5355 => "10001000",5356 => "10000001",5357 => "00011101",5358 => "10111100",5359 => "11110110",5360 => "01001100",5361 => "00110011",5362 => "10110111",5363 => "11110011",5364 => "11000010",5365 => "10010001",5366 => "10000011",5367 => "00100100",5368 => "00110101",5369 => "01000011",5370 => "01101010",5371 => "01110000",5372 => "00000110",5373 => "11110000",5374 => "01010011",5375 => "01000101",5376 => "00010101",5377 => "11101100",5378 => "01100001",5379 => "00010011",5380 => "01011001",5381 => "01101011",5382 => "10111001",5383 => "10010001",5384 => "00001111",5385 => "01001001",5386 => "00001110",5387 => "01010110",5388 => "11000000",5389 => "11100011",5390 => "10011110",5391 => "11000111",5392 => "10100010",5393 => "01000111",5394 => "10100111",5395 => "11100111",5396 => "01110000",5397 => "01100011",5398 => "00011011",5399 => "01000000",5400 => "01111011",5401 => "11010001",5402 => "00110100",5403 => "00101010",5404 => "01100100",5405 => "10001100",5406 => "01101101",5407 => "11010100",5408 => "01101011",5409 => "01010110",5410 => "10011101",5411 => "10000101",5412 => "11001111",5413 => "11001011",5414 => "11111110",5415 => "01100011",5416 => "00010100",5417 => "11001000",5418 => "00001011",5419 => "00010111",5420 => "00110111",5421 => "01011010",5422 => "10111011",5423 => "00100101",5424 => "01110111",5425 => "01011001",5426 => "11110111",5427 => "10011011",5428 => "00101110",5429 => "01000011",5430 => "10111100",5431 => "10011100",5432 => "00010010",5433 => "01000110",5434 => "10001011",5435 => "11110110",5436 => "11110011",5437 => "01000000",5438 => "10010110",5439 => "10010100",5440 => "11011011",5441 => "11110010",5442 => "10011101",5443 => "00010001",5444 => "11000111",5445 => "00111000",5446 => "11001111",5447 => "11011100",5448 => "01010000",5449 => "10010001",5450 => "11110011",5451 => "11000100",5452 => "11110111",5453 => "00001110",5454 => "10001011",5455 => "01111010",5456 => "00001000",5457 => "00001010",5458 => "10111100",5459 => "01101100",5460 => "11100000",5461 => "11111001",5462 => "01101100",5463 => "10000110",5464 => "01001111",5465 => "01000101",5466 => "00011011",5467 => "11000000",5468 => "01010101",5469 => "11111110",5470 => "11101110",5471 => "11000101",5472 => "00010010",5473 => "00100111",5474 => "00001101",5475 => "10110111",5476 => "01110111",5477 => "10110001",5478 => "00110100",5479 => "10000001",5480 => "00011111",5481 => "11100101",5482 => "00011111",5483 => "01000100",5484 => "00000001",5485 => "11000110",5486 => "01000111",5487 => "01110000",5488 => "01100001",5489 => "10111111",5490 => "01110010",5491 => "00010100",5492 => "01010100",5493 => "10101010",5494 => "11110110",5495 => "10100110",5496 => "00001100",5497 => "00001010",5498 => "11110010",5499 => "00000101",5500 => "01101100",5501 => "10001111",5502 => "11111100",5503 => "10011010",5504 => "01001100",5505 => "00000000",5506 => "00100010",5507 => "01010101",5508 => "01100001",5509 => "00111011",5510 => "00011010",5511 => "10101001",5512 => "01100001",5513 => "00110010",5514 => "10101100",5515 => "10010001",5516 => "11000000",5517 => "11000011",5518 => "11111101",5519 => "01000010",5520 => "00010010",5521 => "10001011",5522 => "01010100",5523 => "01011110",5524 => "00011110",5525 => "10011101",5526 => "01000011",5527 => "01000000",5528 => "10001100",5529 => "10101001",5530 => "00101011",5531 => "00100111",5532 => "11101010",5533 => "00100100",5534 => "10000110",5535 => "01000110",5536 => "00110100",5537 => "00110101",5538 => "01000100",5539 => "11010101",5540 => "00101101",5541 => "00010111",5542 => "01001000",5543 => "10011000",5544 => "10011000",5545 => "00010000",5546 => "01011100",5547 => "01101111",5548 => "00111100",5549 => "11101011",5550 => "00100110",5551 => "01001101",5552 => "00010110",5553 => "00010010",5554 => "10101010",5555 => "10110001",5556 => "00010101",5557 => "01100100",5558 => "11100011",5559 => "01010110",5560 => "00010011",5561 => "01101101",5562 => "00001010",5563 => "11101111",5564 => "11101101",5565 => "01011000",5566 => "10101000",5567 => "01000111",5568 => "11001100",5569 => "01011111",5570 => "10001001",5571 => "00110001",5572 => "00100111",5573 => "01001000",5574 => "01001100",5575 => "00110001",5576 => "00001011",5577 => "11000110",5578 => "00100011",5579 => "00111100",5580 => "00001101",5581 => "01111110",5582 => "11101111",5583 => "01100000",5584 => "11001000",5585 => "11011100",5586 => "11001010",5587 => "11000111",5588 => "11100101",5589 => "10110111",5590 => "11110010",5591 => "11100010",5592 => "00101110",5593 => "01101110",5594 => "11011011",5595 => "10011111",5596 => "11101000",5597 => "10111110",5598 => "11010111",5599 => "11001010",5600 => "11011101",5601 => "11101011",5602 => "11001010",5603 => "11010010",5604 => "01001111",5605 => "10010000",5606 => "10100000",5607 => "01000010",5608 => "10101011",5609 => "10100011",5610 => "11110001",5611 => "11010011",5612 => "10000110",5613 => "00100001",5614 => "10011110",5615 => "11010110",5616 => "11100001",5617 => "11101110",5618 => "01111111",5619 => "11111011",5620 => "10000001",5621 => "01001010",5622 => "00100110",5623 => "01010100",5624 => "11101011",5625 => "01010111",5626 => "01010110",5627 => "00001010",5628 => "01001110",5629 => "11100111",5630 => "11001110",5631 => "01001010",5632 => "01000110",5633 => "01101010",5634 => "10101000",5635 => "00111101",5636 => "01100100",5637 => "10111101",5638 => "01100010",5639 => "01001010",5640 => "11111000",5641 => "00000111",5642 => "00000010",5643 => "11100110",5644 => "00001001",5645 => "01111000",5646 => "01000100",5647 => "01001001",5648 => "00100111",5649 => "00000101",5650 => "00111010",5651 => "11011100",5652 => "01110100",5653 => "10101000",5654 => "00010010",5655 => "01001001",5656 => "01110000",5657 => "00101000",5658 => "00011111",5659 => "00111101",5660 => "00001110",5661 => "00101111",5662 => "00100001",5663 => "10110010",5664 => "01011000",5665 => "11000111",5666 => "11000100",5667 => "00111101",5668 => "00101001",5669 => "01111001",5670 => "00000000",5671 => "10001101",5672 => "10110001",5673 => "01000010",5674 => "10001000",5675 => "01111000",5676 => "01001011",5677 => "00101000",5678 => "10010111",5679 => "11101110",5680 => "00010011",5681 => "00000001",5682 => "11010010",5683 => "10001010",5684 => "01111011",5685 => "01101111",5686 => "11111111",5687 => "01011001",5688 => "11001000",5689 => "01100001",5690 => "10101101",5691 => "10000010",5692 => "01101111",5693 => "00100111",5694 => "00001011",5695 => "01001101",5696 => "00101010",5697 => "10001100",5698 => "11100011",5699 => "01101001",5700 => "11111111",5701 => "10011001",5702 => "01101100",5703 => "00011101",5704 => "01111111",5705 => "11010100",5706 => "10011011",5707 => "00110101",5708 => "01010101",5709 => "10001000",5710 => "11011010",5711 => "11011111",5712 => "11001000",5713 => "11100101",5714 => "11011000",5715 => "11011001",5716 => "11101111",5717 => "01110100",5718 => "01011010",5719 => "01101100",5720 => "00011011",5721 => "01111000",5722 => "00010110",5723 => "01001101",5724 => "10001000",5725 => "10111011",5726 => "11011101",5727 => "11101011",5728 => "01111010",5729 => "01111001",5730 => "11000110",5731 => "01000110",5732 => "10100111",5733 => "11010100",5734 => "00000001",5735 => "00101010",5736 => "11100101",5737 => "01011100",5738 => "11101000",5739 => "10001000",5740 => "00101010",5741 => "10010100",5742 => "10111100",5743 => "01110101",5744 => "10100100",5745 => "01111101",5746 => "01011011",5747 => "00001111",5748 => "10000111",5749 => "11011110",5750 => "10111011",5751 => "11000111",5752 => "00100010",5753 => "00011010",5754 => "10111010",5755 => "01000110",5756 => "00111100",5757 => "10110110",5758 => "00010111",5759 => "10100011",5760 => "11111010",5761 => "01001101",5762 => "11011000",5763 => "00110000",5764 => "10001000",5765 => "01000010",5766 => "01111000",5767 => "11100110",5768 => "10100000",5769 => "10100010",5770 => "01001111",5771 => "00101010",5772 => "01111000",5773 => "11010110",5774 => "11001100",5775 => "01001111",5776 => "01100001",5777 => "01100100",5778 => "11001110",5779 => "10101000",5780 => "11110110",5781 => "11011111",5782 => "10010000",5783 => "11010111",5784 => "10010010",5785 => "10011000",5786 => "10100100",5787 => "00101011",5788 => "11111010",5789 => "11000111",5790 => "00000011",5791 => "10100101",5792 => "11001101",5793 => "00000001",5794 => "11110000",5795 => "01001110",5796 => "00100010",5797 => "00100100",5798 => "11100101",5799 => "00011110",5800 => "10000000",5801 => "00011010",5802 => "11100010",5803 => "10000110",5804 => "10011111",5805 => "00101100",5806 => "00011110",5807 => "11111101",5808 => "01111100",5809 => "00000001",5810 => "00001101",5811 => "11101011",5812 => "00101000",5813 => "01111001",5814 => "00100101",5815 => "10110101",5816 => "00110010",5817 => "01101101",5818 => "00010000",5819 => "10101100",5820 => "10001010",5821 => "01000100",5822 => "01111101",5823 => "01010011",5824 => "00100101",5825 => "11001100",5826 => "11010011",5827 => "11100110",5828 => "01100010",5829 => "11100001",5830 => "01110011",5831 => "01101011",5832 => "11100010",5833 => "11010001",5834 => "10110100",5835 => "10001111",5836 => "11101010",5837 => "10111111",5838 => "10011111",5839 => "00011010",5840 => "11100001",5841 => "00000000",5842 => "10010010",5843 => "01010001",5844 => "10010101",5845 => "01101010",5846 => "01100010",5847 => "10101111",5848 => "11000101",5849 => "11000011",5850 => "11111111",5851 => "00110110",5852 => "00011101",5853 => "01110001",5854 => "00110110",5855 => "01000101",5856 => "10011111",5857 => "01011101",5858 => "00100100",5859 => "01010010",5860 => "10100110",5861 => "11111010",5862 => "00000000",5863 => "11100110",5864 => "10010011",5865 => "10001000",5866 => "00100010",5867 => "10000110",5868 => "11101000",5869 => "11110110",5870 => "10000011",5871 => "11000011",5872 => "11110010",5873 => "11010100",5874 => "00001100",5875 => "01001110",5876 => "01011010",5877 => "01100100",5878 => "10011010",5879 => "11111001",5880 => "01101111",5881 => "11011101",5882 => "01000101",5883 => "00000110",5884 => "01000000",5885 => "00100100",5886 => "01111011",5887 => "10011100",5888 => "01000001",5889 => "11000000",5890 => "01011111",5891 => "01101101",5892 => "11000001",5893 => "10010010",5894 => "11001010",5895 => "10001000",5896 => "00110111",5897 => "10011000",5898 => "10100101",5899 => "10100000",5900 => "01101110",5901 => "00111110",5902 => "01110001",5903 => "11110011",5904 => "00001011",5905 => "11000111",5906 => "01001111",5907 => "00011100",5908 => "10100111",5909 => "01000000",5910 => "10000011",5911 => "10011011",5912 => "11000100",5913 => "00110110",5914 => "00000001",5915 => "01010011",5916 => "10101100",5917 => "01101110",5918 => "00111101",5919 => "10000100",5920 => "10111111",5921 => "00000011",5922 => "11011010",5923 => "01010101",5924 => "11110101",5925 => "01110111",5926 => "11111010",5927 => "00100001",5928 => "00111110",5929 => "10000100",5930 => "01011100",5931 => "10111110",5932 => "01100000",5933 => "00110100",5934 => "11000110",5935 => "00010111",5936 => "10100000",5937 => "00000011",5938 => "11001011",5939 => "01101100",5940 => "00101001",5941 => "10010011",5942 => "10011010",5943 => "01110001",5944 => "10111110",5945 => "00111011",5946 => "01100110",5947 => "11101001",5948 => "00101001",5949 => "00111011",5950 => "10000010",5951 => "10100111",5952 => "01100110",5953 => "00101011",5954 => "01111110",5955 => "11100000",5956 => "10111110",5957 => "10010010",5958 => "00000011",5959 => "01011100",5960 => "00100110",5961 => "00101010",5962 => "01011010",5963 => "01011111",5964 => "11000000",5965 => "01001111",5966 => "10100110",5967 => "01000100",5968 => "00000110",5969 => "11100110",5970 => "00000000",5971 => "11011110",5972 => "01001011",5973 => "10010001",5974 => "11010011",5975 => "11010101",5976 => "11110101",5977 => "00010100",5978 => "11111001",5979 => "01011111",5980 => "11100011",5981 => "00100100",5982 => "11100100",5983 => "00100101",5984 => "01110100",5985 => "10000010",5986 => "10001101",5987 => "10001011",5988 => "00111110",5989 => "00011111",5990 => "00001111",5991 => "01010111",5992 => "10101001",5993 => "00001110",5994 => "10001111",5995 => "11000000",5996 => "01111010",5997 => "10110000",5998 => "10101111",5999 => "11001010",6000 => "00010011",6001 => "10101001",6002 => "11100010",6003 => "00010010",6004 => "00100010",6005 => "01000011",6006 => "10100000",6007 => "00111100",6008 => "10101001",6009 => "00110010",6010 => "00011110",6011 => "10000110",6012 => "11001110",6013 => "00000101",6014 => "11100010",6015 => "11111001",6016 => "00000010",6017 => "11100110",6018 => "01000001",6019 => "01100100",6020 => "11101100",6021 => "01110001",6022 => "01101000",6023 => "00000011",6024 => "00111001",6025 => "11100000",6026 => "11000111",6027 => "10001111",6028 => "00110101",6029 => "11110000",6030 => "00000010",6031 => "10110001",6032 => "00000100",6033 => "01000001",6034 => "00010100",6035 => "01000000",6036 => "11110111",6037 => "01111101",6038 => "11100101",6039 => "11001111",6040 => "00000111",6041 => "01010111",6042 => "11001110",6043 => "00010001",6044 => "11001100",6045 => "10110110",6046 => "01010111",6047 => "01001100",6048 => "10001100",6049 => "10011110",6050 => "11010101",6051 => "11000101",6052 => "00110111",6053 => "11010100",6054 => "11000100",6055 => "01001101",6056 => "11101111",6057 => "00010010",6058 => "01011010",6059 => "00110011",6060 => "10111101",6061 => "00110001",6062 => "11000000",6063 => "00101110",6064 => "00110101",6065 => "10111000",6066 => "10110001",6067 => "00111100",6068 => "10011110",6069 => "00011100",6070 => "00110010",6071 => "10111000",6072 => "01011100",6073 => "10000011",6074 => "00010010",6075 => "00000000",6076 => "11000111",6077 => "00000010",6078 => "00011111",6079 => "00001001",6080 => "00100101",6081 => "10101001",6082 => "01100110",6083 => "01010011",6084 => "00000100",6085 => "01111000",6086 => "11011101",6087 => "10100011",6088 => "01011000",6089 => "00110001",6090 => "00110100",6091 => "01000110",6092 => "01111100",6093 => "11000001",6094 => "00111001",6095 => "10001111",6096 => "01000100",6097 => "01011000",6098 => "00010001",6099 => "00111101",6100 => "10001110",6101 => "10001010",6102 => "11010111",6103 => "00011000",6104 => "11111100",6105 => "00000000",6106 => "00010011",6107 => "10001001",6108 => "10110100",6109 => "10000010",6110 => "00100111",6111 => "10010100",6112 => "01010111",6113 => "00101000",6114 => "00111000",6115 => "10111001",6116 => "10101110",6117 => "01010111",6118 => "11101110",6119 => "10111000",6120 => "10111000",6121 => "11100001",6122 => "01101001",6123 => "01000011",6124 => "10011101",6125 => "00100100",6126 => "01101010",6127 => "01011001",6128 => "01100110",6129 => "10001011",6130 => "11001011",6131 => "01101011",6132 => "01100001",6133 => "00100000",6134 => "01010101",6135 => "10000101",6136 => "10111101",6137 => "01010100",6138 => "01010111",6139 => "01110011",6140 => "00110000",6141 => "10000000",6142 => "11010001",6143 => "00111100",6144 => "01011001",6145 => "01001101",6146 => "01101000",6147 => "11110001",6148 => "10110101",6149 => "00001101",6150 => "00111100",6151 => "01110101",6152 => "10111101",6153 => "01100111",6154 => "00111100",6155 => "01101011",6156 => "01101010",6157 => "00000111",6158 => "01100100",6159 => "01111110",6160 => "11110111",6161 => "00010011",6162 => "10100111",6163 => "00101000",6164 => "00010110",6165 => "10011101",6166 => "10100110",6167 => "01011110",6168 => "11001111",6169 => "00001101",6170 => "10010010",6171 => "01101000",6172 => "11111100",6173 => "00100001",6174 => "11111011",6175 => "10110110",6176 => "11001000",6177 => "11000011",6178 => "11100110",6179 => "01110100",6180 => "11000111",6181 => "10110001",6182 => "11010011",6183 => "11101001",6184 => "10001010",6185 => "01001001",6186 => "10101100",6187 => "10100010",6188 => "00111011",6189 => "01110100",6190 => "00101110",6191 => "11000100",6192 => "00010111",6193 => "11111010",6194 => "11011011",6195 => "10101100",6196 => "00111100",6197 => "01100101",6198 => "11011101",6199 => "01100111",6200 => "00000110",6201 => "01000100",6202 => "01001101",6203 => "10110011",6204 => "00100100",6205 => "10001101",6206 => "11100110",6207 => "01000010",6208 => "00101111",6209 => "10001101",6210 => "11110110",6211 => "11110101",6212 => "00111001",6213 => "11100000",6214 => "11011011",6215 => "01110001",6216 => "11100000",6217 => "11100000",6218 => "00100100",6219 => "00100111",6220 => "11010001",6221 => "11001111",6222 => "00100010",6223 => "00100000",6224 => "10001001",6225 => "01100110",6226 => "01100001",6227 => "00100010",6228 => "11100111",6229 => "01101101",6230 => "10010111",6231 => "11010101",6232 => "01011000",6233 => "00110100",6234 => "10110111",6235 => "10100110",6236 => "10100111",6237 => "10110010",6238 => "11000011",6239 => "10111010",6240 => "01011111",6241 => "00110001",6242 => "10110011",6243 => "01001010",6244 => "01101110",6245 => "10010100",6246 => "00110110",6247 => "10100001",6248 => "00001110",6249 => "01010110",6250 => "10111011",6251 => "10111001",6252 => "01001000",6253 => "01101101",6254 => "11011000",6255 => "01111001",6256 => "11101100",6257 => "01010111",6258 => "11101010",6259 => "11010010",6260 => "00010011",6261 => "00000001",6262 => "01010110",6263 => "11000011",6264 => "01000111",6265 => "10101000",6266 => "01110000",6267 => "11001010",6268 => "00010111",6269 => "00110110",6270 => "01111100",6271 => "01001110",6272 => "10110110",6273 => "01101000",6274 => "01111001",6275 => "11001000",6276 => "10001111",6277 => "00110001",6278 => "10111111",6279 => "11100110",6280 => "11101101",6281 => "11010011",6282 => "10101010",6283 => "00000001",6284 => "10000010",6285 => "11001011",6286 => "01111011",6287 => "01110010",6288 => "10101010",6289 => "10010010",6290 => "10001101",6291 => "11010111",6292 => "10101010",6293 => "10101011",6294 => "00001000",6295 => "01010101",6296 => "10010100",6297 => "00111011",6298 => "01000001",6299 => "00000001",6300 => "01001100",6301 => "11101000",6302 => "00011010",6303 => "01001000",6304 => "11000011",6305 => "10001110",6306 => "00111111",6307 => "10101001",6308 => "00111000",6309 => "10001001",6310 => "11100110",6311 => "11101011",6312 => "01000100",6313 => "01110010",6314 => "10111001",6315 => "01000100",6316 => "11001101",6317 => "10110100",6318 => "00101110",6319 => "11001110",6320 => "10000000",6321 => "00011101",6322 => "11011111",6323 => "10100100",6324 => "01000010",6325 => "00100011",6326 => "01000001",6327 => "01011011",6328 => "01001110",6329 => "01110110",6330 => "11001000",6331 => "01101010",6332 => "10110110",6333 => "10110101",6334 => "11100110",6335 => "11011101",6336 => "11001111",6337 => "00100100",6338 => "01101000",6339 => "01111100",6340 => "10101101",6341 => "10011101",6342 => "00000111",6343 => "11111001",6344 => "00011100",6345 => "10100010",6346 => "11111111",6347 => "01011111",6348 => "10101101",6349 => "11111010",6350 => "00001000",6351 => "01010100",6352 => "10101110",6353 => "01110000",6354 => "00110011",6355 => "00011001",6356 => "01111101",6357 => "11110011",6358 => "00000100",6359 => "11111011",6360 => "11011010",6361 => "10101000",6362 => "10001011",6363 => "11010101",6364 => "00001110",6365 => "01010101",6366 => "00011011",6367 => "11010101",6368 => "01110110",6369 => "11100010",6370 => "00011010",6371 => "10011101",6372 => "01101111",6373 => "10111110",6374 => "11101110",6375 => "00011111",6376 => "10101011",6377 => "00010101",6378 => "00101010",6379 => "01100011",6380 => "10000111",6381 => "00000011",6382 => "10111100",6383 => "11001011",6384 => "01101010",6385 => "01100011",6386 => "00111111",6387 => "01100001",6388 => "00100101",6389 => "00011001",6390 => "11110110",6391 => "00000011",6392 => "10000110",6393 => "10010010",6394 => "10010110",6395 => "11001100",6396 => "10001000",6397 => "11111001",6398 => "00010011",6399 => "10001000",6400 => "01110110",6401 => "00011000",6402 => "00000011",6403 => "11001100",6404 => "01010001",6405 => "00000001",6406 => "10011101",6407 => "01011010",6408 => "11010000",6409 => "11110000",6410 => "11011110",6411 => "10101011",6412 => "10110001",6413 => "00000110",6414 => "01000100",6415 => "11001011",6416 => "11100111",6417 => "00101110",6418 => "11111111",6419 => "00010000",6420 => "10000110",6421 => "01101010",6422 => "00110111",6423 => "11000011",6424 => "11110110",6425 => "00110010",6426 => "00100100",6427 => "11000111",6428 => "11000001",6429 => "10010110",6430 => "10001101",6431 => "11100111",6432 => "00100100",6433 => "11001001",6434 => "11111110",6435 => "00011100",6436 => "01001100",6437 => "11101011",6438 => "00111010",6439 => "10001001",6440 => "00100111",6441 => "01011111",6442 => "01000101",6443 => "00100100",6444 => "01101010",6445 => "00100101",6446 => "10001011",6447 => "00111000",6448 => "01111010",6449 => "11010110",6450 => "00101001",6451 => "00010011",6452 => "00011111",6453 => "11001000",6454 => "00001111",6455 => "00010000",6456 => "11101100",6457 => "10100101",6458 => "11000111",6459 => "01010110",6460 => "00101011",6461 => "10001010",6462 => "11000111",6463 => "00000011",6464 => "11000011",6465 => "00110101",6466 => "00110100",6467 => "00011000",6468 => "00001000",6469 => "01111001",6470 => "11001100",6471 => "10100010",6472 => "11111010",6473 => "11100001",6474 => "01001011",6475 => "00010000",6476 => "10101001",6477 => "11101000",6478 => "10010011",6479 => "11001011",6480 => "10011000",6481 => "11100100",6482 => "00101010",6483 => "01110110",6484 => "10011010",6485 => "10010100",6486 => "10110101",6487 => "00101111",6488 => "10111001",6489 => "00111011",6490 => "11000010",6491 => "11001111",6492 => "00111010",6493 => "11000000",6494 => "11010110",6495 => "11110100",6496 => "01110110",6497 => "00011001",6498 => "10110001",6499 => "10111010",6500 => "11001011",6501 => "00111011",6502 => "00000111",6503 => "01000001",6504 => "10111011",6505 => "11101111",6506 => "01111101",6507 => "10000101",6508 => "00111000",6509 => "01011011",6510 => "10010101",6511 => "11110011",6512 => "10110101",6513 => "01010110",6514 => "11000010",6515 => "10011000",6516 => "11001110",6517 => "10001000",6518 => "00100001",6519 => "00111100",6520 => "11000010",6521 => "01010100",6522 => "01010111",6523 => "01110000",6524 => "11100011",6525 => "00001101",6526 => "10010100",6527 => "00111011",6528 => "11111000",6529 => "00001111",6530 => "01111000",6531 => "00010100",6532 => "10011110",6533 => "00110000",6534 => "00101010",6535 => "01100100",6536 => "11111111",6537 => "11101111",6538 => "01000011",6539 => "10000000",6540 => "00110001",6541 => "11110101",6542 => "10101111",6543 => "11000111",6544 => "00101000",6545 => "01110100",6546 => "11011001",6547 => "01100101",6548 => "01010000",6549 => "01111000",6550 => "00101101",6551 => "11001011",6552 => "10001011",6553 => "10111001",6554 => "11101011",6555 => "10110110",6556 => "00000000",6557 => "01011111",6558 => "01011010",6559 => "00101011",6560 => "10011011",6561 => "10011101",6562 => "00001111",6563 => "00111101",6564 => "01011011",6565 => "11111101",6566 => "11111011",6567 => "11110111",6568 => "01110001",6569 => "00010100",6570 => "11111101",6571 => "11000001",6572 => "00000110",6573 => "00101110",6574 => "01101010",6575 => "10011001",6576 => "00101111",6577 => "00010100",6578 => "01100101",6579 => "10110000",6580 => "11010110",6581 => "01010101",6582 => "11000110",6583 => "01010001",6584 => "00100101",6585 => "00001101",6586 => "01001111",6587 => "10000110",6588 => "00110101",6589 => "11011011",6590 => "10000110",6591 => "10111110",6592 => "00001001",6593 => "00101001",6594 => "01011000",6595 => "00110111",6596 => "01011000",6597 => "10100110",6598 => "10100011",6599 => "10110000",6600 => "10010111",6601 => "00001100",6602 => "11110111",6603 => "00000010",6604 => "01011111",6605 => "00010000",6606 => "10000000",6607 => "00011101",6608 => "00011101",6609 => "11100011",6610 => "10011101",6611 => "00110010",6612 => "10110111",6613 => "11011000",6614 => "01110100",6615 => "00111010",6616 => "00100010",6617 => "10000000",6618 => "01111010",6619 => "11100001",6620 => "01011101",6621 => "11100011",6622 => "00010110",6623 => "00011000",6624 => "00010000",6625 => "00000000",6626 => "01110100",6627 => "11010010",6628 => "00110000",6629 => "00000100",6630 => "10001011",6631 => "01101111",6632 => "00100001",6633 => "01111010",6634 => "11100000",6635 => "11010100",6636 => "00100010",6637 => "01111100",6638 => "01110011",6639 => "01001001",6640 => "01000000",6641 => "11110010",6642 => "00001100",6643 => "00011110",6644 => "11100010",6645 => "01110011",6646 => "01001100",6647 => "01100011",6648 => "00110001",6649 => "00100010",6650 => "11101110",6651 => "00010100",6652 => "00001101",6653 => "11111001",6654 => "01110111",6655 => "11011001",6656 => "00101011",6657 => "00110010",6658 => "10111100",6659 => "10000010",6660 => "01110010",6661 => "01101100",6662 => "01110000",6663 => "01000010",6664 => "10001110",6665 => "10110101",6666 => "01110100",6667 => "10101010",6668 => "00000110",6669 => "01011000",6670 => "01011000",6671 => "10111110",6672 => "11100001",6673 => "10010010",6674 => "11010001",6675 => "01001000",6676 => "11101010",6677 => "10110000",6678 => "01101100",6679 => "10111110",6680 => "01110000",6681 => "10001100",6682 => "11101100",6683 => "00101101",6684 => "10001101",6685 => "01111001",6686 => "00011100",6687 => "10010000",6688 => "10000111",6689 => "00111000",6690 => "10110010",6691 => "11110110",6692 => "00100111",6693 => "10111011",6694 => "01101010",6695 => "10100100",6696 => "00001000",6697 => "00011001",6698 => "10011011",6699 => "11010011",6700 => "00010000",6701 => "00110000",6702 => "11110111",6703 => "01001010",6704 => "00010110",6705 => "01110100",6706 => "11101100",6707 => "10001001",6708 => "00011111",6709 => "01001100",6710 => "00010011",6711 => "01000100",6712 => "01110011",6713 => "01100001",6714 => "11001011",6715 => "11001110",6716 => "01000111",6717 => "11100111",6718 => "10011000",6719 => "00101100",6720 => "00111110",6721 => "01001000",6722 => "11100011",6723 => "10010101",6724 => "10111111",6725 => "11101101",6726 => "11100010",6727 => "10111101",6728 => "01000110",6729 => "00011110",6730 => "11110100",6731 => "11111011",6732 => "00001000",6733 => "10110010",6734 => "11110100",6735 => "11000011",6736 => "11111010",6737 => "10111101",6738 => "10110011",6739 => "01100000",6740 => "01111001",6741 => "11001001",6742 => "10100101",6743 => "11011000",6744 => "10000011",6745 => "11101011",6746 => "01110000",6747 => "11111001",6748 => "00011000",6749 => "10001100",6750 => "10010111",6751 => "11011111",6752 => "00001110",6753 => "10011011",6754 => "00101100",6755 => "11001100",6756 => "01111101",6757 => "10000111",6758 => "11101100",6759 => "00010011",6760 => "11000101",6761 => "10011011",6762 => "01110001",6763 => "00000010",6764 => "01111001",6765 => "11010110",6766 => "00000100",6767 => "11101011",6768 => "10100100",6769 => "10011010",6770 => "00011111",6771 => "00100011",6772 => "10000100",6773 => "01001000",6774 => "01001100",6775 => "01101111",6776 => "10100111",6777 => "11010101",6778 => "00000010",6779 => "01101000",6780 => "10001000",6781 => "10001110",6782 => "10001100",6783 => "00011100",6784 => "11011011",6785 => "01001110",6786 => "00101110",6787 => "00111011",6788 => "01000110",6789 => "10001011",6790 => "00111101",6791 => "00100100",6792 => "10001100",6793 => "11001000",6794 => "01010101",6795 => "01111110",6796 => "10111000",6797 => "01010000",6798 => "11011110",6799 => "10011011",6800 => "10101101",6801 => "01001000",6802 => "01111011",6803 => "00110111",6804 => "01001110",6805 => "01100000",6806 => "01110111",6807 => "00101001",6808 => "11111010",6809 => "00010000",6810 => "10100010",6811 => "11001110",6812 => "00001011",6813 => "11110101",6814 => "00000010",6815 => "11000111",6816 => "01001111",6817 => "10111010",6818 => "01100001",6819 => "10110100",6820 => "01010110",6821 => "10110010",6822 => "10111110",6823 => "01111000",6824 => "10000001",6825 => "11011111",6826 => "11101001",6827 => "11101000",6828 => "10111011",6829 => "11010101",6830 => "11100110",6831 => "10101110",6832 => "10000001",6833 => "01110011",6834 => "11101010",6835 => "11000011",6836 => "10000010",6837 => "00100111",6838 => "10001100",6839 => "11000001",6840 => "11001001",6841 => "00010001",6842 => "10001101",6843 => "10011011",6844 => "11110000",6845 => "00111011",6846 => "01101111",6847 => "10000010",6848 => "11011001",6849 => "00001001",6850 => "00011111",6851 => "10100101",6852 => "10001010",6853 => "01000101",6854 => "00010000",6855 => "10111110",6856 => "01110110",6857 => "01010110",6858 => "10011010",6859 => "11010000",6860 => "11101010",6861 => "00111000",6862 => "01101101",6863 => "01011100",6864 => "00001011",6865 => "10101010",6866 => "11000000",6867 => "10000100",6868 => "10111000",6869 => "01101011",6870 => "01111101",6871 => "10010000",6872 => "00110111",6873 => "10011011",6874 => "10101110",6875 => "11100010",6876 => "01011101",6877 => "01000001",6878 => "01110001",6879 => "00111110",6880 => "01000001",6881 => "01110010",6882 => "01110010",6883 => "01011000",6884 => "11000010",6885 => "01011011",6886 => "11010010",6887 => "11110000",6888 => "11010101",6889 => "00101011",6890 => "00011110",6891 => "11110100",6892 => "00011111",6893 => "10100000",6894 => "11111111",6895 => "01101011",6896 => "11110101",6897 => "10010000",6898 => "01101110",6899 => "11001001",6900 => "11011101",6901 => "10001111",6902 => "11000100",6903 => "01011101",6904 => "01001100",6905 => "00111101",6906 => "00010110",6907 => "01000000",6908 => "10100000",6909 => "00110011",6910 => "11010001",6911 => "00101111",6912 => "01001100",6913 => "01101111",6914 => "00101100",6915 => "00000100",6916 => "10101101",6917 => "11101000",6918 => "11100000",6919 => "10101110",6920 => "11001000",6921 => "11001111",6922 => "10101110",6923 => "00101111",6924 => "00010000",6925 => "01100001",6926 => "10111110",6927 => "00001001",6928 => "01010001",6929 => "00110100",6930 => "10101000",6931 => "11000101",6932 => "11000010",6933 => "10010110",6934 => "11000101",6935 => "01101001",6936 => "11100100",6937 => "11011110",6938 => "10100001",6939 => "11111001",6940 => "01000111",6941 => "01001100",6942 => "10100010",6943 => "10001001",6944 => "11101101",6945 => "01001101",6946 => "01110001",6947 => "10101010",6948 => "01001110",6949 => "10101100",6950 => "10001000",6951 => "10011111",6952 => "00100100",6953 => "01101000",6954 => "00011000",6955 => "10111011",6956 => "11100010",6957 => "00100110",6958 => "11101010",6959 => "10111111",6960 => "01110010",6961 => "01110001",6962 => "00010110",6963 => "10110100",6964 => "00000110",6965 => "11111001",6966 => "00111101",6967 => "11111100",6968 => "00011110",6969 => "01011001",6970 => "10010110",6971 => "00001000",6972 => "10010110",6973 => "00110110",6974 => "00011111",6975 => "10000100",6976 => "01001011",6977 => "11111110",6978 => "00110111",6979 => "00000110",6980 => "11010000",6981 => "00111010",6982 => "11111111",6983 => "11000100",6984 => "01011000",6985 => "10110001",6986 => "11000100",6987 => "01000111",6988 => "10000011",6989 => "01110011",6990 => "01010110",6991 => "10001111",6992 => "00100011",6993 => "00101010",6994 => "10011110",6995 => "01110111",6996 => "00010110",6997 => "00100000",6998 => "10101101",6999 => "00111011",7000 => "10101000",7001 => "00001100",7002 => "01000001",7003 => "01010101",7004 => "10011110",7005 => "01111101",7006 => "00001111",7007 => "10000110",7008 => "10000111",7009 => "10010101",7010 => "00111101",7011 => "00111101",7012 => "00011011",7013 => "11011100",7014 => "00011100",7015 => "00100000",7016 => "10011110",7017 => "00111011",7018 => "10001000",7019 => "11011110",7020 => "00100110",7021 => "00110111",7022 => "10111000",7023 => "01101000",7024 => "00100111",7025 => "01010101",7026 => "01100111",7027 => "11000111",7028 => "11111111",7029 => "00110010",7030 => "00100111",7031 => "11010100",7032 => "11000001",7033 => "10011010",7034 => "11111010",7035 => "10011010",7036 => "10010110",7037 => "00011000",7038 => "01101110",7039 => "00111110",7040 => "10001100",7041 => "10010010",7042 => "01101110",7043 => "10011101",7044 => "01100011",7045 => "01110001",7046 => "01101000",7047 => "11000010",7048 => "00111011",7049 => "01110110",7050 => "11100101",7051 => "00101001",7052 => "11010010",7053 => "11010110",7054 => "01000101",7055 => "10010000",7056 => "10101110",7057 => "00110110",7058 => "01001011",7059 => "10010111",7060 => "01000110",7061 => "11001101",7062 => "10011011",7063 => "10001010",7064 => "01111110",7065 => "11001011",7066 => "11101010",7067 => "11111101",7068 => "00110100",7069 => "10010001",7070 => "10000100",7071 => "11000000",7072 => "00110011",7073 => "11111100",7074 => "00100010",7075 => "00011000",7076 => "10001010",7077 => "01110010",7078 => "10000100",7079 => "11000101",7080 => "01111111",7081 => "10100000",7082 => "11111001",7083 => "01101001",7084 => "01010010",7085 => "11101100",7086 => "11000110",7087 => "10110101",7088 => "11111010",7089 => "10110111",7090 => "00010010",7091 => "01110110",7092 => "10101001",7093 => "01010101",7094 => "11111101",7095 => "10010100",7096 => "11001100",7097 => "01100110",7098 => "10101110",7099 => "11011101",7100 => "00000101",7101 => "01001011",7102 => "01101001",7103 => "11100110",7104 => "11110110",7105 => "00000000",7106 => "00000101",7107 => "10000111",7108 => "00100101",7109 => "11010011",7110 => "00110111",7111 => "01101101",7112 => "11001101",7113 => "10110001",7114 => "00010111",7115 => "11011001",7116 => "10111100",7117 => "01000110",7118 => "01111100",7119 => "01111011",7120 => "10100111",7121 => "11001001",7122 => "11101110",7123 => "01100110",7124 => "11011101",7125 => "11111100",7126 => "11111011",7127 => "01100000",7128 => "11100111",7129 => "01000011",7130 => "11111101",7131 => "01010110",7132 => "00110110",7133 => "01000011",7134 => "11100101",7135 => "10010100",7136 => "01001100",7137 => "10101011",7138 => "00110100",7139 => "00010000",7140 => "11101011",7141 => "10011001",7142 => "00010110",7143 => "10011010",7144 => "00000101",7145 => "00110101",7146 => "11101011",7147 => "10010111",7148 => "00001000",7149 => "11010111",7150 => "11110011",7151 => "10101010",7152 => "11001100",7153 => "10101111",7154 => "11101110",7155 => "10100111",7156 => "00011100",7157 => "01110100",7158 => "10011100",7159 => "10010001",7160 => "00000101",7161 => "01001010",7162 => "00001111",7163 => "01111001",7164 => "00000101",7165 => "00100001",7166 => "11011000",7167 => "11001010",7168 => "00000010",7169 => "11001101",7170 => "00001101",7171 => "11110011",7172 => "10000111",7173 => "00100101",7174 => "11011011",7175 => "01110100",7176 => "10100001",7177 => "00001010",7178 => "11101011",7179 => "10100111",7180 => "01001111",7181 => "00000111",7182 => "10001111",7183 => "10011111",7184 => "00111100",7185 => "01110010",7186 => "10000101",7187 => "10101001",7188 => "00000101",7189 => "10100110",7190 => "01010010",7191 => "11100011",7192 => "10010011",7193 => "00011100",7194 => "11010011",7195 => "01110000",7196 => "01010111",7197 => "10000100",7198 => "01001110",7199 => "01001101",7200 => "01111000",7201 => "01100000",7202 => "11010011",7203 => "11001010",7204 => "11000010",7205 => "10011000",7206 => "01011001",7207 => "01101011",7208 => "11110010",7209 => "01000010",7210 => "00001101",7211 => "00010000",7212 => "01100011",7213 => "11010110",7214 => "11001011",7215 => "11101101",7216 => "01111110",7217 => "01110111",7218 => "10010000",7219 => "10011101",7220 => "00011010",7221 => "11001001",7222 => "11000110",7223 => "01000000",7224 => "01010111",7225 => "11110110",7226 => "01011000",7227 => "01011110",7228 => "11001110",7229 => "11101110",7230 => "11111010",7231 => "00010111",7232 => "11011011",7233 => "11110001",7234 => "10001111",7235 => "10101000",7236 => "00101011",7237 => "10110101",7238 => "10100000",7239 => "10011010",7240 => "10100000",7241 => "01110010",7242 => "01011110",7243 => "11101000",7244 => "11111110",7245 => "01000110",7246 => "00001110",7247 => "00110101",7248 => "01100011",7249 => "11001001",7250 => "10010101",7251 => "01011100",7252 => "00110000",7253 => "10110011",7254 => "10110000",7255 => "00100000",7256 => "10001011",7257 => "11011010",7258 => "01000001",7259 => "01011000",7260 => "00111010",7261 => "11001010",7262 => "11000000",7263 => "11101010",7264 => "00000101",7265 => "01010101",7266 => "01000010",7267 => "01100110",7268 => "01110101",7269 => "11000101",7270 => "01011111",7271 => "00000101",7272 => "10001000",7273 => "00100101",7274 => "00110110",7275 => "11100111",7276 => "11010101",7277 => "00001110",7278 => "10100011",7279 => "11111111",7280 => "10011101",7281 => "01101111",7282 => "01010110",7283 => "01101001",7284 => "00111001",7285 => "01111001",7286 => "00001100",7287 => "01111110",7288 => "11001101",7289 => "00110000",7290 => "11110000",7291 => "10010000",7292 => "01111010",7293 => "10010000",7294 => "01110001",7295 => "11001100",7296 => "11011111",7297 => "00101001",7298 => "10101100",7299 => "00010010",7300 => "00111010",7301 => "01101111",7302 => "11101010",7303 => "10010101",7304 => "00011011",7305 => "10100000",7306 => "11011100",7307 => "01100101",7308 => "10011010",7309 => "01100111",7310 => "11100000",7311 => "01111011",7312 => "10100010",7313 => "01101110",7314 => "11001110",7315 => "11001100",7316 => "11011010",7317 => "01100001",7318 => "01110100",7319 => "10010010",7320 => "00001100",7321 => "00111000",7322 => "01010011",7323 => "01000001",7324 => "00011100",7325 => "11110101",7326 => "01111101",7327 => "10010111",7328 => "01110111",7329 => "00011110",7330 => "10110111",7331 => "00000111",7332 => "10010101",7333 => "10001000",7334 => "11000001",7335 => "10100110",7336 => "10000101",7337 => "10000111",7338 => "01111100",7339 => "11101000",7340 => "10101111",7341 => "00100010",7342 => "00111010",7343 => "11110000",7344 => "11111001",7345 => "11111001",7346 => "11110100",7347 => "01010011",7348 => "01000011",7349 => "11010100",7350 => "00101101",7351 => "01101110",7352 => "10011111",7353 => "11001110",7354 => "01100110",7355 => "10110111",7356 => "10000100",7357 => "10101101",7358 => "01001111",7359 => "01100101",7360 => "00000001",7361 => "01001010",7362 => "01011101",7363 => "10011100",7364 => "11001011",7365 => "01100111",7366 => "00000000",7367 => "10010110",7368 => "00000000",7369 => "11111000",7370 => "11101000",7371 => "11110100",7372 => "10100001",7373 => "10101100",7374 => "10111101",7375 => "11001001",7376 => "10000011",7377 => "10010100",7378 => "00110101",7379 => "01100100",7380 => "10000010",7381 => "10011100",7382 => "10100010",7383 => "10010111",7384 => "10110100",7385 => "11101011",7386 => "10010100",7387 => "00101110",7388 => "10101100",7389 => "00101101",7390 => "10011101",7391 => "01001100",7392 => "10000110",7393 => "01111000",7394 => "11010101",7395 => "11100001",7396 => "01100101",7397 => "01011000",7398 => "10010010",7399 => "10000000",7400 => "01001111",7401 => "00010101",7402 => "11011110",7403 => "11101011",7404 => "01001100",7405 => "10110000",7406 => "11100011",7407 => "00111011",7408 => "11100010",7409 => "10001011",7410 => "01000001",7411 => "00101001",7412 => "00011110",7413 => "01000110",7414 => "11111110",7415 => "11110100",7416 => "00100100",7417 => "11111000",7418 => "10000111",7419 => "01100101",7420 => "11010100",7421 => "11110111",7422 => "10111111",7423 => "11011100",7424 => "10001110",7425 => "10101101",7426 => "10010010",7427 => "11101011",7428 => "01011111",7429 => "01101111",7430 => "01000011",7431 => "10111010",7432 => "11101001",7433 => "10111110",7434 => "11001001",7435 => "10011011",7436 => "01000110",7437 => "11100001",7438 => "11110011",7439 => "11101010",7440 => "00101111",7441 => "11000100",7442 => "10011101",7443 => "00001110",7444 => "11110000",7445 => "10110010",7446 => "01101011",7447 => "01110010",7448 => "10100011",7449 => "11110010",7450 => "11010011",7451 => "00000001",7452 => "10110101",7453 => "11010110",7454 => "00011101",7455 => "11100010",7456 => "00101101",7457 => "11010001",7458 => "11100011",7459 => "11001011",7460 => "00101010",7461 => "11001110",7462 => "01011101",7463 => "01111001",7464 => "10001010",7465 => "01011100",7466 => "11011101",7467 => "01101000",7468 => "00100000",7469 => "01111100",7470 => "00111000",7471 => "01011110",7472 => "11001110",7473 => "11111011",7474 => "11110110",7475 => "11010011",7476 => "11100000",7477 => "11101111",7478 => "00001010",7479 => "01110010",7480 => "11111100",7481 => "01000001",7482 => "01100101",7483 => "00110111",7484 => "10010111",7485 => "01010010",7486 => "00110011",7487 => "00001011",7488 => "00100010",7489 => "11100111",7490 => "11110101",7491 => "10101100",7492 => "11111011",7493 => "10011011",7494 => "00000000",7495 => "01101101",7496 => "11100111",7497 => "00101101",7498 => "11100111",7499 => "01111000",7500 => "00100010",7501 => "01111101",7502 => "11000011",7503 => "01100110",7504 => "10111111",7505 => "00110000",7506 => "11101100",7507 => "11000010",7508 => "11000110",7509 => "01110100",7510 => "00111011",7511 => "10000100",7512 => "11000000",7513 => "10100110",7514 => "11111001",7515 => "01101110",7516 => "10001001",7517 => "01110000",7518 => "01110110",7519 => "11100000",7520 => "00000101",7521 => "00100001",7522 => "11010100",7523 => "01101010",7524 => "00101100",7525 => "01011001",7526 => "01000101",7527 => "01001000",7528 => "11110010",7529 => "01100101",7530 => "00000000",7531 => "11101110",7532 => "10010111",7533 => "00010000",7534 => "10101100",7535 => "01101011",7536 => "01100000",7537 => "11111000",7538 => "01011000",7539 => "11101000",7540 => "01100110",7541 => "01111001",7542 => "10011000",7543 => "01111111",7544 => "11001101",7545 => "10011110",7546 => "10110110",7547 => "00100001",7548 => "11000101",7549 => "00010000",7550 => "11100000",7551 => "11010000",7552 => "01000111",7553 => "10010101",7554 => "10000011",7555 => "00101011",7556 => "10010001",7557 => "00100001",7558 => "10110010",7559 => "01010101",7560 => "10000110",7561 => "01011000",7562 => "11011100",7563 => "11110000",7564 => "00111001",7565 => "00001001",7566 => "11000111",7567 => "10010010",7568 => "01000101",7569 => "10001111",7570 => "00101000",7571 => "00100011",7572 => "00000001",7573 => "01110101",7574 => "01001010",7575 => "00010001",7576 => "01000101",7577 => "01011100",7578 => "11011010",7579 => "11110000",7580 => "11001001",7581 => "01011001",7582 => "11100000",7583 => "00001001",7584 => "10000110",7585 => "11111011",7586 => "11000111",7587 => "00100010",7588 => "10011000",7589 => "00100111",7590 => "10010010",7591 => "00110000",7592 => "11001011",7593 => "00011011",7594 => "10010110",7595 => "01111101",7596 => "11010110",7597 => "00010111",7598 => "11011100",7599 => "01000111",7600 => "01101111",7601 => "10000001",7602 => "10001011",7603 => "11110101",7604 => "00011100",7605 => "00110011",7606 => "00110000",7607 => "01101100",7608 => "00110011",7609 => "00001010",7610 => "10000010",7611 => "11110010",7612 => "01101110",7613 => "01101010",7614 => "11010101",7615 => "01110100",7616 => "10110110",7617 => "10100011",7618 => "01111001",7619 => "00101101",7620 => "10000000",7621 => "01000000",7622 => "00001011",7623 => "10010010",7624 => "11010111",7625 => "10111110",7626 => "10010000",7627 => "00000110",7628 => "00110100",7629 => "01101101",7630 => "10110010",7631 => "00111111",7632 => "11000100",7633 => "00000000",7634 => "00010101",7635 => "00011011",7636 => "10000010",7637 => "00101001",7638 => "00100101",7639 => "11000011",7640 => "00110010",7641 => "00010011",7642 => "01100111",7643 => "11011111",7644 => "00000110",7645 => "00110100",7646 => "00100111",7647 => "11010111",7648 => "01000110",7649 => "11100111",7650 => "10011100",7651 => "00100001",7652 => "01100001",7653 => "01001000",7654 => "10000000",7655 => "01100000",7656 => "00110111",7657 => "10111001",7658 => "01100111",7659 => "01000110",7660 => "11100110",7661 => "10101000",7662 => "11011001",7663 => "01110010",7664 => "01111101",7665 => "10001010",7666 => "10000101",7667 => "10001000",7668 => "10110110",7669 => "11110001",7670 => "01110011",7671 => "11111011",7672 => "10000111",7673 => "01101001",7674 => "00101110",7675 => "11011011",7676 => "10011111",7677 => "01010111",7678 => "00100101",7679 => "01111111",7680 => "10001000",7681 => "00000000",7682 => "00101001",7683 => "01011010",7684 => "11011111",7685 => "10010011",7686 => "01011101",7687 => "10100010",7688 => "10011001",7689 => "00010011",7690 => "10010001",7691 => "01100000",7692 => "10000000",7693 => "01100110",7694 => "10111010",7695 => "10011100",7696 => "11010000",7697 => "10101001",7698 => "10111000",7699 => "11011011",7700 => "01110101",7701 => "00100001",7702 => "01111100",7703 => "11100100",7704 => "00010101",7705 => "11011110",7706 => "01111010",7707 => "10011101",7708 => "11101110",7709 => "01110101",7710 => "00101001",7711 => "10001100",7712 => "00100100",7713 => "11101001",7714 => "00000110",7715 => "10011110",7716 => "00000000",7717 => "11101001",7718 => "11011010",7719 => "00000001",7720 => "00101010",7721 => "10010001",7722 => "11001110",7723 => "11011000",7724 => "01000111",7725 => "10010010",7726 => "01010111",7727 => "01000100",7728 => "00001111",7729 => "10010110",7730 => "11010111",7731 => "00001111",7732 => "01001001",7733 => "11011101",7734 => "11101000",7735 => "11101111",7736 => "00001100",7737 => "11100111",7738 => "10001111",7739 => "00110110",7740 => "00111100",7741 => "00010101",7742 => "11000000",7743 => "11010010",7744 => "00101010",7745 => "11011000",7746 => "10110010",7747 => "11010100",7748 => "00000011",7749 => "01010001",7750 => "00000001",7751 => "00000111",7752 => "11111100",7753 => "10001001",7754 => "11001111",7755 => "01001111",7756 => "01101100",7757 => "01011100",7758 => "01110001",7759 => "00100110",7760 => "01110011",7761 => "10011100",7762 => "01010110",7763 => "10010110",7764 => "10100011",7765 => "00110010",7766 => "00101101",7767 => "01001011",7768 => "01011101",7769 => "10100001",7770 => "01000101",7771 => "10100000",7772 => "00010111",7773 => "11011000",7774 => "10101100",7775 => "00111011",7776 => "01101100",7777 => "00100011",7778 => "11111011",7779 => "10000110",7780 => "01101100",7781 => "10011011",7782 => "11111111",7783 => "10110111",7784 => "11101101",7785 => "00111100",7786 => "01110000",7787 => "00111001",7788 => "01101001",7789 => "01111101",7790 => "10111110",7791 => "10000100",7792 => "11101001",7793 => "01001010",7794 => "01101010",7795 => "11001011",7796 => "10101001",7797 => "10101001",7798 => "10101001",7799 => "01010100",7800 => "10110110",7801 => "10010110",7802 => "11001000",7803 => "01011010",7804 => "10011110",7805 => "00101101",7806 => "11000110",7807 => "00011100",7808 => "01110000",7809 => "00101101",7810 => "10011111",7811 => "11110111",7812 => "00010111",7813 => "00000001",7814 => "00110011",7815 => "01100100",7816 => "11110000",7817 => "10001110",7818 => "00001100",7819 => "10110000",7820 => "01111000",7821 => "00101101",7822 => "11010111",7823 => "11101000",7824 => "10000001",7825 => "00000110",7826 => "01110011",7827 => "01101110",7828 => "10010110",7829 => "00010001",7830 => "10000111",7831 => "00001001",7832 => "01111110",7833 => "01000101",7834 => "00100011",7835 => "01111110",7836 => "11111110",7837 => "10011111",7838 => "11111100",7839 => "10101001",7840 => "01111110",7841 => "11100010",7842 => "10011110",7843 => "10100100",7844 => "10001110",7845 => "01101001",7846 => "10011001",7847 => "00001101",7848 => "00001010",7849 => "11001111",7850 => "00111001",7851 => "00110111",7852 => "00000011",7853 => "10111110",7854 => "00110011",7855 => "11010101",7856 => "10100000",7857 => "00110010",7858 => "11011101",7859 => "11100100",7860 => "11011000",7861 => "01110001",7862 => "10111011",7863 => "01011001",7864 => "00000010",7865 => "00000111",7866 => "00000110",7867 => "10100101",7868 => "11111110",7869 => "11101100",7870 => "00001110",7871 => "10000110",7872 => "01100101",7873 => "01010011",7874 => "10100001",7875 => "11110100",7876 => "11110010",7877 => "01011110",7878 => "11001111",7879 => "01111010",7880 => "11110001",7881 => "11110111",7882 => "11100000",7883 => "11010000",7884 => "11011101",7885 => "00101011",7886 => "11110111",7887 => "00010101",7888 => "01100001",7889 => "00010011",7890 => "11100111",7891 => "10110100",7892 => "11101001",7893 => "11010011",7894 => "01001011",7895 => "10000011",7896 => "01000110",7897 => "01100000",7898 => "00101110",7899 => "01100101",7900 => "11001111",7901 => "10000101",7902 => "00000001",7903 => "10010000",7904 => "10111001",7905 => "01111000",7906 => "01111110",7907 => "11111111",7908 => "01010011",7909 => "10000100",7910 => "10100110",7911 => "01110101",7912 => "11100010",7913 => "11010101",7914 => "11110000",7915 => "00001010",7916 => "00111111",7917 => "00111100",7918 => "10101110",7919 => "00011101",7920 => "01001011",7921 => "01011001",7922 => "10010010",7923 => "01000011",7924 => "10011100",7925 => "01011100",7926 => "01011010",7927 => "11010110",7928 => "11001001",7929 => "00110000",7930 => "01111111",7931 => "10111011",7932 => "00110111",7933 => "01011110",7934 => "00010101",7935 => "11100111",7936 => "00100101",7937 => "00100001",7938 => "01100001",7939 => "00101010",7940 => "01111010",7941 => "10100000",7942 => "00010110",7943 => "11101001",7944 => "11110101",7945 => "11001110",7946 => "01100111",7947 => "01001011",7948 => "01001011",7949 => "11010100",7950 => "10011000",7951 => "11100110",7952 => "00110011",7953 => "01000111",7954 => "11001000",7955 => "00111000",7956 => "10011011",7957 => "11011000",7958 => "01011000",7959 => "00101010",7960 => "00100110",7961 => "10011101",7962 => "00100000",7963 => "00100111",7964 => "11011101",7965 => "00010010",7966 => "00101000",7967 => "10111010",7968 => "10111100",7969 => "01001101",7970 => "11010000",7971 => "11001101",7972 => "11001010",7973 => "11011100",7974 => "11011101",7975 => "10111010",7976 => "11010000",7977 => "11110100",7978 => "10010011",7979 => "11110101",7980 => "01000111",7981 => "00110100",7982 => "01000100",7983 => "11110100",7984 => "10001001",7985 => "01110101",7986 => "00101110",7987 => "11001000",7988 => "01110010",7989 => "10000101",7990 => "00000010",7991 => "00100101",7992 => "01111011",7993 => "11001001",7994 => "10111011",7995 => "00100001",7996 => "01111110",7997 => "11110101",7998 => "00000101",7999 => "01100010",8000 => "00101001",8001 => "10100101",8002 => "10111000",8003 => "01001101",8004 => "10001101",8005 => "00110001",8006 => "01100010",8007 => "10110110",8008 => "01101010",8009 => "00100111",8010 => "01011110",8011 => "01100110",8012 => "01001011",8013 => "00001110",8014 => "10101101",8015 => "01111111",8016 => "01110001",8017 => "11000111",8018 => "00110111",8019 => "10000101",8020 => "01100100",8021 => "01100001",8022 => "01001101",8023 => "00110011",8024 => "01101010",8025 => "01101100",8026 => "10010110",8027 => "00110011",8028 => "01101010",8029 => "00111001",8030 => "11001001",8031 => "01111010",8032 => "10101100",8033 => "00101110",8034 => "01001011",8035 => "11101110",8036 => "11000110",8037 => "01010001",8038 => "11100110",8039 => "10000101",8040 => "00100001",8041 => "00001110",8042 => "01110111",8043 => "00010110",8044 => "11101100",8045 => "01111111",8046 => "01110010",8047 => "11001000",8048 => "01110111",8049 => "01011110",8050 => "11010100",8051 => "10000110",8052 => "00011011",8053 => "11110100",8054 => "11001110",8055 => "11100111",8056 => "10100001",8057 => "00100000",8058 => "01101011",8059 => "11010111",8060 => "00110101",8061 => "01100110",8062 => "11101001",8063 => "10001011",8064 => "11010001",8065 => "11111110",8066 => "01000111",8067 => "10110110",8068 => "00111100",8069 => "10001000",8070 => "10000101",8071 => "10110100",8072 => "01010101",8073 => "10101101",8074 => "11101101",8075 => "01101110",8076 => "11011000",8077 => "01011011",8078 => "00011010",8079 => "01010110",8080 => "10110010",8081 => "10100011",8082 => "10011110",8083 => "01110110",8084 => "10100111",8085 => "10010000",8086 => "10100111",8087 => "11110011",8088 => "11111101",8089 => "01110100",8090 => "01010111",8091 => "11001111",8092 => "00100101",8093 => "01001011",8094 => "10100110",8095 => "10110000",8096 => "11110000",8097 => "10011011",8098 => "10111111",8099 => "11011000",8100 => "11010000",8101 => "01000110",8102 => "11101000",8103 => "10011100",8104 => "10110001",8105 => "10000100",8106 => "11010001",8107 => "11000111",8108 => "01000010",8109 => "10000111",8110 => "00110100",8111 => "00110110",8112 => "11110000",8113 => "10100110",8114 => "10110010",8115 => "00000100",8116 => "01110111",8117 => "10111011",8118 => "01001101",8119 => "10000110",8120 => "11010100",8121 => "10010000",8122 => "00110110",8123 => "00010000",8124 => "11110110",8125 => "10001001",8126 => "10011001",8127 => "11111010",8128 => "10000011",8129 => "00100110",8130 => "01101000",8131 => "10001010",8132 => "10110101",8133 => "00010111",8134 => "10000000",8135 => "10011101",8136 => "10110001",8137 => "01011001",8138 => "10000010",8139 => "01111010",8140 => "00010001",8141 => "10000111",8142 => "01111110",8143 => "00100100",8144 => "11110111",8145 => "10110000",8146 => "01000011",8147 => "01101100",8148 => "10001000",8149 => "01001001",8150 => "00000111",8151 => "01011000",8152 => "11100101",8153 => "01010111",8154 => "11100101",8155 => "01001101",8156 => "10000100",8157 => "11100010",8158 => "11111010",8159 => "11011100",8160 => "00011011",8161 => "11101011",8162 => "01101100",8163 => "01010111",8164 => "10100011",8165 => "10011111",8166 => "10101110",8167 => "00111100",8168 => "01110101",8169 => "01001110",8170 => "01110110",8171 => "10011001",8172 => "01011110",8173 => "10100001",8174 => "10010100",8175 => "00001000",8176 => "11111000",8177 => "10110000",8178 => "11001111",8179 => "01100100",8180 => "01101101",8181 => "01100001",8182 => "10010100",8183 => "01100110",8184 => "01001101",8185 => "00001000",8186 => "10101100",8187 => "01010000",8188 => "10001111",8189 => "00000001",8190 => "11101011",8191 => "10111011",8192 => "01100010",8193 => "00110001",8194 => "11100000",8195 => "00110100",8196 => "01111110",8197 => "00100111",8198 => "00110100",8199 => "11000100",8200 => "01010000",8201 => "11011011",8202 => "01001010",8203 => "00110101",8204 => "10100100",8205 => "11111010",8206 => "11100101",8207 => "00000101",8208 => "01011010",8209 => "11101000",8210 => "11110110",8211 => "00100000",8212 => "11001111",8213 => "11100010",8214 => "00010100",8215 => "10001100",8216 => "01010001",8217 => "10111000",8218 => "10000101",8219 => "10110101",8220 => "00000100",8221 => "01111111",8222 => "00110001",8223 => "01101111",8224 => "11111011",8225 => "01101101",8226 => "11100011",8227 => "11000100",8228 => "10100011",8229 => "01100011",8230 => "01011001",8231 => "11001000",8232 => "10011110",8233 => "00010000",8234 => "11110100",8235 => "00101010",8236 => "00100011",8237 => "10100111",8238 => "01000001",8239 => "00011000",8240 => "11100111",8241 => "10110111",8242 => "01010001",8243 => "11111010",8244 => "00101001",8245 => "10010000",8246 => "11001100",8247 => "10101011",8248 => "11000101",8249 => "10111011",8250 => "01111111",8251 => "00011001",8252 => "01110010",8253 => "11011110",8254 => "11000001",8255 => "10011000",8256 => "01110001",8257 => "10101011",8258 => "00100010",8259 => "01100110",8260 => "00011110",8261 => "01101011",8262 => "10000100",8263 => "10110101",8264 => "00110111",8265 => "11001110",8266 => "00110001",8267 => "01001100",8268 => "10101001",8269 => "01100111",8270 => "10101010",8271 => "11101010",8272 => "10010000",8273 => "01010101",8274 => "10100010",8275 => "10110101",8276 => "00100100",8277 => "00100100",8278 => "11011101",8279 => "11111000",8280 => "00010110",8281 => "00111010",8282 => "00000000",8283 => "10011000",8284 => "11010000",8285 => "01100101",8286 => "10011100",8287 => "11100010",8288 => "01110110",8289 => "11001011",8290 => "10011011",8291 => "00100100",8292 => "01001101",8293 => "01110010",8294 => "11100000",8295 => "10010001",8296 => "10111010",8297 => "01100001",8298 => "01001110",8299 => "10000100",8300 => "01011011",8301 => "00011110",8302 => "11100111",8303 => "01000111",8304 => "11100101",8305 => "00110001",8306 => "11010011",8307 => "00101000",8308 => "00111111",8309 => "00010110",8310 => "00001011",8311 => "11110000",8312 => "01101110",8313 => "11001011",8314 => "01011110",8315 => "00100001",8316 => "00001000",8317 => "01101111",8318 => "01111100",8319 => "01001111",8320 => "11000111",8321 => "00101111",8322 => "01111001",8323 => "01011110",8324 => "00000000",8325 => "10000001",8326 => "01011001",8327 => "10110011",8328 => "11010101",8329 => "10000011",8330 => "11011101",8331 => "00011000",8332 => "01101000",8333 => "11011101",8334 => "10110011",8335 => "01010110",8336 => "11001101",8337 => "11111011",8338 => "10011110",8339 => "00101100",8340 => "01011110",8341 => "00001101",8342 => "01101101",8343 => "01010001",8344 => "11111001",8345 => "00100001",8346 => "00100010",8347 => "01000110",8348 => "10001101",8349 => "10111110",8350 => "01100110",8351 => "01000101",8352 => "11011010",8353 => "00000100",8354 => "10101010",8355 => "00000010",8356 => "00101110",8357 => "10111100",8358 => "10110000",8359 => "10101010",8360 => "10000101",8361 => "11000101",8362 => "00110010",8363 => "11011101",8364 => "00001011",8365 => "01000011",8366 => "11111111",8367 => "01111101",8368 => "11001001",8369 => "00010101",8370 => "11111001",8371 => "00101110",8372 => "10011001",8373 => "01011001",8374 => "11111110",8375 => "00000011",8376 => "00000010",8377 => "00000000",8378 => "11100001",8379 => "01100000",8380 => "11110001",8381 => "10111110",8382 => "01011011",8383 => "10110000",8384 => "00010010",8385 => "01001011",8386 => "10011011",8387 => "10100100",8388 => "01100010",8389 => "11101100",8390 => "10110010",8391 => "00001110",8392 => "01011001",8393 => "11010100",8394 => "00111101",8395 => "10000101",8396 => "10010111",8397 => "10110100",8398 => "00010010",8399 => "01111011",8400 => "10011110",8401 => "00001110",8402 => "01000110",8403 => "01111000",8404 => "00000110",8405 => "10101101",8406 => "01010000",8407 => "01101101",8408 => "00110110",8409 => "01000111",8410 => "01111001",8411 => "01000110",8412 => "00111111",8413 => "00010001",8414 => "00010101",8415 => "00100111",8416 => "11011111",8417 => "11101000",8418 => "00011100",8419 => "01001000",8420 => "11000010",8421 => "01001100",8422 => "01000000",8423 => "01001110",8424 => "11011100",8425 => "10101110",8426 => "10111011",8427 => "10001101",8428 => "00001011",8429 => "00010111",8430 => "00111101",8431 => "01001110",8432 => "10100111",8433 => "10101101",8434 => "01010010",8435 => "00010010",8436 => "00010100",8437 => "00000010",8438 => "00000111",8439 => "11001110",8440 => "00101110",8441 => "10001001",8442 => "11010001",8443 => "10100111",8444 => "11100011",8445 => "10110000",8446 => "00101110",8447 => "11000100",8448 => "10110110",8449 => "01101010",8450 => "00011010",8451 => "11110111",8452 => "10100101",8453 => "11110111",8454 => "10110011",8455 => "11100011",8456 => "00101001",8457 => "11000110",8458 => "11110101",8459 => "10011011",8460 => "11011101",8461 => "10100011",8462 => "10001010",8463 => "11101101",8464 => "00000000",8465 => "00011010",8466 => "11111111",8467 => "01000100",8468 => "00000011",8469 => "11101011",8470 => "01100100",8471 => "00000000",8472 => "01001001",8473 => "00110111",8474 => "10101010",8475 => "00011110",8476 => "01000001",8477 => "01111110",8478 => "11101001",8479 => "00001000",8480 => "11100000",8481 => "00101011",8482 => "10101001",8483 => "10001101",8484 => "11110111",8485 => "01001100",8486 => "01000000",8487 => "01000111",8488 => "00111000",8489 => "10101000",8490 => "10011111",8491 => "01101011",8492 => "00011000",8493 => "10011100",8494 => "10011111",8495 => "00100010",8496 => "01001001",8497 => "01011010",8498 => "00101100",8499 => "11101100",8500 => "11001000",8501 => "11111001",8502 => "00001110",8503 => "10100100",8504 => "01001100",8505 => "11111100",8506 => "00110110",8507 => "00010100",8508 => "11101100",8509 => "10010010",8510 => "00111010",8511 => "10100110",8512 => "01101001",8513 => "10111001",8514 => "01010010",8515 => "10111000",8516 => "00110011",8517 => "10100000",8518 => "10101001",8519 => "11100011",8520 => "11000101",8521 => "01100010",8522 => "01101000",8523 => "11100010",8524 => "10100000",8525 => "01110100",8526 => "00110101",8527 => "10001111",8528 => "11101111",8529 => "11100100",8530 => "10010100",8531 => "01101100",8532 => "01011111",8533 => "10000010",8534 => "01000010",8535 => "11001011",8536 => "00001101",8537 => "10100111",8538 => "11101010",8539 => "01101111",8540 => "10001000",8541 => "01010111",8542 => "00111110",8543 => "11100110",8544 => "11010111",8545 => "01000011",8546 => "10100001",8547 => "11001010",8548 => "01100001",8549 => "01111010",8550 => "11111100",8551 => "01011011",8552 => "00011101",8553 => "11011100",8554 => "01100001",8555 => "01000110",8556 => "11101001",8557 => "10000011",8558 => "01100000",8559 => "11000111",8560 => "00110000",8561 => "01100000",8562 => "11111100",8563 => "10010001",8564 => "01000101",8565 => "11101101",8566 => "10111010",8567 => "00110001",8568 => "01011000",8569 => "11001011",8570 => "00100001",8571 => "10111011",8572 => "11001100",8573 => "00111111",8574 => "11110101",8575 => "10111000",8576 => "01000010",8577 => "11011110",8578 => "10111011",8579 => "01110101",8580 => "10111010",8581 => "11110010",8582 => "00111011",8583 => "10110110",8584 => "00010100",8585 => "01010100",8586 => "01010100",8587 => "11101101",8588 => "11001001",8589 => "10011010",8590 => "00000010",8591 => "11010011",8592 => "01010000",8593 => "01010101",8594 => "01100000",8595 => "11110000",8596 => "01011101",8597 => "11011001",8598 => "00101100",8599 => "11010000",8600 => "00111001",8601 => "10101100",8602 => "00010101",8603 => "00000010",8604 => "00100100",8605 => "00111011",8606 => "01110001",8607 => "01011101",8608 => "01101111",8609 => "01001110",8610 => "01001111",8611 => "10101011",8612 => "11000111",8613 => "00010011",8614 => "11101100",8615 => "01111110",8616 => "00101111",8617 => "01101000",8618 => "10110001",8619 => "00001011",8620 => "11100101",8621 => "01111011",8622 => "00111010",8623 => "01010101",8624 => "00111000",8625 => "11101011",8626 => "10000001",8627 => "01100010",8628 => "10100110",8629 => "10011011",8630 => "10011011",8631 => "10100101",8632 => "01001001",8633 => "11000100",8634 => "11101001",8635 => "00101101",8636 => "01000110",8637 => "01010101",8638 => "11110010",8639 => "00000100",8640 => "01110011",8641 => "01001010",8642 => "11101001",8643 => "10001010",8644 => "10100001",8645 => "00010111",8646 => "01110000",8647 => "10110010",8648 => "00111001",8649 => "00010101",8650 => "10101110",8651 => "11110111",8652 => "10101001",8653 => "11111000",8654 => "01001101",8655 => "01000100",8656 => "11111111",8657 => "11011110",8658 => "11101000",8659 => "00100100",8660 => "01100000",8661 => "01000111",8662 => "00101011",8663 => "10000100",8664 => "00011011",8665 => "11001101",8666 => "11110111",8667 => "10000110",8668 => "01001011",8669 => "10000111",8670 => "10101010",8671 => "10000101",8672 => "11011011",8673 => "11110111",8674 => "01110100",8675 => "11110000",8676 => "01111101",8677 => "01010100",8678 => "10000100",8679 => "01101001",8680 => "10101100",8681 => "01110100",8682 => "00100011",8683 => "01000101",8684 => "01110110",8685 => "01101011",8686 => "01100000",8687 => "00100000",8688 => "00100111",8689 => "00001110",8690 => "00111010",8691 => "10010100",8692 => "11010001",8693 => "01101000",8694 => "00001110",8695 => "11010110",8696 => "11101011",8697 => "11110111",8698 => "10000111",8699 => "10110100",8700 => "00111011",8701 => "11000100",8702 => "00110001",8703 => "00110001",8704 => "00000101",8705 => "11101110",8706 => "10111011",8707 => "00110000",8708 => "11110100",8709 => "11001011",8710 => "11011110",8711 => "10100001",8712 => "10010100",8713 => "10101010",8714 => "00101010",8715 => "01010001",8716 => "11000000",8717 => "10001100",8718 => "00011101",8719 => "01111111",8720 => "01001111",8721 => "11010101",8722 => "01110111",8723 => "01110100",8724 => "11101101",8725 => "01011010",8726 => "01010001",8727 => "11011010",8728 => "11000011",8729 => "10111110",8730 => "01011011",8731 => "00101011",8732 => "11011011",8733 => "00110100",8734 => "01001101",8735 => "00010100",8736 => "11100010",8737 => "01101111",8738 => "11110100",8739 => "11110111",8740 => "10001100",8741 => "01101000",8742 => "00101011",8743 => "00011110",8744 => "01110111",8745 => "10000000",8746 => "11000011",8747 => "11001011",8748 => "01100010",8749 => "11110011",8750 => "01110111",8751 => "10101111",8752 => "01001000",8753 => "10100001",8754 => "10000101",8755 => "00110101",8756 => "00000011",8757 => "11001111",8758 => "00011001",8759 => "10101110",8760 => "10111010",8761 => "10010101",8762 => "01010001",8763 => "11001111",8764 => "11001001",8765 => "10111001",8766 => "00101011",8767 => "10100010",8768 => "10100110",8769 => "10000101",8770 => "00111101",8771 => "10011001",8772 => "11101101",8773 => "10101111",8774 => "11001001",8775 => "10001111",8776 => "00011000",8777 => "00010100",8778 => "00011100",8779 => "01011111",8780 => "11111010",8781 => "10011111",8782 => "10100110",8783 => "01010001",8784 => "01011000",8785 => "00101110",8786 => "11101110",8787 => "01111111",8788 => "01111001",8789 => "00100100",8790 => "00000110",8791 => "01000111",8792 => "10111011",8793 => "00111111",8794 => "01101001",8795 => "00101000",8796 => "01110110",8797 => "00011101",8798 => "10101111",8799 => "01110100",8800 => "10000110",8801 => "11000100",8802 => "11011111",8803 => "11110000",8804 => "01010010",8805 => "01011110",8806 => "11001111",8807 => "00010011",8808 => "00100011",8809 => "10000100",8810 => "00101000",8811 => "01001001",8812 => "10001100",8813 => "01111010",8814 => "00111000",8815 => "01111001",8816 => "10001011",8817 => "01101001",8818 => "10100001",8819 => "11110110",8820 => "11010001",8821 => "01100101",8822 => "00110111",8823 => "00110010",8824 => "01010000",8825 => "00111111",8826 => "11010100",8827 => "10101111",8828 => "01101110",8829 => "10000010",8830 => "01111101",8831 => "11010111",8832 => "00111101",8833 => "11010101",8834 => "01100100",8835 => "01110011",8836 => "10111101",8837 => "11101100",8838 => "10101101",8839 => "00000000",8840 => "01100011",8841 => "01001000",8842 => "10101011",8843 => "00101001",8844 => "00110110",8845 => "01011110",8846 => "10000001",8847 => "01101100",8848 => "00100001",8849 => "10001101",8850 => "00101111",8851 => "01011101",8852 => "11010101",8853 => "01011000",8854 => "00001101",8855 => "00100110",8856 => "00101001",8857 => "01100000",8858 => "10111000",8859 => "00011011",8860 => "00110011",8861 => "11101010",8862 => "10000110",8863 => "11100010",8864 => "01100111",8865 => "00001100",8866 => "11111101",8867 => "10011010",8868 => "00100100",8869 => "11001100",8870 => "11010111",8871 => "01000011",8872 => "00010011",8873 => "01100110",8874 => "10101100",8875 => "00111110",8876 => "11001000",8877 => "01001001",8878 => "00010100",8879 => "10000110",8880 => "01101110",8881 => "11011001",8882 => "01100011",8883 => "11111101",8884 => "01001110",8885 => "11000110",8886 => "01111000",8887 => "01100001",8888 => "10100101",8889 => "11001101",8890 => "01100110",8891 => "00111011",8892 => "11000101",8893 => "01101000",8894 => "10101100",8895 => "11000111",8896 => "11101001",8897 => "00111111",8898 => "01000111",8899 => "11011001",8900 => "00100011",8901 => "11100101",8902 => "10000001",8903 => "01010010",8904 => "01000001",8905 => "11100010",8906 => "11001111",8907 => "11001100",8908 => "10000000",8909 => "00110111",8910 => "01101101",8911 => "11011010",8912 => "00000100",8913 => "01101101",8914 => "10000010",8915 => "00010101",8916 => "10001000",8917 => "00110001",8918 => "00101011",8919 => "11110010",8920 => "01010000",8921 => "01001100",8922 => "10110010",8923 => "01110011",8924 => "01101001",8925 => "01011101",8926 => "00110111",8927 => "11011111",8928 => "11010100",8929 => "10001101",8930 => "10110111",8931 => "00110100",8932 => "10101100",8933 => "10000110",8934 => "00101001",8935 => "00100111",8936 => "00110101",8937 => "11100110",8938 => "10010101",8939 => "01100000",8940 => "11110100",8941 => "01101110",8942 => "00011100",8943 => "01001100",8944 => "01111110",8945 => "10010000",8946 => "01101100",8947 => "00000101",8948 => "00111001",8949 => "10011100",8950 => "11001101",8951 => "10100111",8952 => "10000001",8953 => "10111010",8954 => "00011010",8955 => "00001010",8956 => "00111011",8957 => "11110000",8958 => "10011000",8959 => "11110110",8960 => "10100100",8961 => "01100010",8962 => "01100110",8963 => "11110000",8964 => "00100101",8965 => "01100111",8966 => "01011010",8967 => "11100110",8968 => "11101110",8969 => "00010100",8970 => "00001010",8971 => "11110100",8972 => "01111010",8973 => "11011111",8974 => "11011010",8975 => "11011100",8976 => "00011111",8977 => "01110011",8978 => "10010001",8979 => "11010011",8980 => "11000111",8981 => "01000100",8982 => "01011100",8983 => "10111110",8984 => "11000110",8985 => "11100101",8986 => "01110011",8987 => "00001001",8988 => "11000010",8989 => "01010000",8990 => "00001010",8991 => "00001110",8992 => "11000000",8993 => "11111001",8994 => "00101000",8995 => "11110101",8996 => "01001110",8997 => "11101110",8998 => "01001010",8999 => "10011011",9000 => "11110100",9001 => "11111110",9002 => "01101101",9003 => "10000101",9004 => "00001010",9005 => "10100010",9006 => "01011011",9007 => "01001110",9008 => "01111010",9009 => "10101101",9010 => "11111111",9011 => "00110011",9012 => "10001111",9013 => "01011101",9014 => "00011101",9015 => "11110110",9016 => "00011100",9017 => "11110111",9018 => "11100000",9019 => "11010110",9020 => "00111111",9021 => "01100000",9022 => "01010110",9023 => "10000111",9024 => "10001100",9025 => "01111011",9026 => "01011110",9027 => "00110000",9028 => "10011100",9029 => "10100100",9030 => "11010101",9031 => "10010111",9032 => "11011010",9033 => "10010110",9034 => "01100100",9035 => "11010110",9036 => "11001011",9037 => "00010001",9038 => "01010010",9039 => "00001001",9040 => "00001010",9041 => "11000101",9042 => "01000000",9043 => "11111111",9044 => "01101101",9045 => "10111100",9046 => "11101011",9047 => "11010100",9048 => "10010101",9049 => "10011110",9050 => "11111000",9051 => "00100000",9052 => "10101110",9053 => "01111111",9054 => "11001110",9055 => "01100101",9056 => "01000010",9057 => "11000111",9058 => "10101111",9059 => "01011000",9060 => "10101111",9061 => "01111000",9062 => "01011101",9063 => "11100100",9064 => "00000011",9065 => "01110110",9066 => "11010011",9067 => "10111110",9068 => "01011011",9069 => "10011110",9070 => "11101111",9071 => "01011010",9072 => "01101001",9073 => "00000010",9074 => "10110011",9075 => "01101101",9076 => "00100000",9077 => "11100001",9078 => "11001001",9079 => "10000111",9080 => "00110011",9081 => "11010100",9082 => "11001110",9083 => "10001101",9084 => "00110010",9085 => "10100000",9086 => "00001001",9087 => "00101101",9088 => "11000011",9089 => "11111001",9090 => "10111000",9091 => "10101011",9092 => "00001100",9093 => "00101011",9094 => "01110110",9095 => "10100001",9096 => "10010111",9097 => "01000011",9098 => "11000010",9099 => "01011111",9100 => "10011100",9101 => "11001110",9102 => "10100010",9103 => "01000111",9104 => "10010111",9105 => "10111111",9106 => "01001111",9107 => "10001001",9108 => "01101101",9109 => "10000011",9110 => "10111111",9111 => "01001110",9112 => "10110010",9113 => "11110001",9114 => "01101011",9115 => "11011001",9116 => "11001010",9117 => "11100000",9118 => "01110100",9119 => "10011010",9120 => "11101001",9121 => "01100101",9122 => "01011011",9123 => "10110110",9124 => "11100000",9125 => "00101101",9126 => "10001010",9127 => "00111111",9128 => "11001000",9129 => "01100100",9130 => "11101001",9131 => "01011100",9132 => "01011010",9133 => "10111111",9134 => "11110000",9135 => "10101000",9136 => "10010110",9137 => "11011010",9138 => "00110111",9139 => "01001100",9140 => "11100101",9141 => "10011100",9142 => "01101100",9143 => "01111011",9144 => "11101100",9145 => "11110100",9146 => "00000011",9147 => "11000111",9148 => "11111110",9149 => "11100001",9150 => "00101100",9151 => "00110001",9152 => "11010011",9153 => "11111111",9154 => "01010000",9155 => "10110110",9156 => "10111011",9157 => "10011001",9158 => "00010100",9159 => "10011001",9160 => "10110001",9161 => "10101101",9162 => "00001101",9163 => "01001100",9164 => "00001011",9165 => "00011111",9166 => "10000110",9167 => "00101000",9168 => "00110000",9169 => "00111100",9170 => "10010000",9171 => "01111100",9172 => "01110000",9173 => "10101000",9174 => "00100000",9175 => "10101101",9176 => "10010100",9177 => "11010101",9178 => "11000010",9179 => "11110101",9180 => "01000111",9181 => "10000100",9182 => "00100011",9183 => "00110100",9184 => "00111110",9185 => "01011001",9186 => "00111101",9187 => "11110101",9188 => "01110000",9189 => "00100000",9190 => "11000000",9191 => "10110011",9192 => "11010000",9193 => "00000101",9194 => "11001101",9195 => "00110000",9196 => "01111011",9197 => "01100110",9198 => "01100000",9199 => "10011100",9200 => "00100100",9201 => "10100011",9202 => "01111101",9203 => "01110111",9204 => "00100010",9205 => "11001010",9206 => "11010100",9207 => "01010101",9208 => "10101111",9209 => "11100001",9210 => "00100001",9211 => "10010101",9212 => "01101011",9213 => "01000001",9214 => "01000010",9215 => "00101101",9216 => "00101110",9217 => "01100010",9218 => "10000010",9219 => "11001110",9220 => "01000101",9221 => "00111000",9222 => "10001101",9223 => "11101001",9224 => "10010101",9225 => "01010100",9226 => "01100110",9227 => "00111100",9228 => "00110001",9229 => "01000110",9230 => "11101011",9231 => "10101011",9232 => "10001011",9233 => "10011011",9234 => "00110011",9235 => "10010101",9236 => "01011101",9237 => "01001101",9238 => "00100010",9239 => "01000001",9240 => "00011111",9241 => "01111111",9242 => "11111101",9243 => "01001011",9244 => "10001101",9245 => "10100011",9246 => "00011110",9247 => "01001010",9248 => "01100100",9249 => "10100101",9250 => "11110110",9251 => "11111001",9252 => "00001101",9253 => "10111000",9254 => "01100101",9255 => "11011101",9256 => "11001100",9257 => "00100101",9258 => "00100110",9259 => "01100111",9260 => "00001010",9261 => "01001110",9262 => "11000000",9263 => "00000110",9264 => "01101111",9265 => "10110100",9266 => "01100010",9267 => "11111010",9268 => "01011111",9269 => "10011011",9270 => "10110111",9271 => "01010100",9272 => "11011101",9273 => "01000000",9274 => "10011001",9275 => "01000110",9276 => "11100000",9277 => "10001110",9278 => "11001000",9279 => "10101011",9280 => "00111110",9281 => "00100001",9282 => "01001101",9283 => "01111010",9284 => "00111000",9285 => "00001111",9286 => "01110111",9287 => "01111000",9288 => "00011000",9289 => "10011011",9290 => "10101101",9291 => "01010101",9292 => "11000011",9293 => "11100010",9294 => "01011101",9295 => "10100101",9296 => "10111110",9297 => "00001111",9298 => "00011101",9299 => "11000101",9300 => "00111010",9301 => "01100101",9302 => "01100100",9303 => "01001100",9304 => "10010001",9305 => "10111100",9306 => "11110000",9307 => "10111110",9308 => "11011001",9309 => "10001001",9310 => "10000110",9311 => "11110010",9312 => "01101110",9313 => "01101111",9314 => "11101011",9315 => "11111111",9316 => "11110100",9317 => "10110100",9318 => "11010001",9319 => "10111101",9320 => "10101101",9321 => "00110101",9322 => "00000100",9323 => "11000101",9324 => "01100111",9325 => "11101011",9326 => "01010011",9327 => "11101100",9328 => "11110010",9329 => "11110010",9330 => "01111000",9331 => "11111011",9332 => "10111100",9333 => "01110000",9334 => "10001100",9335 => "01110010",9336 => "10101100",9337 => "10001101",9338 => "10001001",9339 => "10100111",9340 => "00011110",9341 => "01110110",9342 => "11101010",9343 => "11000110",9344 => "00010100",9345 => "00110100",9346 => "01010100",9347 => "11111010",9348 => "11001111",9349 => "01001111",9350 => "01011111",9351 => "00010001",9352 => "00001110",9353 => "00011011",9354 => "10110001",9355 => "11001011",9356 => "10110101",9357 => "11111001",9358 => "01111100",9359 => "00001100",9360 => "00101011",9361 => "01011101",9362 => "11000100",9363 => "11110010",9364 => "11100100",9365 => "01011011",9366 => "11010100",9367 => "10001100",9368 => "01100011",9369 => "11111000",9370 => "10110100",9371 => "10101100",9372 => "10001000",9373 => "10110011",9374 => "11100101",9375 => "01110110",9376 => "01110010",9377 => "00111101",9378 => "01101111",9379 => "00010001",9380 => "01000110",9381 => "11010001",9382 => "00110110",9383 => "00110111",9384 => "01111011",9385 => "00110110",9386 => "01011011",9387 => "01100001",9388 => "00101111",9389 => "00101010",9390 => "11001001",9391 => "01111000",9392 => "11100000",9393 => "00010100",9394 => "00110101",9395 => "11010100",9396 => "11100010",9397 => "10101111",9398 => "11100100",9399 => "00111001",9400 => "10000000",9401 => "01010110",9402 => "01101001",9403 => "01101111",9404 => "11011110",9405 => "01000100",9406 => "10101010",9407 => "11001010",9408 => "11100111",9409 => "01010000",9410 => "00011011",9411 => "10110101",9412 => "11100100",9413 => "11110001",9414 => "00010101",9415 => "00001000",9416 => "11111001",9417 => "01000001",9418 => "11010111",9419 => "00001001",9420 => "11011100",9421 => "01111111",9422 => "11001010",9423 => "00111001",9424 => "01011101",9425 => "01111011",9426 => "11010000",9427 => "11100010",9428 => "11000000",9429 => "00111100",9430 => "01111010",9431 => "00000101",9432 => "01001110",9433 => "11010100",9434 => "00111101",9435 => "11011100",9436 => "01001110",9437 => "11110110",9438 => "01110000",9439 => "10111000",9440 => "00001011",9441 => "00100110",9442 => "01110001",9443 => "01101000",9444 => "10011011",9445 => "10100111",9446 => "01001100",9447 => "10111010",9448 => "11011100",9449 => "00110100",9450 => "00011000",9451 => "10001010",9452 => "01111011",9453 => "01101101",9454 => "10011010",9455 => "00011101",9456 => "11011101",9457 => "11010101",9458 => "01100000",9459 => "11100101",9460 => "01110110",9461 => "00011100",9462 => "11111101",9463 => "00011110",9464 => "11100111",9465 => "00110011",9466 => "01011111",9467 => "01101111",9468 => "10011100",9469 => "01101000",9470 => "00110001",9471 => "01000101",9472 => "10110110",9473 => "11101011",9474 => "01010110",9475 => "10101010",9476 => "00011000",9477 => "10110111",9478 => "01110101",9479 => "01010010",9480 => "10001010",9481 => "00001101",9482 => "00011000",9483 => "00110100",9484 => "01001001",9485 => "01110101",9486 => "11101100",9487 => "11100001",9488 => "11100011",9489 => "01101111",9490 => "10011110",9491 => "10100111",9492 => "10110011",9493 => "10001100",9494 => "00110010",9495 => "01000110",9496 => "01010110",9497 => "01101011",9498 => "11110111",9499 => "01010001",9500 => "01111100",9501 => "10101100",9502 => "10111001",9503 => "11000110",9504 => "01100101",9505 => "00000001",9506 => "11101010",9507 => "00000011",9508 => "10000110",9509 => "10011000",9510 => "01010110",9511 => "00001000",9512 => "10000111",9513 => "10011111",9514 => "11000111",9515 => "00100100",9516 => "00000000",9517 => "10000001",9518 => "11010000",9519 => "00000101",9520 => "10001010",9521 => "10001100",9522 => "11101100",9523 => "11001010",9524 => "10110010",9525 => "11111011",9526 => "00110011",9527 => "11100000",9528 => "11010011",9529 => "00110110",9530 => "01010010",9531 => "10101100",9532 => "00011010",9533 => "11100010",9534 => "00101000",9535 => "01111110",9536 => "11101010",9537 => "01110010",9538 => "01011101",9539 => "10000110",9540 => "00011011",9541 => "10010101",9542 => "10010011",9543 => "10010001",9544 => "11111111",9545 => "00110111",9546 => "10101111",9547 => "10000100",9548 => "11111110",9549 => "00101011",9550 => "11011111",9551 => "10110001",9552 => "10011011",9553 => "01010000",9554 => "00101110",9555 => "00100101",9556 => "01110010",9557 => "10010111",9558 => "10101111",9559 => "01001111",9560 => "11011111",9561 => "10000110",9562 => "11000111",9563 => "01100101",9564 => "01111101",9565 => "01110011",9566 => "01111000",9567 => "10010000",9568 => "10011110",9569 => "00000011",9570 => "11000100",9571 => "10010010",9572 => "00101001",9573 => "11111011",9574 => "00110001",9575 => "11001101",9576 => "11000011",9577 => "00000110",9578 => "11100100",9579 => "10101111",9580 => "01101110",9581 => "10110100",9582 => "11100111",9583 => "10011011",9584 => "01011101",9585 => "11110010",9586 => "01111100",9587 => "10000010",9588 => "10110111",9589 => "00010110",9590 => "10101011",9591 => "01101101",9592 => "11011100",9593 => "01111100",9594 => "10000010",9595 => "00111011",9596 => "00101010",9597 => "11111010",9598 => "00011011",9599 => "01010010",9600 => "01111111",9601 => "11011001",9602 => "00101010",9603 => "01100100",9604 => "11010010",9605 => "01001001",9606 => "01011111",9607 => "00000100",9608 => "11011110",9609 => "11101001",9610 => "00001100",9611 => "01001101",9612 => "00101110",9613 => "01111011",9614 => "01101110",9615 => "01010111",9616 => "11000001",9617 => "11100010",9618 => "00110110",9619 => "01011010",9620 => "10001100",9621 => "10011111",9622 => "01001101",9623 => "01011010",9624 => "00011011",9625 => "11011011",9626 => "10100001",9627 => "01000100",9628 => "10111101",9629 => "00101010",9630 => "01111010",9631 => "10010101",9632 => "01110111",9633 => "01110011",9634 => "00010100",9635 => "00100101",9636 => "01100101",9637 => "00101100",9638 => "11110000",9639 => "10000010",9640 => "10110000",9641 => "01110111",9642 => "01011100",9643 => "00010001",9644 => "01100011",9645 => "01001000",9646 => "00011100",9647 => "01110111",9648 => "10100111",9649 => "11100100",9650 => "00010101",9651 => "10101000",9652 => "11000101",9653 => "10000100",9654 => "01000011",9655 => "01110010",9656 => "10100101",9657 => "10101010",9658 => "11001000",9659 => "00011001",9660 => "11110111",9661 => "10110100",9662 => "10000110",9663 => "11100101",9664 => "11000110",9665 => "11111000",9666 => "00111011",9667 => "01001011",9668 => "01110101",9669 => "10101111",9670 => "10001110",9671 => "11111111",9672 => "11110110",9673 => "00100111",9674 => "11001011",9675 => "10110011",9676 => "11100101",9677 => "11010001",9678 => "10100101",9679 => "10101101",9680 => "01101110",9681 => "11011011",9682 => "10111110",9683 => "00111110",9684 => "11100100",9685 => "11001111",9686 => "01011100",9687 => "00101010",9688 => "11011110",9689 => "00111000",9690 => "10011110",9691 => "01000111",9692 => "11011000",9693 => "10011111",9694 => "10100100",9695 => "11011101",9696 => "10000110",9697 => "10001010",9698 => "11101011",9699 => "01100000",9700 => "10011011",9701 => "00010100",9702 => "00111011",9703 => "00110011",9704 => "00101111",9705 => "11101001",9706 => "10011111",9707 => "01000101",9708 => "01101111",9709 => "00000101",9710 => "11000010",9711 => "10110110",9712 => "11101111",9713 => "11101010",9714 => "10100000",9715 => "00111010",9716 => "10110101",9717 => "01010010",9718 => "00011101",9719 => "11100001",9720 => "01100010",9721 => "00100001",9722 => "11111010",9723 => "01101011",9724 => "10001100",9725 => "11100111",9726 => "01011000",9727 => "10010110",9728 => "10000001",9729 => "10000000",9730 => "01111000",9731 => "11110010",9732 => "00011111",9733 => "11010101",9734 => "11110110",9735 => "01110101",9736 => "01001001",9737 => "00111110",9738 => "10110000",9739 => "11000100",9740 => "11110100",9741 => "01000001",9742 => "11011000",9743 => "01100011",9744 => "01011110",9745 => "10001111",9746 => "10110010",9747 => "10101001",9748 => "10101001",9749 => "01001011",9750 => "11000101",9751 => "11111101",9752 => "00100001",9753 => "01010111",9754 => "01101100",9755 => "01111001",9756 => "00110100",9757 => "11001110",9758 => "11000111",9759 => "10100011",9760 => "00111011",9761 => "01001000",9762 => "11110100",9763 => "10011010",9764 => "11001010",9765 => "01110011",9766 => "01110100",9767 => "01101000",9768 => "00110101",9769 => "01101000",9770 => "01110000",9771 => "00011001",9772 => "01101010",9773 => "10101000",9774 => "00011000",9775 => "10101110",9776 => "01011100",9777 => "11111100",9778 => "01111100",9779 => "10000100",9780 => "10010101",9781 => "00001111",9782 => "11110000",9783 => "00011111",9784 => "01000110",9785 => "00010101",9786 => "01110000",9787 => "11101111",9788 => "11011001",9789 => "01001100",9790 => "10101010",9791 => "00101011",9792 => "11010011",9793 => "11100011",9794 => "10100010",9795 => "00011001",9796 => "10011010",9797 => "11000000",9798 => "10111100",9799 => "01101100",9800 => "10101100",9801 => "11011100",9802 => "11010101",9803 => "00100010",9804 => "11100000",9805 => "11001010",9806 => "01011001",9807 => "10110011",9808 => "01000010",9809 => "00110000",9810 => "01001100",9811 => "00111110",9812 => "01101001",9813 => "00101110",9814 => "01001001",9815 => "11000010",9816 => "00100111",9817 => "10101010",9818 => "01101010",9819 => "00001011",9820 => "00011110",9821 => "11000001",9822 => "10110001",9823 => "00100111",9824 => "00000101",9825 => "10100010",9826 => "10111100",9827 => "01011111",9828 => "00001111",9829 => "10000111",9830 => "00001110",9831 => "10010011",9832 => "00100111",9833 => "00000101",9834 => "01100001",9835 => "10101011",9836 => "00110111",9837 => "11110001",9838 => "01100011",9839 => "00011110",9840 => "11111011",9841 => "10101111",9842 => "00111101",9843 => "10010110",9844 => "00011100",9845 => "10110001",9846 => "00110101",9847 => "11110110",9848 => "01100010",9849 => "00110000",9850 => "11110111",9851 => "11000111",9852 => "01100101",9853 => "01101110",9854 => "10000101",9855 => "01010100",9856 => "01000100",9857 => "00000010",9858 => "00001111",9859 => "01010111",9860 => "11100001",9861 => "10001110",9862 => "00110101",9863 => "00110101",9864 => "01110101",9865 => "10001000",9866 => "11101010",9867 => "11011000",9868 => "11011101",9869 => "10111110",9870 => "00011101",9871 => "11100101",9872 => "10101010",9873 => "00001100",9874 => "01100001",9875 => "11010000",9876 => "11111111",9877 => "11111001",9878 => "00111100",9879 => "10011100",9880 => "11011111",9881 => "01110011",9882 => "01001001",9883 => "01111101",9884 => "10011010",9885 => "00000101",9886 => "11111110",9887 => "10101100",9888 => "11001010",9889 => "00110111",9890 => "00011110",9891 => "01001110",9892 => "00111010",9893 => "11101001",9894 => "01110100",9895 => "10101100",9896 => "11011100",9897 => "10011001",9898 => "01000101",9899 => "00001111",9900 => "10110101",9901 => "01101000",9902 => "11111001",9903 => "10000111",9904 => "10100111",9905 => "00111111",9906 => "11100001",9907 => "00100100",9908 => "11010101",9909 => "01100000",9910 => "00001101",9911 => "10111100",9912 => "11111000",9913 => "01101111",9914 => "11111101",9915 => "00100011",9916 => "10110010",9917 => "01111010",9918 => "11110111",9919 => "11100110",9920 => "01111010",9921 => "11001000",9922 => "00010111",9923 => "00111101",9924 => "11011100",9925 => "00011101",9926 => "10111000",9927 => "10111011",9928 => "01011111",9929 => "10011000",9930 => "11111111",9931 => "00101100",9932 => "01001100",9933 => "10001010",9934 => "10110101",9935 => "00111001",9936 => "11101000",9937 => "10001011",9938 => "01100010",9939 => "01000011",9940 => "11001110",9941 => "10011010",9942 => "01101100",9943 => "10111001",9944 => "11001001",9945 => "11011110",9946 => "10110111",9947 => "10000001",9948 => "11001001",9949 => "10010100",9950 => "10111100",9951 => "10100111",9952 => "10011011",9953 => "11110000",9954 => "01100011",9955 => "10000000",9956 => "10101100",9957 => "11111010",9958 => "10010101",9959 => "00001000",9960 => "00011111",9961 => "10101010",9962 => "00000100",9963 => "11111000",9964 => "00001000",9965 => "10100111",9966 => "11000000",9967 => "11100101",9968 => "10110101",9969 => "00111100",9970 => "01001111",9971 => "11001010",9972 => "11010101",9973 => "11011011",9974 => "10011101",9975 => "00110010",9976 => "00000011",9977 => "00010110",9978 => "00101011",9979 => "10000011",9980 => "00101100",9981 => "10101011",9982 => "11000010",9983 => "00010100",9984 => "01101001",9985 => "01101001",9986 => "01110011",9987 => "00010001",9988 => "01111011",9989 => "01111011",9990 => "11011001",9991 => "10101111",9992 => "10111010",9993 => "00011000",9994 => "10110110",9995 => "01010101",9996 => "11000110",9997 => "10100101",9998 => "00011001",9999 => "01000110",10000 => "00010110",10001 => "01001110",10002 => "11011011",10003 => "00011000",10004 => "01111000",10005 => "10101011",10006 => "00011100",10007 => "01100111",10008 => "01010101",10009 => "10000011",10010 => "00011000",10011 => "00011011",10012 => "11010010",10013 => "00111100",10014 => "10001011",10015 => "00000011",10016 => "11101101",10017 => "10111111",10018 => "01101001",10019 => "00000010",10020 => "00111110",10021 => "00101110",10022 => "00010001",10023 => "11001011",10024 => "10110001",10025 => "11001010",10026 => "11010010",10027 => "10000011",10028 => "10101010",10029 => "10101000",10030 => "01100100",10031 => "11001100",10032 => "01000000",10033 => "11011101",10034 => "01100110",10035 => "10111110",10036 => "10000101",10037 => "00111000",10038 => "10010010",10039 => "01100011",10040 => "11011100",10041 => "11011010",10042 => "00000101",10043 => "00000110",10044 => "10100000",10045 => "11010111",10046 => "11010001",10047 => "11010010",10048 => "11101010",10049 => "10101001",10050 => "11010001",10051 => "00111000",10052 => "10010100",10053 => "11011110",10054 => "10111100",10055 => "10110100",10056 => "01001010",10057 => "10011001",10058 => "10111110",10059 => "11110110",10060 => "11110101",10061 => "01011110",10062 => "11100111",10063 => "10001000",10064 => "10000001",10065 => "00001011",10066 => "01000111",10067 => "01011001",10068 => "00100100",10069 => "01111011",10070 => "01011001",10071 => "00111110",10072 => "01000011",10073 => "10001011",10074 => "01000111",10075 => "00011001",10076 => "00011000",10077 => "01100101",10078 => "11001011",10079 => "01111100",10080 => "01000100",10081 => "10111110",10082 => "11010111",10083 => "00100110",10084 => "01011001",10085 => "00001001",10086 => "00011011",10087 => "11101011",10088 => "01001010",10089 => "11110100",10090 => "01010010",10091 => "00011110",10092 => "11111101",10093 => "10000011",10094 => "11110010",10095 => "10110010",10096 => "10110100",10097 => "00010011",10098 => "10111111",10099 => "10100010",10100 => "11011000",10101 => "11110001",10102 => "11101110",10103 => "10101011",10104 => "11101010",10105 => "10000000",10106 => "00000100",10107 => "00111000",10108 => "01010110",10109 => "00001100",10110 => "01110111",10111 => "11000001",10112 => "10111000",10113 => "11111111",10114 => "10001101",10115 => "01111000",10116 => "10011101",10117 => "11000011",10118 => "00110110",10119 => "01001010",10120 => "10010101",10121 => "11000110",10122 => "10000110",10123 => "00111010",10124 => "00111100",10125 => "10011011",10126 => "10010101",10127 => "00011011",10128 => "00101111",10129 => "10101110",10130 => "11110010",10131 => "11100100",10132 => "10110001",10133 => "01000100",10134 => "11000101",10135 => "11011001",10136 => "00111101",10137 => "00001011",10138 => "10000011",10139 => "10101010",10140 => "11101111",10141 => "00001111",10142 => "01101110",10143 => "01000101",10144 => "11110010",10145 => "01110110",10146 => "10111000",10147 => "01100001",10148 => "00101011",10149 => "11011111",10150 => "00101111",10151 => "11010110",10152 => "01000011",10153 => "00100010",10154 => "01100010",10155 => "11100011",10156 => "00011001",10157 => "01010011",10158 => "01101001",10159 => "00101100",10160 => "00100111",10161 => "11100010",10162 => "10010010",10163 => "10000101",10164 => "10000110",10165 => "01111010",10166 => "00011110",10167 => "10101111",10168 => "11010001",10169 => "10010101",10170 => "00011011",10171 => "10110010",10172 => "01000000",10173 => "10001011",10174 => "00111110",10175 => "10010011",10176 => "01101001",10177 => "11101010",10178 => "10101011",10179 => "00100111",10180 => "00101010",10181 => "00011101",10182 => "01100001",10183 => "10011100",10184 => "00101001",10185 => "11000001",10186 => "10100011",10187 => "00010000",10188 => "11101111",10189 => "01101011",10190 => "01111100",10191 => "10101100",10192 => "01001101",10193 => "01110011",10194 => "00101110",10195 => "10010110",10196 => "11010111",10197 => "11100101",10198 => "11001011",10199 => "00100010",10200 => "11010110",10201 => "01110110",10202 => "11001111",10203 => "10010000",10204 => "01111001",10205 => "11111110",10206 => "00010000",10207 => "11111101",10208 => "01011111",10209 => "11000010",10210 => "01010111",10211 => "11011011",10212 => "00000001",10213 => "10100111",10214 => "00111000",10215 => "00100111",10216 => "00111101",10217 => "00110010",10218 => "10001111",10219 => "10011011",10220 => "00111101",10221 => "00010000",10222 => "11010000",10223 => "01001010",10224 => "01111111",10225 => "10100011",10226 => "10011001",10227 => "00011011",10228 => "10000110",10229 => "00111001",10230 => "01000100",10231 => "11010111",10232 => "00110110",10233 => "01011001",10234 => "00010001",10235 => "11000100",10236 => "00010001",10237 => "11111110",10238 => "11101010",10239 => "11111001",10240 => "01101101",10241 => "11000101",10242 => "00100100",10243 => "11101011",10244 => "01001010",10245 => "11000010",10246 => "00011001",10247 => "01011110",10248 => "01011001",10249 => "11101000",10250 => "00000011",10251 => "11101101",10252 => "11101011",10253 => "10001001",10254 => "01111111",10255 => "10101010",10256 => "01110010",10257 => "11011001",10258 => "00110000",10259 => "11001100",10260 => "10000000",10261 => "11101110",10262 => "10110111",10263 => "00100011",10264 => "00110110",10265 => "00000010",10266 => "10101000",10267 => "11110011",10268 => "01001110",10269 => "11011110",10270 => "10001000",10271 => "00101011",10272 => "00001110",10273 => "00001001",10274 => "01011100",10275 => "01101111",10276 => "11111001",10277 => "11010101",10278 => "01010111",10279 => "10011000",10280 => "10101000",10281 => "11110111",10282 => "01011110",10283 => "01110111",10284 => "11011110",10285 => "11011101",10286 => "00100001",10287 => "00010111",10288 => "01110110",10289 => "01010111",10290 => "10001101",10291 => "01011101",10292 => "00111000",10293 => "10100010",10294 => "10100011",10295 => "01001011",10296 => "11001000",10297 => "11111000",10298 => "11101001",10299 => "10000101",10300 => "00111101",10301 => "11111001",10302 => "01110101",10303 => "01000001",10304 => "10110110",10305 => "01011010",10306 => "01101100",10307 => "01000000",10308 => "10100010",10309 => "10111111",10310 => "10111100",10311 => "00111100",10312 => "00100000",10313 => "11101001",10314 => "11111100",10315 => "00000101",10316 => "11000000",10317 => "01101110",10318 => "10010001",10319 => "10000111",10320 => "11110000",10321 => "01100001",10322 => "10101110",10323 => "11011010",10324 => "11110100",10325 => "10000100",10326 => "10111011",10327 => "10110010",10328 => "01101101",10329 => "11110101",10330 => "11001110",10331 => "10001101",10332 => "00100011",10333 => "01110101",10334 => "00011100",10335 => "01101011",10336 => "10010100",10337 => "10001111",10338 => "01101010",10339 => "00010010",10340 => "10010101",10341 => "10000101",10342 => "00000100",10343 => "01100010",10344 => "11110110",10345 => "11101111",10346 => "00100000",10347 => "11100000",10348 => "10101110",10349 => "10110001",10350 => "11111101",10351 => "11101100",10352 => "00000011",10353 => "01101010",10354 => "11100110",10355 => "10011010",10356 => "00001000",10357 => "11111111",10358 => "10000001",10359 => "10010000",10360 => "00010000",10361 => "00111001",10362 => "10111111",10363 => "11110011",10364 => "10000100",10365 => "11001101",10366 => "10111001",10367 => "10100011",10368 => "00100010",10369 => "10011010",10370 => "01001001",10371 => "11001001",10372 => "01100011",10373 => "00100001",10374 => "11011010",10375 => "01111100",10376 => "11110101",10377 => "00110000",10378 => "01011100",10379 => "11011010",10380 => "10010011",10381 => "11101100",10382 => "00001100",10383 => "00000010",10384 => "11100010",10385 => "00011000",10386 => "10111001",10387 => "00011100",10388 => "00111010",10389 => "01011000",10390 => "00101101",10391 => "01000010",10392 => "00000011",10393 => "01100001",10394 => "10101101",10395 => "10100100",10396 => "00001000",10397 => "01100010",10398 => "01100000",10399 => "10111101",10400 => "01001110",10401 => "11010111",10402 => "11010100",10403 => "11100101",10404 => "00100010",10405 => "01101000",10406 => "11101010",10407 => "01110010",10408 => "10011110",10409 => "00000011",10410 => "10111100",10411 => "01010111",10412 => "11101011",10413 => "00001110",10414 => "00100101",10415 => "11010001",10416 => "11001010",10417 => "00000101",10418 => "10110111",10419 => "01101110",10420 => "10110110",10421 => "11011110",10422 => "01011110",10423 => "00000100",10424 => "11111110",10425 => "11001100",10426 => "01010100",10427 => "10001000",10428 => "01100111",10429 => "10101011",10430 => "10110101",10431 => "01110110",10432 => "01100110",10433 => "11111100",10434 => "10011001",10435 => "11011100",10436 => "10010010",10437 => "01111100",10438 => "11111100",10439 => "11000011",10440 => "01101001",10441 => "01001010",10442 => "01111001",10443 => "01100011",10444 => "01110111",10445 => "11110000",10446 => "11110100",10447 => "01101110",10448 => "01010000",10449 => "10100010",10450 => "11101000",10451 => "00110010",10452 => "11010000",10453 => "11111110",10454 => "01111110",10455 => "00111010",10456 => "11110101",10457 => "10111010",10458 => "00010011",10459 => "11010010",10460 => "11101111",10461 => "01100010",10462 => "11100010",10463 => "00100011",10464 => "00111111",10465 => "00111110",10466 => "00000110",10467 => "00100110",10468 => "01111011",10469 => "10011101",10470 => "00101000",10471 => "10110101",10472 => "11011110",10473 => "11011010",10474 => "00000101",10475 => "10010001",10476 => "11101011",10477 => "11011100",10478 => "00101010",10479 => "00100110",10480 => "10100100",10481 => "00001000",10482 => "11100111",10483 => "10111001",10484 => "00010111",10485 => "10000000",10486 => "00010010",10487 => "01010111",10488 => "01010111",10489 => "10000111",10490 => "10000111",10491 => "11101010",10492 => "10011000",10493 => "10111101",10494 => "00011000",10495 => "11111110",10496 => "10000001",10497 => "01001000",10498 => "10010101",10499 => "00001100",10500 => "00110100",10501 => "10011001",10502 => "10100000",10503 => "11010100",10504 => "10011001",10505 => "10001111",10506 => "00010110",10507 => "10111110",10508 => "10100011",10509 => "00011001",10510 => "11111101",10511 => "01010110",10512 => "11001101",10513 => "11011110",10514 => "10011100",10515 => "10110001",10516 => "11111010",10517 => "10000001",10518 => "10011101",10519 => "10100010",10520 => "00010110",10521 => "11000110",10522 => "00000001",10523 => "11100101",10524 => "11011001",10525 => "10100011",10526 => "00100000",10527 => "01101000",10528 => "11001011",10529 => "10110010",10530 => "01011110",10531 => "01111011",10532 => "10110110",10533 => "10011110",10534 => "00101101",10535 => "11110110",10536 => "11010010",10537 => "00010111",10538 => "11010000",10539 => "00001110",10540 => "11010111",10541 => "10110110",10542 => "10111001",10543 => "00000101",10544 => "00111001",10545 => "11111010",10546 => "00000000",10547 => "10000000",10548 => "10010100",10549 => "11100011",10550 => "11010110",10551 => "11010101",10552 => "01010011",10553 => "01000110",10554 => "00010000",10555 => "00111011",10556 => "00100111",10557 => "11111000",10558 => "10001001",10559 => "10111111",10560 => "11011011",10561 => "00001001",10562 => "11001100",10563 => "01110000",10564 => "10111010",10565 => "01011101",10566 => "01111110",10567 => "10111111",10568 => "00000000",10569 => "11101111",10570 => "01011001",10571 => "00010010",10572 => "00101001",10573 => "00011000",10574 => "01110011",10575 => "10000100",10576 => "10101100",10577 => "00110100",10578 => "10010010",10579 => "00111101",10580 => "00000100",10581 => "01001010",10582 => "01001010",10583 => "10101001",10584 => "11111100",10585 => "10000010",10586 => "11000000",10587 => "01001111",10588 => "11110100",10589 => "01111111",10590 => "11110011",10591 => "11000001",10592 => "01101110",10593 => "11111110",10594 => "11001001",10595 => "01011010",10596 => "00000000",10597 => "10010001",10598 => "01100010",10599 => "01111100",10600 => "01100110",10601 => "10100001",10602 => "11111101",10603 => "00111111",10604 => "01011011",10605 => "11111110",10606 => "11011100",10607 => "00100110",10608 => "11001000",10609 => "10100110",10610 => "00111010",10611 => "11100110",10612 => "01101110",10613 => "11001010",10614 => "10100010",10615 => "11100001",10616 => "11000000",10617 => "01111111",10618 => "01010110",10619 => "01110110",10620 => "01110001",10621 => "00110011",10622 => "10111110",10623 => "10101000",10624 => "00010110",10625 => "01010100",10626 => "10110011",10627 => "11110100",10628 => "00001111",10629 => "01000101",10630 => "00010001",10631 => "00011111",10632 => "10101011",10633 => "00111010",10634 => "00101111",10635 => "10011110",10636 => "10101010",10637 => "11010011",10638 => "01110000",10639 => "01001000",10640 => "10100111",10641 => "00100101",10642 => "00111011",10643 => "00101011",10644 => "11111101",10645 => "11000011",10646 => "11010011",10647 => "01010100",10648 => "01111110",10649 => "00111100",10650 => "10001011",10651 => "01000001",10652 => "00100110",10653 => "10010011",10654 => "10010010",10655 => "11011011",10656 => "00100110",10657 => "11000001",10658 => "11101100",10659 => "11011001",10660 => "00101101",10661 => "01101101",10662 => "11110101",10663 => "10111101",10664 => "00110111",10665 => "01000100",10666 => "00111100",10667 => "10101001",10668 => "00000110",10669 => "10111010",10670 => "00101010",10671 => "11110110",10672 => "00010101",10673 => "10100110",10674 => "11000110",10675 => "11110101",10676 => "00100100",10677 => "11000010",10678 => "01100001",10679 => "01110101",10680 => "00000100",10681 => "11000110",10682 => "01101110",10683 => "10100111",10684 => "10001111",10685 => "01000110",10686 => "11010101",10687 => "11110001",10688 => "01011110",10689 => "11011110",10690 => "00000100",10691 => "00011111",10692 => "10000010",10693 => "00111000",10694 => "10001010",10695 => "11111110",10696 => "11100111",10697 => "01000110",10698 => "01001010",10699 => "01001000",10700 => "01110011",10701 => "00101100",10702 => "10010010",10703 => "00000011",10704 => "01011000",10705 => "10001001",10706 => "10000000",10707 => "01010101",10708 => "10001010",10709 => "01011010",10710 => "10011100",10711 => "11011110",10712 => "11001101",10713 => "11100100",10714 => "10111010",10715 => "10010010",10716 => "11110000",10717 => "11100110",10718 => "11100100",10719 => "01101010",10720 => "11000001",10721 => "10111001",10722 => "01001111",10723 => "01110110",10724 => "01010111",10725 => "01100000",10726 => "00011011",10727 => "10101000",10728 => "10001011",10729 => "10111100",10730 => "10000101",10731 => "11110010",10732 => "00011100",10733 => "00001000",10734 => "11000101",10735 => "11110000",10736 => "10111000",10737 => "10100000",10738 => "00011110",10739 => "11110101",10740 => "10001011",10741 => "01001010",10742 => "10001101",10743 => "10010110",10744 => "11011100",10745 => "10001000",10746 => "11100100",10747 => "11001010",10748 => "00011001",10749 => "11111010",10750 => "11110001",10751 => "00100000",10752 => "11110111",10753 => "00101100",10754 => "01100001",10755 => "00110101",10756 => "10100110",10757 => "10111000",10758 => "01111000",10759 => "00011001",10760 => "11010101",10761 => "01010110",10762 => "10110001",10763 => "10100101",10764 => "10001111",10765 => "11011010",10766 => "10101001",10767 => "01010110",10768 => "00001101",10769 => "10110110",10770 => "10010100",10771 => "11101000",10772 => "00011000",10773 => "11111011",10774 => "11010000",10775 => "10101001",10776 => "01110100",10777 => "00100100",10778 => "01101100",10779 => "00110100",10780 => "01101001",10781 => "00101000",10782 => "01110001",10783 => "11011100",10784 => "11001000",10785 => "00110110",10786 => "00000001",10787 => "11100000",10788 => "10001111",10789 => "10001011",10790 => "00000010",10791 => "01010110",10792 => "10010010",10793 => "10101101",10794 => "01101101",10795 => "01111011",10796 => "00101010",10797 => "01010000",10798 => "11010001",10799 => "00100000",10800 => "11011101",10801 => "00101110",10802 => "01101011",10803 => "00000000",10804 => "11111010",10805 => "10100101",10806 => "00101110",10807 => "10011011",10808 => "11010110",10809 => "10011001",10810 => "01011111",10811 => "10100110",10812 => "11001010",10813 => "00010110",10814 => "00110001",10815 => "10111001",10816 => "10011001",10817 => "01101100",10818 => "01110000",10819 => "11101000",10820 => "00100100",10821 => "01100100",10822 => "11000011",10823 => "01011100",10824 => "11000001",10825 => "01101010",10826 => "11001110",10827 => "01000000",10828 => "10010000",10829 => "00110100",10830 => "00000001",10831 => "11111000",10832 => "10111100",10833 => "10001100",10834 => "01011110",10835 => "11000001",10836 => "00010011",10837 => "11010110",10838 => "01000001",10839 => "11111100",10840 => "11110101",10841 => "01110011",10842 => "01010101",10843 => "10011011",10844 => "11110110",10845 => "10001101",10846 => "01011011",10847 => "01010101",10848 => "10101100",10849 => "01000111",10850 => "01110001",10851 => "11011010",10852 => "01000001",10853 => "11111101",10854 => "11110101",10855 => "10100101",10856 => "00110010",10857 => "10011111",10858 => "11000110",10859 => "00101101",10860 => "00000000",10861 => "11000011",10862 => "11110000",10863 => "10100111",10864 => "01111010",10865 => "10110101",10866 => "11110111",10867 => "00010011",10868 => "10010000",10869 => "10110100",10870 => "10110111",10871 => "01100010",10872 => "10101111",10873 => "00011100",10874 => "01111100",10875 => "01111010",10876 => "11000100",10877 => "00110100",10878 => "10110001",10879 => "10101000",10880 => "01001001",10881 => "10001101",10882 => "10001101",10883 => "01111100",10884 => "01001000",10885 => "10000101",10886 => "10000001",10887 => "00101000",10888 => "10110011",10889 => "11110011",10890 => "00011100",10891 => "11100010",10892 => "00100110",10893 => "01101000",10894 => "11010000",10895 => "10110010",10896 => "01101110",10897 => "01011101",10898 => "10011001",10899 => "00100100",10900 => "01110101",10901 => "00001100",10902 => "10011100",10903 => "01110100",10904 => "11110110",10905 => "10011100",10906 => "11010101",10907 => "10101110",10908 => "01011000",10909 => "11111100",10910 => "10100010",10911 => "11010111",10912 => "10111010",10913 => "01111011",10914 => "01100011",10915 => "10011011",10916 => "11001101",10917 => "01010010",10918 => "00110100",10919 => "00111111",10920 => "01010000",10921 => "01011000",10922 => "11000111",10923 => "10101110",10924 => "11101100",10925 => "00110001",10926 => "11110110",10927 => "00010110",10928 => "00101101",10929 => "01000000",10930 => "00011011",10931 => "00000110",10932 => "11100000",10933 => "01011011",10934 => "11100001",10935 => "11000011",10936 => "11110110",10937 => "11101110",10938 => "01011110",10939 => "11101000",10940 => "01001011",10941 => "00101010",10942 => "00100110",10943 => "11001100",10944 => "10110000",10945 => "01000111",10946 => "00010011",10947 => "01001110",10948 => "10000010",10949 => "11101011",10950 => "01011100",10951 => "11100001",10952 => "00000101",10953 => "01000000",10954 => "11101010",10955 => "10100011",10956 => "11000100",10957 => "11100110",10958 => "11001000",10959 => "01001011",10960 => "00111001",10961 => "10100100",10962 => "00101011",10963 => "00010101",10964 => "00110011",10965 => "00101010",10966 => "11101010",10967 => "01010011",10968 => "11011110",10969 => "00001101",10970 => "10001100",10971 => "00110001",10972 => "10100101",10973 => "00011101",10974 => "00110011",10975 => "11100000",10976 => "10010010",10977 => "11011110",10978 => "00110110",10979 => "10101011",10980 => "10101101",10981 => "01010011",10982 => "11100000",10983 => "01010110",10984 => "00101000",10985 => "10011101",10986 => "10101011",10987 => "01101011",10988 => "10000010",10989 => "11110011",10990 => "11101100",10991 => "11100011",10992 => "11011110",10993 => "01111001",10994 => "00111010",10995 => "10001001",10996 => "01100110",10997 => "01111011",10998 => "11111110",10999 => "01100000",11000 => "00010010",11001 => "00110010",11002 => "10010101",11003 => "01011110",11004 => "00011001",11005 => "00110011",11006 => "11100110",11007 => "11111000",11008 => "00111000",11009 => "01100001",11010 => "00001101",11011 => "11101101",11012 => "10100100",11013 => "01100011",11014 => "10101011",11015 => "00010011",11016 => "00111100",11017 => "00000000",11018 => "11101011",11019 => "10011101",11020 => "10111011",11021 => "11111100",11022 => "01110100",11023 => "01001110",11024 => "10101110",11025 => "10110100",11026 => "11101000",11027 => "01011000",11028 => "10010011",11029 => "00100111",11030 => "10100010",11031 => "11000100",11032 => "11101011",11033 => "00101111",11034 => "01001101",11035 => "01010111",11036 => "00110000",11037 => "10111101",11038 => "10111011",11039 => "01010111",11040 => "00110110",11041 => "10000100",11042 => "11100101",11043 => "00001100",11044 => "11001110",11045 => "11000000",11046 => "10101000",11047 => "11011101",11048 => "11000111",11049 => "01101110",11050 => "10000111",11051 => "01100011",11052 => "11111111",11053 => "10010110",11054 => "10001001",11055 => "10101001",11056 => "01000101",11057 => "11000011",11058 => "01001101",11059 => "00100011",11060 => "00101100",11061 => "11111100",11062 => "01111100",11063 => "11000110",11064 => "00010010",11065 => "10100011",11066 => "00001000",11067 => "10011010",11068 => "11000110",11069 => "11000000",11070 => "11000110",11071 => "01100100",11072 => "10100001",11073 => "01111110",11074 => "01100000",11075 => "11000000",11076 => "00000001",11077 => "10010100",11078 => "10011000",11079 => "01010001",11080 => "00101101",11081 => "00111001",11082 => "00101011",11083 => "01001101",11084 => "00000111",11085 => "00010110",11086 => "01010010",11087 => "01011100",11088 => "10101010",11089 => "00101000",11090 => "11000010",11091 => "10100001",11092 => "11111001",11093 => "01011101",11094 => "10111100",11095 => "01010001",11096 => "00110100",11097 => "11101010",11098 => "01100001",11099 => "10100110",11100 => "01101011",11101 => "10010110",11102 => "11101101",11103 => "10010111",11104 => "10000000",11105 => "10001111",11106 => "10101100",11107 => "00001001",11108 => "10011100",11109 => "01011110",11110 => "01011100",11111 => "00110000",11112 => "00010101",11113 => "10000000",11114 => "11110101",11115 => "01101011",11116 => "11010000",11117 => "11001011",11118 => "11010101",11119 => "01100100",11120 => "10010011",11121 => "01111001",11122 => "10111001",11123 => "11111101",11124 => "11110010",11125 => "11010110",11126 => "11101000",11127 => "11110001",11128 => "00001100",11129 => "01100101",11130 => "10111100",11131 => "11010100",11132 => "10111101",11133 => "11000000",11134 => "11011001",11135 => "11001001",11136 => "10001001",11137 => "11111100",11138 => "00010111",11139 => "01010110",11140 => "10011100",11141 => "10101010",11142 => "11110111",11143 => "01010100",11144 => "01101110",11145 => "01010011",11146 => "01001110",11147 => "10011111",11148 => "11100010",11149 => "10011101",11150 => "11110110",11151 => "10011111",11152 => "10110100",11153 => "11101010",11154 => "00110101",11155 => "00001110",11156 => "01101011",11157 => "11110100",11158 => "01101100",11159 => "01010001",11160 => "01000110",11161 => "11011001",11162 => "10010100",11163 => "10100000",11164 => "01001101",11165 => "10111101",11166 => "11110100",11167 => "00011011",11168 => "10010111",11169 => "10110101",11170 => "00110001",11171 => "00100010",11172 => "10011001",11173 => "01000010",11174 => "01000011",11175 => "11011000",11176 => "11110101",11177 => "10100101",11178 => "00001110",11179 => "10111101",11180 => "00111110",11181 => "11110010",11182 => "00111010",11183 => "11101011",11184 => "01000011",11185 => "00101111",11186 => "01110111",11187 => "00000010",11188 => "01110010",11189 => "01001110",11190 => "10100111",11191 => "00011101",11192 => "01111111",11193 => "11001101",11194 => "00111011",11195 => "00101101",11196 => "11100101",11197 => "10000110",11198 => "01111010",11199 => "00011011",11200 => "11101110",11201 => "11101111",11202 => "11011010",11203 => "01101100",11204 => "10100010",11205 => "10110001",11206 => "01111110",11207 => "10111101",11208 => "11110000",11209 => "11011100",11210 => "00011111",11211 => "11001111",11212 => "00000101",11213 => "01100100",11214 => "10001101",11215 => "10000101",11216 => "10101000",11217 => "10011110",11218 => "01111100",11219 => "10000111",11220 => "10000101",11221 => "01101011",11222 => "11001010",11223 => "10001011",11224 => "01101001",11225 => "11011111",11226 => "00110101",11227 => "11001100",11228 => "10111011",11229 => "11001100",11230 => "11101001",11231 => "11101111",11232 => "10011111",11233 => "01011000",11234 => "10110001",11235 => "10100011",11236 => "11000001",11237 => "10101100",11238 => "00101000",11239 => "10110111",11240 => "11111110",11241 => "00010001",11242 => "01100010",11243 => "11001111",11244 => "11111101",11245 => "01110100",11246 => "11111110",11247 => "00001001",11248 => "11001101",11249 => "00110111",11250 => "10010110",11251 => "00111100",11252 => "11110000",11253 => "00010100",11254 => "00010001",11255 => "00000101",11256 => "11001000",11257 => "01000010",11258 => "11110111",11259 => "11010101",11260 => "11100000",11261 => "00001000",11262 => "01000000",11263 => "10001010",11264 => "00100010",11265 => "01010001",11266 => "10111110",11267 => "01100000",11268 => "00110001",11269 => "11100111",11270 => "00011100",11271 => "10110011",11272 => "10111100",11273 => "11000101",11274 => "10001000",11275 => "10010110",11276 => "00010101",11277 => "01011110",11278 => "01011011",11279 => "01011010",11280 => "01011110",11281 => "00110010",11282 => "10101000",11283 => "00100111",11284 => "01001011",11285 => "01100010",11286 => "00001001",11287 => "11110110",11288 => "00110000",11289 => "00001000",11290 => "11100110",11291 => "01101110",11292 => "01100110",11293 => "01110110",11294 => "10110011",11295 => "00111000",11296 => "00110001",11297 => "11111010",11298 => "10110011",11299 => "01111010",11300 => "01100000",11301 => "11001000",11302 => "10100110",11303 => "00111100",11304 => "10100010",11305 => "10111010",11306 => "11010011",11307 => "11100100",11308 => "00110111",11309 => "01000001",11310 => "10111011",11311 => "00011011",11312 => "10111001",11313 => "00001001",11314 => "10101110",11315 => "11101010",11316 => "11010010",11317 => "11011100",11318 => "11100011",11319 => "00101110",11320 => "01010011",11321 => "01100110",11322 => "00100101",11323 => "01110101",11324 => "11001001",11325 => "10100000",11326 => "01110000",11327 => "00011001",11328 => "11010000",11329 => "01100110",11330 => "10010011",11331 => "10100100",11332 => "01000001",11333 => "10110110",11334 => "00110010",11335 => "01001001",11336 => "11000110",11337 => "01111000",11338 => "10011110",11339 => "11000001",11340 => "01100110",11341 => "01001010",11342 => "00110110",11343 => "10110010",11344 => "01001001",11345 => "10101011",11346 => "00001000",11347 => "01000000",11348 => "00001000",11349 => "11100010",11350 => "00110011",11351 => "11100010",11352 => "01111001",11353 => "10101101",11354 => "11010011",11355 => "00000000",11356 => "10011100",11357 => "00110110",11358 => "01100111",11359 => "11110111",11360 => "00110011",11361 => "10010010",11362 => "10010000",11363 => "00011010",11364 => "11100110",11365 => "11001000",11366 => "00001111",11367 => "11111001",11368 => "11010111",11369 => "01111010",11370 => "11111011",11371 => "01000001",11372 => "11111011",11373 => "01110010",11374 => "11101101",11375 => "11000010",11376 => "00101011",11377 => "01101000",11378 => "00111101",11379 => "10111010",11380 => "11011111",11381 => "10100011",11382 => "11001100",11383 => "01110100",11384 => "11010100",11385 => "00011010",11386 => "01101101",11387 => "11110001",11388 => "10010100",11389 => "11111001",11390 => "00110010",11391 => "01101101",11392 => "00110101",11393 => "11110001",11394 => "00111001",11395 => "01010011",11396 => "11101001",11397 => "11000001",11398 => "11011010",11399 => "11101101",11400 => "00011110",11401 => "01110001",11402 => "11111010",11403 => "11010111",11404 => "00101010",11405 => "10111010",11406 => "10001100",11407 => "11101011",11408 => "00001001",11409 => "11010011",11410 => "10000010",11411 => "11010000",11412 => "00010000",11413 => "11101100",11414 => "00100000",11415 => "01011011",11416 => "00111100",11417 => "11000001",11418 => "00110000",11419 => "00001110",11420 => "01001101",11421 => "10011001",11422 => "01011001",11423 => "00111001",11424 => "01100011",11425 => "00000101",11426 => "11000011",11427 => "10000111",11428 => "11111011",11429 => "10100000",11430 => "10110011",11431 => "10101111",11432 => "11110110",11433 => "10011001",11434 => "00110001",11435 => "10011011",11436 => "00100010",11437 => "01111111",11438 => "10010100",11439 => "10011101",11440 => "01100010",11441 => "11110110",11442 => "10110011",11443 => "10011010",11444 => "11001000",11445 => "11100101",11446 => "01101000",11447 => "00110010",11448 => "10100011",11449 => "11000101",11450 => "00001110",11451 => "01111111",11452 => "00001000",11453 => "11100100",11454 => "01100000",11455 => "11111000",11456 => "01010101",11457 => "10101001",11458 => "00011100",11459 => "11000111",11460 => "10111110",11461 => "01100101",11462 => "01000111",11463 => "00011110",11464 => "00111110",11465 => "01000010",11466 => "00110100",11467 => "11110010",11468 => "10011110",11469 => "10001100",11470 => "11101101",11471 => "10000001",11472 => "01011111",11473 => "10101001",11474 => "01011010",11475 => "11010101",11476 => "11111000",11477 => "01101000",11478 => "01001110",11479 => "01111100",11480 => "11011111",11481 => "00000011",11482 => "11010101",11483 => "00000110",11484 => "01111010",11485 => "10010011",11486 => "01010010",11487 => "01011011",11488 => "11100011",11489 => "10100011",11490 => "10001110",11491 => "11001100",11492 => "00101011",11493 => "01100111",11494 => "10100101",11495 => "01011001",11496 => "01100100",11497 => "10101101",11498 => "10001110",11499 => "01000011",11500 => "00101010",11501 => "00100010",11502 => "01011110",11503 => "11010100",11504 => "11000100",11505 => "01110110",11506 => "00010001",11507 => "11011110",11508 => "00000011",11509 => "01000101",11510 => "01101101",11511 => "00101110",11512 => "11111101",11513 => "10110100",11514 => "11101011",11515 => "10110001",11516 => "01101001",11517 => "00101100",11518 => "11111001",11519 => "00111000",11520 => "11101011",11521 => "00010000",11522 => "00010001",11523 => "10011100",11524 => "11111111",11525 => "01110110",11526 => "11110100",11527 => "10111100",11528 => "01110110",11529 => "11010000",11530 => "10111111",11531 => "00001000",11532 => "11110000",11533 => "01010010",11534 => "00111101",11535 => "01010011",11536 => "00111000",11537 => "00010110",11538 => "00001100",11539 => "10101010",11540 => "00100000",11541 => "01011110",11542 => "01101000",11543 => "00111111",11544 => "01100110",11545 => "01000100",11546 => "11011110",11547 => "10001111",11548 => "00000011",11549 => "00100101",11550 => "11001011",11551 => "00011110",11552 => "01111101",11553 => "11001000",11554 => "10001101",11555 => "00100101",11556 => "00001101",11557 => "01101001",11558 => "11010100",11559 => "01000010",11560 => "10100011",11561 => "11101001",11562 => "10010111",11563 => "11111111",11564 => "01000001",11565 => "01001010",11566 => "10000101",11567 => "10001011",11568 => "11110000",11569 => "01001110",11570 => "01110000",11571 => "10001101",11572 => "10110100",11573 => "01001001",11574 => "01100011",11575 => "11001100",11576 => "01110001",11577 => "11100011",11578 => "11001100",11579 => "01101000",11580 => "10010100",11581 => "11101011",11582 => "01011100",11583 => "00110011",11584 => "10100011",11585 => "00001110",11586 => "00001011",11587 => "01001110",11588 => "00001000",11589 => "01011000",11590 => "00100101",11591 => "01010101",11592 => "00110001",11593 => "11101111",11594 => "10001110",11595 => "01010111",11596 => "10001101",11597 => "01100000",11598 => "00110001",11599 => "01010010",11600 => "11101100",11601 => "10101010",11602 => "00001011",11603 => "01000111",11604 => "00001010",11605 => "11101110",11606 => "00011111",11607 => "00110110",11608 => "00011100",11609 => "01110111",11610 => "10110111",11611 => "01001110",11612 => "10110000",11613 => "10001000",11614 => "00001010",11615 => "01001010",11616 => "11111101",11617 => "11000000",11618 => "11101111",11619 => "01001111",11620 => "00100010",11621 => "01110001",11622 => "01010001",11623 => "00111111",11624 => "01010011",11625 => "00111101",11626 => "00110101",11627 => "11001010",11628 => "00110110",11629 => "00010101",11630 => "00100011",11631 => "01110011",11632 => "11000010",11633 => "10010100",11634 => "10110110",11635 => "10100010",11636 => "00010010",11637 => "11010011",11638 => "01000001",11639 => "01000101",11640 => "10100110",11641 => "10011011",11642 => "00000101",11643 => "10111110",11644 => "10001010",11645 => "01111100",11646 => "10100110",11647 => "11110111",11648 => "11010111",11649 => "11110101",11650 => "00101011",11651 => "11001100",11652 => "00010101",11653 => "00000111",11654 => "11101101",11655 => "10011001",11656 => "11001000",11657 => "00100001",11658 => "01000100",11659 => "01010110",11660 => "01001001",11661 => "00001001",11662 => "10001011",11663 => "00000111",11664 => "00000001",11665 => "00100110",11666 => "00001000",11667 => "01000110",11668 => "01111001",11669 => "10000011",11670 => "10110001",11671 => "10010011",11672 => "00101011",11673 => "11010010",11674 => "01111111",11675 => "11000101",11676 => "00001000",11677 => "01111001",11678 => "00100110",11679 => "11001011",11680 => "00001001",11681 => "01100000",11682 => "01100100",11683 => "11000101",11684 => "00110011",11685 => "10011100",11686 => "11000000",11687 => "11101001",11688 => "11100110",11689 => "10001010",11690 => "01000011",11691 => "11101111",11692 => "10001110",11693 => "01110100",11694 => "10111001",11695 => "10111001",11696 => "11100001",11697 => "00110010",11698 => "11100010",11699 => "10010111",11700 => "11110000",11701 => "01011001",11702 => "11110000",11703 => "10010100",11704 => "10011010",11705 => "01011000",11706 => "00000111",11707 => "01010111",11708 => "01110101",11709 => "10001110",11710 => "10001011",11711 => "11001101",11712 => "00110100",11713 => "01111110",11714 => "01111010",11715 => "01101010",11716 => "01100111",11717 => "00001100",11718 => "01001001",11719 => "10011100",11720 => "11001100",11721 => "10111100",11722 => "00000100",11723 => "00010010",11724 => "11011101",11725 => "00111000",11726 => "11010110",11727 => "00111011",11728 => "10111010",11729 => "01100101",11730 => "11100100",11731 => "10111101",11732 => "01010001",11733 => "00100100",11734 => "00001111",11735 => "11000011",11736 => "00000111",11737 => "10011111",11738 => "10101011",11739 => "11001101",11740 => "11100011",11741 => "01011100",11742 => "10110011",11743 => "10000111",11744 => "00100110",11745 => "11101010",11746 => "10111010",11747 => "11111011",11748 => "10001000",11749 => "01100111",11750 => "10100101",11751 => "00101001",11752 => "00010001",11753 => "10101010",11754 => "01011010",11755 => "00010111",11756 => "11000010",11757 => "00100001",11758 => "00110010",11759 => "01100110",11760 => "00111001",11761 => "11010110",11762 => "10010110",11763 => "11000010",11764 => "00001011",11765 => "10010001",11766 => "11011001",11767 => "00100010",11768 => "11110101",11769 => "10100000",11770 => "11001001",11771 => "11000100",11772 => "00101000",11773 => "01101110",11774 => "10010001",11775 => "00011000",11776 => "11101000",11777 => "00011101",11778 => "01011100",11779 => "11001111",11780 => "00010111",11781 => "10011011",11782 => "11100000",11783 => "11111111",11784 => "10001000",11785 => "00100111",11786 => "01101000",11787 => "00001001",11788 => "10011001",11789 => "11000111",11790 => "11111110",11791 => "11111010",11792 => "00001101",11793 => "11101111",11794 => "10110110",11795 => "10001011",11796 => "00000011",11797 => "00110111",11798 => "00110100",11799 => "10000110",11800 => "00111110",11801 => "11011100",11802 => "11010100",11803 => "00100100",11804 => "11101011",11805 => "01100100",11806 => "11101001",11807 => "00000010",11808 => "10110110",11809 => "01100101",11810 => "00001100",11811 => "11100011",11812 => "11011000",11813 => "11011110",11814 => "01100110",11815 => "10000101",11816 => "11000100",11817 => "00010000",11818 => "01011101",11819 => "00111111",11820 => "00110111",11821 => "01001001",11822 => "10000010",11823 => "11011011",11824 => "11000101",11825 => "00110010",11826 => "11011111",11827 => "11101101",11828 => "00010100",11829 => "10001011",11830 => "11000111",11831 => "00100000",11832 => "00011100",11833 => "11000011",11834 => "10110110",11835 => "11011001",11836 => "00001010",11837 => "11101010",11838 => "01011101",11839 => "00010100",11840 => "11001001",11841 => "10010100",11842 => "10100110",11843 => "01101011",11844 => "01010001",11845 => "01010111",11846 => "11111001",11847 => "10010100",11848 => "11011010",11849 => "00100101",11850 => "10010010",11851 => "11110001",11852 => "01110001",11853 => "10111111",11854 => "10001100",11855 => "01001011",11856 => "10001110",11857 => "11000011",11858 => "00110100",11859 => "00001110",11860 => "11011001",11861 => "00110011",11862 => "01000100",11863 => "01110111",11864 => "10001011",11865 => "10100010",11866 => "00110101",11867 => "01001100",11868 => "00000001",11869 => "11100001",11870 => "10111010",11871 => "00100110",11872 => "00101100",11873 => "01111011",11874 => "10111101",11875 => "00111011",11876 => "10010001",11877 => "11101100",11878 => "11100110",11879 => "11010010",11880 => "00000111",11881 => "00111001",11882 => "01001000",11883 => "00101011",11884 => "01000101",11885 => "11011101",11886 => "11111011",11887 => "10000011",11888 => "01101011",11889 => "01110111",11890 => "10111110",11891 => "10010100",11892 => "01101001",11893 => "11000111",11894 => "00001110",11895 => "11000101",11896 => "01011101",11897 => "10100100",11898 => "00100101",11899 => "10111000",11900 => "01100101",11901 => "11010000",11902 => "01110010",11903 => "10111011",11904 => "11011010",11905 => "10111000",11906 => "01101101",11907 => "01011010",11908 => "11011100",11909 => "10011011",11910 => "11001001",11911 => "11100001",11912 => "10000111",11913 => "10011010",11914 => "11011101",11915 => "10110010",11916 => "10101100",11917 => "01110111",11918 => "00100101",11919 => "11010111",11920 => "00000110",11921 => "01110000",11922 => "00100000",11923 => "01111110",11924 => "10101100",11925 => "00001001",11926 => "10010011",11927 => "01010001",11928 => "00111100",11929 => "10000010",11930 => "11111100",11931 => "11100111",11932 => "01101111",11933 => "11101100",11934 => "10101000",11935 => "11010110",11936 => "00110010",11937 => "10100001",11938 => "11000000",11939 => "10011110",11940 => "11100111",11941 => "01001000",11942 => "10101011",11943 => "11000011",11944 => "01101010",11945 => "11010110",11946 => "00101111",11947 => "01000011",11948 => "10110001",11949 => "01110010",11950 => "00000010",11951 => "01111000",11952 => "11101110",11953 => "01101111",11954 => "11000000",11955 => "11110100",11956 => "01100101",11957 => "01111111",11958 => "10101100",11959 => "01000111",11960 => "10101000",11961 => "01011001",11962 => "00110111",11963 => "11101010",11964 => "00010010",11965 => "11110111",11966 => "10000101",11967 => "10100100",11968 => "01010101",11969 => "00010010",11970 => "00100111",11971 => "01111011",11972 => "01100100",11973 => "10011000",11974 => "00000000",11975 => "01001011",11976 => "00001010",11977 => "01000110",11978 => "11101000",11979 => "01001010",11980 => "10010111",11981 => "11011101",11982 => "11111100",11983 => "10001000",11984 => "11111101",11985 => "00001001",11986 => "11000011",11987 => "10011011",11988 => "01111100",11989 => "10100110",11990 => "00010100",11991 => "10001011",11992 => "00100101",11993 => "01100010",11994 => "00101101",11995 => "10100000",11996 => "10100100",11997 => "11001001",11998 => "10010101",11999 => "11110110",12000 => "11111010",12001 => "10000101",12002 => "01111000",12003 => "10000100",12004 => "11011110",12005 => "00001101",12006 => "10000110",12007 => "01111000",12008 => "10001101",12009 => "01111000",12010 => "10111100",12011 => "10100011",12012 => "11100001",12013 => "10111100",12014 => "11111111",12015 => "01100011",12016 => "10010000",12017 => "01100010",12018 => "00011011",12019 => "10111100",12020 => "11110110",12021 => "00111101",12022 => "01011100",12023 => "00011111",12024 => "00101110",12025 => "01101110",12026 => "11001011",12027 => "10011111",12028 => "01110101",12029 => "01000000",12030 => "00010111",12031 => "11111000",12032 => "11001011",12033 => "11110000",12034 => "11110001",12035 => "00111010",12036 => "11000010",12037 => "10011110",12038 => "10001100",12039 => "10101011",12040 => "10001110",12041 => "11111010",12042 => "11000111",12043 => "00100011",12044 => "01000010",12045 => "11101000",12046 => "10101011",12047 => "11101010",12048 => "10001000",12049 => "10000111",12050 => "11101011",12051 => "01101100",12052 => "01000011",12053 => "00100101",12054 => "00001011",12055 => "10011100",12056 => "00011101",12057 => "11010001",12058 => "11001010",12059 => "00111100",12060 => "01001111",12061 => "10010111",12062 => "10111100",12063 => "00101011",12064 => "01101101",12065 => "10010100",12066 => "11110101",12067 => "01111111",12068 => "01011000",12069 => "10010111",12070 => "01000011",12071 => "00111101",12072 => "11001110",12073 => "00110001",12074 => "00111000",12075 => "11101110",12076 => "10100010",12077 => "00010100",12078 => "10100010",12079 => "00001010",12080 => "01100001",12081 => "11101000",12082 => "00011110",12083 => "10000001",12084 => "10011000",12085 => "01000111",12086 => "01010011",12087 => "11101110",12088 => "10000011",12089 => "10011010",12090 => "11000101",12091 => "10101000",12092 => "10111011",12093 => "01000011",12094 => "10110100",12095 => "00001010",12096 => "10011011",12097 => "01000100",12098 => "11000100",12099 => "00100100",12100 => "01000011",12101 => "00000100",12102 => "00100110",12103 => "00010001",12104 => "00111111",12105 => "10111001",12106 => "10001111",12107 => "10000101",12108 => "01001000",12109 => "00001010",12110 => "01011101",12111 => "10100100",12112 => "01011001",12113 => "00110101",12114 => "01011011",12115 => "00110100",12116 => "10010110",12117 => "01111001",12118 => "00011101",12119 => "11000000",12120 => "01100001",12121 => "11001011",12122 => "00111110",12123 => "10100101",12124 => "01000000",12125 => "01110011",12126 => "01111101",12127 => "00100001",12128 => "11001000",12129 => "00110111",12130 => "11100101",12131 => "11000110",12132 => "11000101",12133 => "11101101",12134 => "01000101",12135 => "10100001",12136 => "10110011",12137 => "10101000",12138 => "01000001",12139 => "01000000",12140 => "11001111",12141 => "11001110",12142 => "10101011",12143 => "10110001",12144 => "11110011",12145 => "11001111",12146 => "01000110",12147 => "01110101",12148 => "01111100",12149 => "00011001",12150 => "11100001",12151 => "11000001",12152 => "10100011",12153 => "00010001",12154 => "01001101",12155 => "00111001",12156 => "11111011",12157 => "00110000",12158 => "10110011",12159 => "10101010",12160 => "00101010",12161 => "00111001",12162 => "10110000",12163 => "01101001",12164 => "00000111",12165 => "00110010",12166 => "11011011",12167 => "00011101",12168 => "10001000",12169 => "00111011",12170 => "01111001",12171 => "00100101",12172 => "00110101",12173 => "00010100",12174 => "00101010",12175 => "10100110",12176 => "00100000",12177 => "01101101",12178 => "11000011",12179 => "01100011",12180 => "11011000",12181 => "11100101",12182 => "00001011",12183 => "00111110",12184 => "01110101",12185 => "11010011",12186 => "10111101",12187 => "00011011",12188 => "10100001",12189 => "10110010",12190 => "00110111",12191 => "11101101",12192 => "00101011",12193 => "11111011",12194 => "01111001",12195 => "01110000",12196 => "10100110",12197 => "00011100",12198 => "01100101",12199 => "11000101",12200 => "01100111",12201 => "10100000",12202 => "10001100",12203 => "11111110",12204 => "11001110",12205 => "00010010",12206 => "00100011",12207 => "01101110",12208 => "11010101",12209 => "01011010",12210 => "00110111",12211 => "10000101",12212 => "01001110",12213 => "01101001",12214 => "11100011",12215 => "00101101",12216 => "00011011",12217 => "01000110",12218 => "00001100",12219 => "00001011",12220 => "01110110",12221 => "11101101",12222 => "11110111",12223 => "00000000",12224 => "00110111",12225 => "11000011",12226 => "11011000",12227 => "00001111",12228 => "10000111",12229 => "01101010",12230 => "11010111",12231 => "11010110",12232 => "11101110",12233 => "11110110",12234 => "10000011",12235 => "01011011",12236 => "10101101",12237 => "01110111",12238 => "11111001",12239 => "11110111",12240 => "01111011",12241 => "01100000",12242 => "11001111",12243 => "10101101",12244 => "01111111",12245 => "01000010",12246 => "00100111",12247 => "01000110",12248 => "11010010",12249 => "11100010",12250 => "01010001",12251 => "10111100",12252 => "10101100",12253 => "11100011",12254 => "10000001",12255 => "10011100",12256 => "11111101",12257 => "00101100",12258 => "10110011",12259 => "11101000",12260 => "11001010",12261 => "00010000",12262 => "11111100",12263 => "10011100",12264 => "10010101",12265 => "00111010",12266 => "00010001",12267 => "11101110",12268 => "01011110",12269 => "00111101",12270 => "11010100",12271 => "01011001",12272 => "11001111",12273 => "01010101",12274 => "10011000",12275 => "00011110",12276 => "10110010",12277 => "00001001",12278 => "00110001",12279 => "01101000",12280 => "00010101",12281 => "10011001",12282 => "00011000",12283 => "00110100",12284 => "10011110",12285 => "10001100",12286 => "00111111",12287 => "01100110",12288 => "11000000",12289 => "00001000",12290 => "00000110",12291 => "11010010",12292 => "00011100",12293 => "00000001",12294 => "01011011",12295 => "01011011",12296 => "00000101",12297 => "10111010",12298 => "10011000",12299 => "10001101",12300 => "11011100",12301 => "11001101",12302 => "01001011",12303 => "11001000",12304 => "00001101",12305 => "10010001",12306 => "11011100",12307 => "10111000",12308 => "11110111",12309 => "00011011",12310 => "01100111",12311 => "10011010",12312 => "10011010",12313 => "01000100",12314 => "01010111",12315 => "11001000",12316 => "00000000",12317 => "01101111",12318 => "11100011",12319 => "11100111",12320 => "01000101",12321 => "11001011",12322 => "00000100",12323 => "00000101",12324 => "11101100",12325 => "00000011",12326 => "00011011",12327 => "00111001",12328 => "00110101",12329 => "10100000",12330 => "10101011",12331 => "10000000",12332 => "11111000",12333 => "01100110",12334 => "01000101",12335 => "11010000",12336 => "10101001",12337 => "11010110",12338 => "10001010",12339 => "01010011",12340 => "00110001",12341 => "11000000",12342 => "01000101",12343 => "11101110",12344 => "00011010",12345 => "01110100",12346 => "01111110",12347 => "11101010",12348 => "01011110",12349 => "10011100",12350 => "10010111",12351 => "00010100",12352 => "10000011",12353 => "11100101",12354 => "01110000",12355 => "10101010",12356 => "01010001",12357 => "00101000",12358 => "00001011",12359 => "10010111",12360 => "01101000",12361 => "11011001",12362 => "01001110",12363 => "10111010",12364 => "01011000",12365 => "11111110",12366 => "10011011",12367 => "10001001",12368 => "11011011",12369 => "11100001",12370 => "01111000",12371 => "11011000",12372 => "11110110",12373 => "00101001",12374 => "11110000",12375 => "10110101",12376 => "00101110",12377 => "01000111",12378 => "01101010",12379 => "00011100",12380 => "00011111",12381 => "11001000",12382 => "01110001",12383 => "11111011",12384 => "01001100",12385 => "11111101",12386 => "00110001",12387 => "01000000",12388 => "11101111",12389 => "01101110",12390 => "11010010",12391 => "01000101",12392 => "11001011",12393 => "01110101",12394 => "10011011",12395 => "00100111",12396 => "01001110",12397 => "11010100",12398 => "11101100",12399 => "00100100",12400 => "10010110",12401 => "00000101",12402 => "00111001",12403 => "01010001",12404 => "11010101",12405 => "00111010",12406 => "10000001",12407 => "01010101",12408 => "11111110",12409 => "10010001",12410 => "10100000",12411 => "01101000",12412 => "11101001",12413 => "01001101",12414 => "01001101",12415 => "10001101",12416 => "10110100",12417 => "01000111",12418 => "11010111",12419 => "01111001",12420 => "11000010",12421 => "01110101",12422 => "00100001",12423 => "11100010",12424 => "10011110",12425 => "10000000",12426 => "00000011",12427 => "00110011",12428 => "00000101",12429 => "10110000",12430 => "10001110",12431 => "01110001",12432 => "11111111",12433 => "00010001",12434 => "00111010",12435 => "01100011",12436 => "10001001",12437 => "11000011",12438 => "10000011",12439 => "11000110",12440 => "10110100",12441 => "00011001",12442 => "11101000",12443 => "10000011",12444 => "10100110",12445 => "00010001",12446 => "10111101",12447 => "01111111",12448 => "01100111",12449 => "11111101",12450 => "01100000",12451 => "00101101",12452 => "00011110",12453 => "01100011",12454 => "00110100",12455 => "01111010",12456 => "00011101",12457 => "01100110",12458 => "10100111",12459 => "11011011",12460 => "11011110",12461 => "10010000",12462 => "10111101",12463 => "11101100",12464 => "11010001",12465 => "01100011",12466 => "11111000",12467 => "01110001",12468 => "01111100",12469 => "11010000",12470 => "10001011",12471 => "10001101",12472 => "01000111",12473 => "11110011",12474 => "00101101",12475 => "01101011",12476 => "01110110",12477 => "00110011",12478 => "10100111",12479 => "10001001",12480 => "10001010",12481 => "10010011",12482 => "10011000",12483 => "00000011",12484 => "01010100",12485 => "01101011",12486 => "10110111",12487 => "01100001",12488 => "11100111",12489 => "00111101",12490 => "01000111",12491 => "10001101",12492 => "11010101",12493 => "10010011",12494 => "11111001",12495 => "01001110",12496 => "01010110",12497 => "00000110",12498 => "11010110",12499 => "00111011",12500 => "00110100",12501 => "11100100",12502 => "11001011",12503 => "10000010",12504 => "01111111",12505 => "10011011",12506 => "01010001",12507 => "01111111",12508 => "00011011",12509 => "11010011",12510 => "01011100",12511 => "11011111",12512 => "00000100",12513 => "11000110",12514 => "10110000",12515 => "01100011",12516 => "01101010",12517 => "01111000",12518 => "10101010",12519 => "11000110",12520 => "11110100",12521 => "01111000",12522 => "10010000",12523 => "00111010",12524 => "01011000",12525 => "00000100",12526 => "00001011",12527 => "01101110",12528 => "00001001",12529 => "10000011",12530 => "11001010",12531 => "00001000",12532 => "10001100",12533 => "01111100",12534 => "00111001",12535 => "01110101",12536 => "00010011",12537 => "11001100",12538 => "10110101",12539 => "01011101",12540 => "00001001",12541 => "00001110",12542 => "10001111",12543 => "00111110",12544 => "10111110",12545 => "11101001",12546 => "10110100",12547 => "10000100",12548 => "00011100",12549 => "01111110",12550 => "11001010",12551 => "11110101",12552 => "01001110",12553 => "10100000",12554 => "11011000",12555 => "10010000",12556 => "10101010",12557 => "10010000",12558 => "00101001",12559 => "01111100",12560 => "00100001",12561 => "01010100",12562 => "10110001",12563 => "11011100",12564 => "01000111",12565 => "11110001",12566 => "01110011",12567 => "11000010",12568 => "11111010",12569 => "00001110",12570 => "00110001",12571 => "11000011",12572 => "11100010",12573 => "01001111",12574 => "00101101",12575 => "01101001",12576 => "00100010",12577 => "11100000",12578 => "01000001",12579 => "10111001",12580 => "00001110",12581 => "10001001",12582 => "10101010",12583 => "10001011",12584 => "00111011",12585 => "11101011",12586 => "01101000",12587 => "00111100",12588 => "10110110",12589 => "00111110",12590 => "11000110",12591 => "01101001",12592 => "11100101",12593 => "01000110",12594 => "11110111",12595 => "10110000",12596 => "00100100",12597 => "01111010",12598 => "00000110",12599 => "00110000",12600 => "11011110",12601 => "00000011",12602 => "11001001",12603 => "00001110",12604 => "10000101",12605 => "10011000",12606 => "11001011",12607 => "00010100",12608 => "01001100",12609 => "00111000",12610 => "11000010",12611 => "01011011",12612 => "11101010",12613 => "00110101",12614 => "00111001",12615 => "10000111",12616 => "01110010",12617 => "10111010",12618 => "10011011",12619 => "01000010",12620 => "10110111",12621 => "11100111",12622 => "10101011",12623 => "00101101",12624 => "00000111",12625 => "11110001",12626 => "10101111",12627 => "11000011",12628 => "01000110",12629 => "11000100",12630 => "11110111",12631 => "11011001",12632 => "10111100",12633 => "11010111",12634 => "01111100",12635 => "01011100",12636 => "01010011",12637 => "11011000",12638 => "00110100",12639 => "01010101",12640 => "01001101",12641 => "11111111",12642 => "11101111",12643 => "10100011",12644 => "00011111",12645 => "00100110",12646 => "11110001",12647 => "11100100",12648 => "01111011",12649 => "11111111",12650 => "10001111",12651 => "10110010",12652 => "01111100",12653 => "10001101",12654 => "10011001",12655 => "00101100",12656 => "10110100",12657 => "01110011",12658 => "00001110",12659 => "11101100",12660 => "01110100",12661 => "01010011",12662 => "01100110",12663 => "10010001",12664 => "00110011",12665 => "00100111",12666 => "10001111",12667 => "11000010",12668 => "11110011",12669 => "00001101",12670 => "11101100",12671 => "11001000",12672 => "10011101",12673 => "10100111",12674 => "01110001",12675 => "11011101",12676 => "00010110",12677 => "11011100",12678 => "11000001",12679 => "11110111",12680 => "01100111",12681 => "11110010",12682 => "11111101",12683 => "01001100",12684 => "00011000",12685 => "01000100",12686 => "11001100",12687 => "10000100",12688 => "11010100",12689 => "10000001",12690 => "00000001",12691 => "01011101",12692 => "00100101",12693 => "01110001",12694 => "01101100",12695 => "11010011",12696 => "01001001",12697 => "11111101",12698 => "10100000",12699 => "11011001",12700 => "00111100",12701 => "10110110",12702 => "10011011",12703 => "01111010",12704 => "10001010",12705 => "11010101",12706 => "11110110",12707 => "10010000",12708 => "10011100",12709 => "01101101",12710 => "11001000",12711 => "11110100",12712 => "00000010",12713 => "01101001",12714 => "11000000",12715 => "00000100",12716 => "01111011",12717 => "11100110",12718 => "10011000",12719 => "01001011",12720 => "00010110",12721 => "10011001",12722 => "11011000",12723 => "10100100",12724 => "01101000",12725 => "10101000",12726 => "01101000",12727 => "10010010",12728 => "10001001",12729 => "00110000",12730 => "01011011",12731 => "10110101",12732 => "00000000",12733 => "10111001",12734 => "10111100",12735 => "11001001",12736 => "11100101",12737 => "00010100",12738 => "00010110",12739 => "10000011",12740 => "00100110",12741 => "10101011",12742 => "11011110",12743 => "01011000",12744 => "00111010",12745 => "00110000",12746 => "10010111",12747 => "11010001",12748 => "01111111",12749 => "10101100",12750 => "10010011",12751 => "00111011",12752 => "10111110",12753 => "10111011",12754 => "01001110",12755 => "10001001",12756 => "00101011",12757 => "11101100",12758 => "01000100",12759 => "01011000",12760 => "01010101",12761 => "11110011",12762 => "10000110",12763 => "00110100",12764 => "11001111",12765 => "00000011",12766 => "10111110",12767 => "01011111",12768 => "11100100",12769 => "01100010",12770 => "10011010",12771 => "00001111",12772 => "10001000",12773 => "00110010",12774 => "11111100",12775 => "01011010",12776 => "00101011",12777 => "11010011",12778 => "01101011",12779 => "11111001",12780 => "00110010",12781 => "01000010",12782 => "10110111",12783 => "11011001",12784 => "01101001",12785 => "10101001",12786 => "00101000",12787 => "10101111",12788 => "00111110",12789 => "10110001",12790 => "01100010",12791 => "10000100",12792 => "01100100",12793 => "10101110",12794 => "01001001",12795 => "11011101",12796 => "00000010",12797 => "01001100",12798 => "10100110",12799 => "00100001",12800 => "11100010",12801 => "01100011",12802 => "10111001",12803 => "01100011",12804 => "01011101",12805 => "10010010",12806 => "00110110",12807 => "00000101",12808 => "01000011",12809 => "11010011",12810 => "11101101",12811 => "11011101",12812 => "01001010",12813 => "10010001",12814 => "10111100",12815 => "01011100",12816 => "00100011",12817 => "01000100",12818 => "01101101",12819 => "01001000",12820 => "00000011",12821 => "10100011",12822 => "00110100",12823 => "10011110",12824 => "00010101",12825 => "01001101",12826 => "01001010",12827 => "00001001",12828 => "01110010",12829 => "10011110",12830 => "11001100",12831 => "10011000",12832 => "10110111",12833 => "11000101",12834 => "01011000",12835 => "00011011",12836 => "01000110",12837 => "01010100",12838 => "00101100",12839 => "01000000",12840 => "10001010",12841 => "10011110",12842 => "11000010",12843 => "11001000",12844 => "10101010",12845 => "01011010",12846 => "00101100",12847 => "11000011",12848 => "10110110",12849 => "00001010",12850 => "10010000",12851 => "01011000",12852 => "10100000",12853 => "01011000",12854 => "10011011",12855 => "11011010",12856 => "01011101",12857 => "11101011",12858 => "11101100",12859 => "00111011",12860 => "11111000",12861 => "01110011",12862 => "01101100",12863 => "01001011",12864 => "11101110",12865 => "01000110",12866 => "11111011",12867 => "00001100",12868 => "10001100",12869 => "01000101",12870 => "00001111",12871 => "11111111",12872 => "10000001",12873 => "00101111",12874 => "10100100",12875 => "01000000",12876 => "11101110",12877 => "01111101",12878 => "01110101",12879 => "00111010",12880 => "11111011",12881 => "01000101",12882 => "00100011",12883 => "10010011",12884 => "01001110",12885 => "11110100",12886 => "10101010",12887 => "01010111",12888 => "10101000",12889 => "11001000",12890 => "10010010",12891 => "10001001",12892 => "01100111",12893 => "10011111",12894 => "11000101",12895 => "00111001",12896 => "10000100",12897 => "01111100",12898 => "00001101",12899 => "01101111",12900 => "01000110",12901 => "10001100",12902 => "10011010",12903 => "00111011",12904 => "01011001",12905 => "11111000",12906 => "01111101",12907 => "00101101",12908 => "10111100",12909 => "00000110",12910 => "01011000",12911 => "00100110",12912 => "00100100",12913 => "00110110",12914 => "00011001",12915 => "10000110",12916 => "10100001",12917 => "01011111",12918 => "00110110",12919 => "10110001",12920 => "11010111",12921 => "10011011",12922 => "10000000",12923 => "10011000",12924 => "10101110",12925 => "00010101",12926 => "00001101",12927 => "00001011",12928 => "00111100",12929 => "11101011",12930 => "01100100",12931 => "01111011",12932 => "01011110",12933 => "01010011",12934 => "00000010",12935 => "10000111",12936 => "01001110",12937 => "01010100",12938 => "10010101",12939 => "00010011",12940 => "11001111",12941 => "11101010",12942 => "10000011",12943 => "00011111",12944 => "11101000",12945 => "01110100",12946 => "01110001",12947 => "01000100",12948 => "00100000",12949 => "10101111",12950 => "01100101",12951 => "11000110",12952 => "01100011",12953 => "11111000",12954 => "11000111",12955 => "11111101",12956 => "10000100",12957 => "10010111",12958 => "10110101",12959 => "11101000",12960 => "11000111",12961 => "00001101",12962 => "11010111",12963 => "11101001",12964 => "00100010",12965 => "10011000",12966 => "10110001",12967 => "10010001",12968 => "00110101",12969 => "11010110",12970 => "01100110",12971 => "01011111",12972 => "01111011",12973 => "01101100",12974 => "01001110",12975 => "11010001",12976 => "00111001",12977 => "10101111",12978 => "01101110",12979 => "00110011",12980 => "10100010",12981 => "10000111",12982 => "11111110",12983 => "10111101",12984 => "00001010",12985 => "01001000",12986 => "00001110",12987 => "01111001",12988 => "00110011",12989 => "10011100",12990 => "00101110",12991 => "01011001",12992 => "11110010",12993 => "01011110",12994 => "11110010",12995 => "00111011",12996 => "10000001",12997 => "00011101",12998 => "11100001",12999 => "01110100",13000 => "10100111",13001 => "01111001",13002 => "00110100",13003 => "11111011",13004 => "00011100",13005 => "11011001",13006 => "00011111",13007 => "01111010",13008 => "10100110",13009 => "11101100",13010 => "10010000",13011 => "01110101",13012 => "00001011",13013 => "11001100",13014 => "01000001",13015 => "11010101",13016 => "01100100",13017 => "11000100",13018 => "01011000",13019 => "10011001",13020 => "10110110",13021 => "00111100",13022 => "10001011",13023 => "00110100",13024 => "11010110",13025 => "10010101",13026 => "10111110",13027 => "01101111",13028 => "00100000",13029 => "11111010",13030 => "00001111",13031 => "00001000",13032 => "11010101",13033 => "11001010",13034 => "10010101",13035 => "11101010",13036 => "00101000",13037 => "01010001",13038 => "11110001",13039 => "01010110",13040 => "10001001",13041 => "11110001",13042 => "01101111",13043 => "10001101",13044 => "00111100",13045 => "10101100",13046 => "00111100",13047 => "11010110",13048 => "01010101",13049 => "11111001",13050 => "01111010",13051 => "10010100",13052 => "00000110",13053 => "01011000",13054 => "01000010",13055 => "10101101",13056 => "10011010",13057 => "01101000",13058 => "00001011",13059 => "11010100",13060 => "10101000",13061 => "10110101",13062 => "00001100",13063 => "11111010",13064 => "11011001",13065 => "10001110",13066 => "01100001",13067 => "11101010",13068 => "11010111",13069 => "00011111",13070 => "10000100",13071 => "00111110",13072 => "00010101",13073 => "01110001",13074 => "10100011",13075 => "00010111",13076 => "00001011",13077 => "11011101",13078 => "11000000",13079 => "01110011",13080 => "11001000",13081 => "01111001",13082 => "00000100",13083 => "01001100",13084 => "01011100",13085 => "10101111",13086 => "00010111",13087 => "00011111",13088 => "00110110",13089 => "11101001",13090 => "00101010",13091 => "00010101",13092 => "11110010",13093 => "11010100",13094 => "10011001",13095 => "00101100",13096 => "00111101",13097 => "00111100",13098 => "00101101",13099 => "10110101",13100 => "11010001",13101 => "10000011",13102 => "01001000",13103 => "11001110",13104 => "01110111",13105 => "10101101",13106 => "10001101",13107 => "00111110",13108 => "10100011",13109 => "11100110",13110 => "10110100",13111 => "00001110",13112 => "00000101",13113 => "00110100",13114 => "00110011",13115 => "11101110",13116 => "00101001",13117 => "01111100",13118 => "00111001",13119 => "00110010",13120 => "00001110",13121 => "10001100",13122 => "00101111",13123 => "00100111",13124 => "01111100",13125 => "01001110",13126 => "01001000",13127 => "11111001",13128 => "01110100",13129 => "10101001",13130 => "00101100",13131 => "10101110",13132 => "10011110",13133 => "01010100",13134 => "00111101",13135 => "10100011",13136 => "01110110",13137 => "00000000",13138 => "10110101",13139 => "10111110",13140 => "01100100",13141 => "11011101",13142 => "01001110",13143 => "00000001",13144 => "11110011",13145 => "11101000",13146 => "10010101",13147 => "00100111",13148 => "00101011",13149 => "10000101",13150 => "01100100",13151 => "10010011",13152 => "10101011",13153 => "01111110",13154 => "01100011",13155 => "11011010",13156 => "01010011",13157 => "01111000",13158 => "11111010",13159 => "00010011",13160 => "00011011",13161 => "00011111",13162 => "11011010",13163 => "00110111",13164 => "10110010",13165 => "00101011",13166 => "00110101",13167 => "11110101",13168 => "01011111",13169 => "01110110",13170 => "00111110",13171 => "11110101",13172 => "10110100",13173 => "01111011",13174 => "11110000",13175 => "00011011",13176 => "00110100",13177 => "11001011",13178 => "01111001",13179 => "01101000",13180 => "00011110",13181 => "00011101",13182 => "01000101",13183 => "11101101",13184 => "00111110",13185 => "10000001",13186 => "11101110",13187 => "10100100",13188 => "10110000",13189 => "01000000",13190 => "00001001",13191 => "11000010",13192 => "01110111",13193 => "01011001",13194 => "10010100",13195 => "01000101",13196 => "00100011",13197 => "10101000",13198 => "00110110",13199 => "10011111",13200 => "11110100",13201 => "00011100",13202 => "00000011",13203 => "11011010",13204 => "01111100",13205 => "01011001",13206 => "10111110",13207 => "11010101",13208 => "10011100",13209 => "11000111",13210 => "01110110",13211 => "00001101",13212 => "01011011",13213 => "11001010",13214 => "01101101",13215 => "01010101",13216 => "10101100",13217 => "01001110",13218 => "01101011",13219 => "11101000",13220 => "10010011",13221 => "00111001",13222 => "10011010",13223 => "00111110",13224 => "00110101",13225 => "10000100",13226 => "11001101",13227 => "11000010",13228 => "01000101",13229 => "00101100",13230 => "00000000",13231 => "10001111",13232 => "01010100",13233 => "01110000",13234 => "10100000",13235 => "01010110",13236 => "10010101",13237 => "00011000",13238 => "10001010",13239 => "10101011",13240 => "01010100",13241 => "10111011",13242 => "01101001",13243 => "10011110",13244 => "11000100",13245 => "10111011",13246 => "00011100",13247 => "10000010",13248 => "10000001",13249 => "01101001",13250 => "00101111",13251 => "11010001",13252 => "10010001",13253 => "10000000",13254 => "11000010",13255 => "01111110",13256 => "11100001",13257 => "01100000",13258 => "10000111",13259 => "00000001",13260 => "00111010",13261 => "00010001",13262 => "00110001",13263 => "00101111",13264 => "11101100",13265 => "00100011",13266 => "10001011",13267 => "00001111",13268 => "01111001",13269 => "01000001",13270 => "11010011",13271 => "11010000",13272 => "10001000",13273 => "11010000",13274 => "10111001",13275 => "01000000",13276 => "01101100",13277 => "00010110",13278 => "10100001",13279 => "01111110",13280 => "01110001",13281 => "11000100",13282 => "11111010",13283 => "11011000",13284 => "00010001",13285 => "00101010",13286 => "00010001",13287 => "11000110",13288 => "10001010",13289 => "11001010",13290 => "01111001",13291 => "11101101",13292 => "11100111",13293 => "00111101",13294 => "01111001",13295 => "10001001",13296 => "10011010",13297 => "01111111",13298 => "00111100",13299 => "11101011",13300 => "00010110",13301 => "11000111",13302 => "10010010",13303 => "01110001",13304 => "01111000",13305 => "10100010",13306 => "11101011",13307 => "00001111",13308 => "10111110",13309 => "01111110",13310 => "01010111",13311 => "01010101",13312 => "11000010",13313 => "10101011",13314 => "01011111",13315 => "01101011",13316 => "10111100",13317 => "10110101",13318 => "00011101",13319 => "00111010",13320 => "11001100",13321 => "00000101",13322 => "10111110",13323 => "00101101",13324 => "10010101",13325 => "00110011",13326 => "11011011",13327 => "01001010",13328 => "11010011",13329 => "00010000",13330 => "01101100",13331 => "10000101",13332 => "01101100",13333 => "10111111",13334 => "01011111",13335 => "01010100",13336 => "11011111",13337 => "10010100",13338 => "00001100",13339 => "11100100",13340 => "00011110",13341 => "11000110",13342 => "10001110",13343 => "01111010",13344 => "11010111",13345 => "01100000",13346 => "11011100",13347 => "11000110",13348 => "10001101",13349 => "10011100",13350 => "01000001",13351 => "10001101",13352 => "00010111",13353 => "01100100",13354 => "11110010",13355 => "11101001",13356 => "00111010",13357 => "00111000",13358 => "00100111",13359 => "00110101",13360 => "11011100",13361 => "11000111",13362 => "11111000",13363 => "10001011",13364 => "01110000",13365 => "11001000",13366 => "00001111",13367 => "11100011",13368 => "11000100",13369 => "00011000",13370 => "10111111",13371 => "10001000",13372 => "11100000",13373 => "10111111",13374 => "00110101",13375 => "00011101",13376 => "11100110",13377 => "01000111",13378 => "00110000",13379 => "01101101",13380 => "10100101",13381 => "01101100",13382 => "00011000",13383 => "00001100",13384 => "00101101",13385 => "00010001",13386 => "10110111",13387 => "00000100",13388 => "11010000",13389 => "11111101",13390 => "10100001",13391 => "10111101",13392 => "01110101",13393 => "11000010",13394 => "10101011",13395 => "01110101",13396 => "01110001",13397 => "01100111",13398 => "00001001",13399 => "10010001",13400 => "00100100",13401 => "00000011",13402 => "11111101",13403 => "00101101",13404 => "00111100",13405 => "01101101",13406 => "10011111",13407 => "00000111",13408 => "01110011",13409 => "11011010",13410 => "00001011",13411 => "11101011",13412 => "10001001",13413 => "00110011",13414 => "11000111",13415 => "00001111",13416 => "01010101",13417 => "00100111",13418 => "00010011",13419 => "00100011",13420 => "00001010",13421 => "10011011",13422 => "10101101",13423 => "11010111",13424 => "10000011",13425 => "11101001",13426 => "10111011",13427 => "11111010",13428 => "01001001",13429 => "11011001",13430 => "11101010",13431 => "00111000",13432 => "11111100",13433 => "11011110",13434 => "10101010",13435 => "01100111",13436 => "00110000",13437 => "10000011",13438 => "11100000",13439 => "10100000",13440 => "01011110",13441 => "01010000",13442 => "00110010",13443 => "10111110",13444 => "00101001",13445 => "11111011",13446 => "01110100",13447 => "11000010",13448 => "01001001",13449 => "11100000",13450 => "11101010",13451 => "11011101",13452 => "10010010",13453 => "11100001",13454 => "00111111",13455 => "00011111",13456 => "10100110",13457 => "00110100",13458 => "00011001",13459 => "11011001",13460 => "10000101",13461 => "00011000",13462 => "10011011",13463 => "11011001",13464 => "01000010",13465 => "10001001",13466 => "11111010",13467 => "10010101",13468 => "00000010",13469 => "11001100",13470 => "10101010",13471 => "01111101",13472 => "01000000",13473 => "11110001",13474 => "10110110",13475 => "10111001",13476 => "01110100",13477 => "11110011",13478 => "00111000",13479 => "01011001",13480 => "11010000",13481 => "10100010",13482 => "11000010",13483 => "11111100",13484 => "10001110",13485 => "10111010",13486 => "00000011",13487 => "00000111",13488 => "00000110",13489 => "10100101",13490 => "00010001",13491 => "11111100",13492 => "10001111",13493 => "00011111",13494 => "11100111",13495 => "01110110",13496 => "01111100",13497 => "01111110",13498 => "11011100",13499 => "11000100",13500 => "01111000",13501 => "01111100",13502 => "10100100",13503 => "11101001",13504 => "00100000",13505 => "11100010",13506 => "01110001",13507 => "01111010",13508 => "10000001",13509 => "10110000",13510 => "11011001",13511 => "00010101",13512 => "00011001",13513 => "10010010",13514 => "10010100",13515 => "11100001",13516 => "10101110",13517 => "00010111",13518 => "00110011",13519 => "11101101",13520 => "10000111",13521 => "10111001",13522 => "01011110",13523 => "01111011",13524 => "00001010",13525 => "00010011",13526 => "10000101",13527 => "10111110",13528 => "01011111",13529 => "00000111",13530 => "00110010",13531 => "11110011",13532 => "01001110",13533 => "00001110",13534 => "10001100",13535 => "10011101",13536 => "01100111",13537 => "10010100",13538 => "10000101",13539 => "11111010",13540 => "11001111",13541 => "11010111",13542 => "01000101",13543 => "11000001",13544 => "10101010",13545 => "00110100",13546 => "01000101",13547 => "10010011",13548 => "11100010",13549 => "01001101",13550 => "11000101",13551 => "10100111",13552 => "00011101",13553 => "00110001",13554 => "11010111",13555 => "00011101",13556 => "10110000",13557 => "10111001",13558 => "01110010",13559 => "11100101",13560 => "00010100",13561 => "11100100",13562 => "00101111",13563 => "00000111",13564 => "11011111",13565 => "01111101",13566 => "11110101",13567 => "00101010",13568 => "11000110",13569 => "00100101",13570 => "11110001",13571 => "00011001",13572 => "00110100",13573 => "10110110",13574 => "10001111",13575 => "01001010",13576 => "00111110",13577 => "10000011",13578 => "01100010",13579 => "11001010",13580 => "01100001",13581 => "01000101",13582 => "00111000",13583 => "01010111",13584 => "00001000",13585 => "00000011",13586 => "10010100",13587 => "00110111",13588 => "01001110",13589 => "11100110",13590 => "00101100",13591 => "11010001",13592 => "10001110",13593 => "00100000",13594 => "01000000",13595 => "01100001",13596 => "01001101",13597 => "11110011",13598 => "11100011",13599 => "00111000",13600 => "11000111",13601 => "11001010",13602 => "01100010",13603 => "10011110",13604 => "10100110",13605 => "01001111",13606 => "10101000",13607 => "11011101",13608 => "00100011",13609 => "10011000",13610 => "00111110",13611 => "00111101",13612 => "00001111",13613 => "11000111",13614 => "10001100",13615 => "11101101",13616 => "01110110",13617 => "00110010",13618 => "00000111",13619 => "11010111",13620 => "11100100",13621 => "11011101",13622 => "01101111",13623 => "11001101",13624 => "10001100",13625 => "01100111",13626 => "00010001",13627 => "10010000",13628 => "00100011",13629 => "11111101",13630 => "10011100",13631 => "11000100",13632 => "11000101",13633 => "00100000",13634 => "11010001",13635 => "00001110",13636 => "00101110",13637 => "01100011",13638 => "10101001",13639 => "01100010",13640 => "00101011",13641 => "01011000",13642 => "10000110",13643 => "11011111",13644 => "10011000",13645 => "00101000",13646 => "01110111",13647 => "10111111",13648 => "10001011",13649 => "10000110",13650 => "01000000",13651 => "10001101",13652 => "11001001",13653 => "01111001",13654 => "11110101",13655 => "00100001",13656 => "11011111",13657 => "10001101",13658 => "00100010",13659 => "11110011",13660 => "01111100",13661 => "10001010",13662 => "00010100",13663 => "10111011",13664 => "10111010",13665 => "10111010",13666 => "00111010",13667 => "01101000",13668 => "11110111",13669 => "01011000",13670 => "10110111",13671 => "00101010",13672 => "01110011",13673 => "10000111",13674 => "11001100",13675 => "11110011",13676 => "10111011",13677 => "10001001",13678 => "11001101",13679 => "01101101",13680 => "10011110",13681 => "10011100",13682 => "01000010",13683 => "11101111",13684 => "11001011",13685 => "11011001",13686 => "11000011",13687 => "00010101",13688 => "11001110",13689 => "11111001",13690 => "01010111",13691 => "11111111",13692 => "10101011",13693 => "11110001",13694 => "11101111",13695 => "10010111",13696 => "01000000",13697 => "11011010",13698 => "01110100",13699 => "01001000",13700 => "01111111",13701 => "01010101",13702 => "10100110",13703 => "01000101",13704 => "01010000",13705 => "00001110",13706 => "01010101",13707 => "00010000",13708 => "00001000",13709 => "01000010",13710 => "10011001",13711 => "01110000",13712 => "11101100",13713 => "00101111",13714 => "01001010",13715 => "00000011",13716 => "00100011",13717 => "10101001",13718 => "10100101",13719 => "10010100",13720 => "00001110",13721 => "00111111",13722 => "00001000",13723 => "00111000",13724 => "11111001",13725 => "00010011",13726 => "11110111",13727 => "11101110",13728 => "10010010",13729 => "00100011",13730 => "11100111",13731 => "11000110",13732 => "01011110",13733 => "10010111",13734 => "01001000",13735 => "01001110",13736 => "11111011",13737 => "11110111",13738 => "10101100",13739 => "11000010",13740 => "01101011",13741 => "11000010",13742 => "10110111",13743 => "10101010",13744 => "10111001",13745 => "11101000",13746 => "10101110",13747 => "10011001",13748 => "01111000",13749 => "01001101",13750 => "11010111",13751 => "11100000",13752 => "11111110",13753 => "00101101",13754 => "11100110",13755 => "10110110",13756 => "00110111",13757 => "01001011",13758 => "01100000",13759 => "11000101",13760 => "00010111",13761 => "11011010",13762 => "01010110",13763 => "01011101",13764 => "11010000",13765 => "11100000",13766 => "01001000",13767 => "01011010",13768 => "10000011",13769 => "10110100",13770 => "01111001",13771 => "00011000",13772 => "00001101",13773 => "01010110",13774 => "10000000",13775 => "00010100",13776 => "11010110",13777 => "01010111",13778 => "11001011",13779 => "10111011",13780 => "00100011",13781 => "00001111",13782 => "00101001",13783 => "01011000",13784 => "10000011",13785 => "10100111",13786 => "11111110",13787 => "00111110",13788 => "00111000",13789 => "10111110",13790 => "01011110",13791 => "10011000",13792 => "00000010",13793 => "10000010",13794 => "10011100",13795 => "11101101",13796 => "10110111",13797 => "01000011",13798 => "01111111",13799 => "01110100",13800 => "11110111",13801 => "10010001",13802 => "10100111",13803 => "11101100",13804 => "00110100",13805 => "00110011",13806 => "00100001",13807 => "10011101",13808 => "10001011",13809 => "11111101",13810 => "11011011",13811 => "00101011",13812 => "01110111",13813 => "00110101",13814 => "10101010",13815 => "00000000",13816 => "01101110",13817 => "01101001",13818 => "01111111",13819 => "01111101",13820 => "01110011",13821 => "10101101",13822 => "11101010",13823 => "11111110",13824 => "00111001",13825 => "10101010",13826 => "00001011",13827 => "10110100",13828 => "11100011",13829 => "10111000",13830 => "00110100",13831 => "10001001",13832 => "00010110",13833 => "11011000",13834 => "01110010",13835 => "01101101",13836 => "01001000",13837 => "01010010",13838 => "11001100",13839 => "10100001",13840 => "11010111",13841 => "01011000",13842 => "00100011",13843 => "11110110",13844 => "01011110",13845 => "11111111",13846 => "10011100",13847 => "10101100",13848 => "11101101",13849 => "01011101",13850 => "11110000",13851 => "11110101",13852 => "01000001",13853 => "11100110",13854 => "01110010",13855 => "10101111",13856 => "11011111",13857 => "01000011",13858 => "10111100",13859 => "11010100",13860 => "10100101",13861 => "11100110",13862 => "10000001",13863 => "10110010",13864 => "11001100",13865 => "01100000",13866 => "11110000",13867 => "11101010",13868 => "10001001",13869 => "11111100",13870 => "00100001",13871 => "10110000",13872 => "01001010",13873 => "10010001",13874 => "00000011",13875 => "11000110",13876 => "00111010",13877 => "01010101",13878 => "01010110",13879 => "10101110",13880 => "00111010",13881 => "00010010",13882 => "00110001",13883 => "00110010",13884 => "11100011",13885 => "00111111",13886 => "11001110",13887 => "01011011",13888 => "10010100",13889 => "00100110",13890 => "10001010",13891 => "01000101",13892 => "10001101",13893 => "00101011",13894 => "10101001",13895 => "10010001",13896 => "11110001",13897 => "10100001",13898 => "11101101",13899 => "10000111",13900 => "01001000",13901 => "10101110",13902 => "10100010",13903 => "01010111",13904 => "11010110",13905 => "10110101",13906 => "10000001",13907 => "00001101",13908 => "01111011",13909 => "10100100",13910 => "10100000",13911 => "00011000",13912 => "10101010",13913 => "11010011",13914 => "11010000",13915 => "01110110",13916 => "01111001",13917 => "10000111",13918 => "11110111",13919 => "11011011",13920 => "01000000",13921 => "11001001",13922 => "10011011",13923 => "11101110",13924 => "10110111",13925 => "01111111",13926 => "00100011",13927 => "01001110",13928 => "00011100",13929 => "01011101",13930 => "11011010",13931 => "00100111",13932 => "10100011",13933 => "00111111",13934 => "11110010",13935 => "00111001",13936 => "01010110",13937 => "01110010",13938 => "01100110",13939 => "01000100",13940 => "11111100",13941 => "11111000",13942 => "00101011",13943 => "00101110",13944 => "00011110",13945 => "10110110",13946 => "11011110",13947 => "00111000",13948 => "00101110",13949 => "11001011",13950 => "01000000",13951 => "00111001",13952 => "01010100",13953 => "11101110",13954 => "00011101",13955 => "11010101",13956 => "01011111",13957 => "01101100",13958 => "00001111",13959 => "10101010",13960 => "00001011",13961 => "11001111",13962 => "10001011",13963 => "10001000",13964 => "00110111",13965 => "01000100",13966 => "10010011",13967 => "11010000",13968 => "00100101",13969 => "10010110",13970 => "01000100",13971 => "11001000",13972 => "00110100",13973 => "00011110",13974 => "01111000",13975 => "01100110",13976 => "00001000",13977 => "01010011",13978 => "00011010",13979 => "00010011",13980 => "00010010",13981 => "00010101",13982 => "01111101",13983 => "01100101",13984 => "11010111",13985 => "10111010",13986 => "11101010",13987 => "01110100",13988 => "01111010",13989 => "00011011",13990 => "00100100",13991 => "01100110",13992 => "00001100",13993 => "11010101",13994 => "01000011",13995 => "00110001",13996 => "01001110",13997 => "10011000",13998 => "10010110",13999 => "01010100",14000 => "01110110",14001 => "00000001",14002 => "10111111",14003 => "01011000",14004 => "00111111",14005 => "00110010",14006 => "01011101",14007 => "00100100",14008 => "01101011",14009 => "11001010",14010 => "10010110",14011 => "00101100",14012 => "11101101",14013 => "11010001",14014 => "10101001",14015 => "10011101",14016 => "10010010",14017 => "01101111",14018 => "11110011",14019 => "10101000",14020 => "01011010",14021 => "00011000",14022 => "00011101",14023 => "11001011",14024 => "00100011",14025 => "11110110",14026 => "10011110",14027 => "10101011",14028 => "10011000",14029 => "01001111",14030 => "01100001",14031 => "10011001",14032 => "01100011",14033 => "00101110",14034 => "11011000",14035 => "11101101",14036 => "11010010",14037 => "11011001",14038 => "11001011",14039 => "11011001",14040 => "11110100",14041 => "01010110",14042 => "11011110",14043 => "00010000",14044 => "01011011",14045 => "01010101",14046 => "11010111",14047 => "01011010",14048 => "11000000",14049 => "00101110",14050 => "01010100",14051 => "01110111",14052 => "01000000",14053 => "00001011",14054 => "00010000",14055 => "10001011",14056 => "10101111",14057 => "11001100",14058 => "11101011",14059 => "00110100",14060 => "11100101",14061 => "10101111",14062 => "11101001",14063 => "11100110",14064 => "10011010",14065 => "01000011",14066 => "11001011",14067 => "00010100",14068 => "01101001",14069 => "01101001",14070 => "00110010",14071 => "10110001",14072 => "11101110",14073 => "10100000",14074 => "01100010",14075 => "11011101",14076 => "10101011",14077 => "11010101",14078 => "11111000",14079 => "11111110",14080 => "11111001",14081 => "11001011",14082 => "01010111",14083 => "00111111",14084 => "11011010",14085 => "10110100",14086 => "11011010",14087 => "01111001",14088 => "00010001",14089 => "10011011",14090 => "00001100",14091 => "01011100",14092 => "01110011",14093 => "11110111",14094 => "10011100",14095 => "01111100",14096 => "00000111",14097 => "11000111",14098 => "01010011",14099 => "10011101",14100 => "11010010",14101 => "11001001",14102 => "00010000",14103 => "00011110",14104 => "11001110",14105 => "00111111",14106 => "00001010",14107 => "01111110",14108 => "00100001",14109 => "00001010",14110 => "01110010",14111 => "10000000",14112 => "11001011",14113 => "01000110",14114 => "11100100",14115 => "10110011",14116 => "00010001",14117 => "00110010",14118 => "11011000",14119 => "00100000",14120 => "11111000",14121 => "10110100",14122 => "00100111",14123 => "00111101",14124 => "00110100",14125 => "10111100",14126 => "00100001",14127 => "00010100",14128 => "11001101",14129 => "00101100",14130 => "10010101",14131 => "00101101",14132 => "00011100",14133 => "11110011",14134 => "11010011",14135 => "11000011",14136 => "10001100",14137 => "00100101",14138 => "00100010",14139 => "11110100",14140 => "00110111",14141 => "10000011",14142 => "01100011",14143 => "01110001",14144 => "01001001",14145 => "01001100",14146 => "00110101",14147 => "01010110",14148 => "00001110",14149 => "11100111",14150 => "01101110",14151 => "10111010",14152 => "10010001",14153 => "10100001",14154 => "00011001",14155 => "10010100",14156 => "00001100",14157 => "01110110",14158 => "00011000",14159 => "01001001",14160 => "00011100",14161 => "10101111",14162 => "11000101",14163 => "11100011",14164 => "00101010",14165 => "01011011",14166 => "11000111",14167 => "10010110",14168 => "11100000",14169 => "10011010",14170 => "10100001",14171 => "10101100",14172 => "11111110",14173 => "00011110",14174 => "00110101",14175 => "10110101",14176 => "10101000",14177 => "11111010",14178 => "10000100",14179 => "11011111",14180 => "00001011",14181 => "11100111",14182 => "01111100",14183 => "10110100",14184 => "01001001",14185 => "11011001",14186 => "01111000",14187 => "00001000",14188 => "01001011",14189 => "10100110",14190 => "01001101",14191 => "10001001",14192 => "10010111",14193 => "11011010",14194 => "11011111",14195 => "01000100",14196 => "01011010",14197 => "00100100",14198 => "01111010",14199 => "00011101",14200 => "11111001",14201 => "01111101",14202 => "01101000",14203 => "00011100",14204 => "10011010",14205 => "01100010",14206 => "01100010",14207 => "01000111",14208 => "00001110",14209 => "00110111",14210 => "10000000",14211 => "11100111",14212 => "00111110",14213 => "01110111",14214 => "00001111",14215 => "10111100",14216 => "00101110",14217 => "01111110",14218 => "11010101",14219 => "10110110",14220 => "00101000",14221 => "11011111",14222 => "00011001",14223 => "11011110",14224 => "11100111",14225 => "01000011",14226 => "01010001",14227 => "00100001",14228 => "01010101",14229 => "10000011",14230 => "10111110",14231 => "00110000",14232 => "11011001",14233 => "10001111",14234 => "00101110",14235 => "01101001",14236 => "00010011",14237 => "01111010",14238 => "11100000",14239 => "01001000",14240 => "01011111",14241 => "11101001",14242 => "11100110",14243 => "10100001",14244 => "01111000",14245 => "00001101",14246 => "10001110",14247 => "11111111",14248 => "01110111",14249 => "01000100",14250 => "10010101",14251 => "01110000",14252 => "00100010",14253 => "00001000",14254 => "11010101",14255 => "10111101",14256 => "11110110",14257 => "01101011",14258 => "00110001",14259 => "10111100",14260 => "10000101",14261 => "00011011",14262 => "01110010",14263 => "00100011",14264 => "10110100",14265 => "10001011",14266 => "01101000",14267 => "10010111",14268 => "10000101",14269 => "00000100",14270 => "11011010",14271 => "10010011",14272 => "01000100",14273 => "01100100",14274 => "10110011",14275 => "10011110",14276 => "11111111",14277 => "10111100",14278 => "11101011",14279 => "10010001",14280 => "00100101",14281 => "10001111",14282 => "10011010",14283 => "11001000",14284 => "01111011",14285 => "10011100",14286 => "10010000",14287 => "00011001",14288 => "00011011",14289 => "01111011",14290 => "11000001",14291 => "00101000",14292 => "10000010",14293 => "11000110",14294 => "01100010",14295 => "10000111",14296 => "10111010",14297 => "11011001",14298 => "11001110",14299 => "00101011",14300 => "00111001",14301 => "01001001",14302 => "11110101",14303 => "10111000",14304 => "00001010",14305 => "00011000",14306 => "11111000",14307 => "11000011",14308 => "01010110",14309 => "01111101",14310 => "11011001",14311 => "01110111",14312 => "01100101",14313 => "00110001",14314 => "11001111",14315 => "11101111",14316 => "01110000",14317 => "11001101",14318 => "01001100",14319 => "11100010",14320 => "01000100",14321 => "10011100",14322 => "01111110",14323 => "10101111",14324 => "01101111",14325 => "00010001",14326 => "11101111",14327 => "10101110",14328 => "10011100",14329 => "10101101",14330 => "01001111",14331 => "00010101",14332 => "10010100",14333 => "00011000",14334 => "11111101",14335 => "11010001",14336 => "01001110",14337 => "10110001",14338 => "10010011",14339 => "00000010",14340 => "11011101",14341 => "01100001",14342 => "00111010",14343 => "10111111",14344 => "01000001",14345 => "01111101",14346 => "00111101",14347 => "01110001",14348 => "01111010",14349 => "01000000",14350 => "11010100",14351 => "00000111",14352 => "00011010",14353 => "00110100",14354 => "10110111",14355 => "11001100",14356 => "01000011",14357 => "10101111",14358 => "00110010",14359 => "01010010",14360 => "11000011",14361 => "11010011",14362 => "01101010",14363 => "01111101",14364 => "10001000",14365 => "11101111",14366 => "10110000",14367 => "01010011",14368 => "11100111",14369 => "11010000",14370 => "11000101",14371 => "10100111",14372 => "00110010",14373 => "11011010",14374 => "11101101",14375 => "01000111",14376 => "10111100",14377 => "00110001",14378 => "10010101",14379 => "01110111",14380 => "10010100",14381 => "01000101",14382 => "00111000",14383 => "01011011",14384 => "00110011",14385 => "10110001",14386 => "00010111",14387 => "10110010",14388 => "10100111",14389 => "10011000",14390 => "00101111",14391 => "11000110",14392 => "10001110",14393 => "11001011",14394 => "11101111",14395 => "11110010",14396 => "01001100",14397 => "00001101",14398 => "10110111",14399 => "00010101",14400 => "00001111",14401 => "11111110",14402 => "10100000",14403 => "11010010",14404 => "10101110",14405 => "11111010",14406 => "11011110",14407 => "00110110",14408 => "10100100",14409 => "01110100",14410 => "11010101",14411 => "00001010",14412 => "10000110",14413 => "10001101",14414 => "01010110",14415 => "01010100",14416 => "01100101",14417 => "11000001",14418 => "01010110",14419 => "10001100",14420 => "00110110",14421 => "11101100",14422 => "10010010",14423 => "10011110",14424 => "00110100",14425 => "01001111",14426 => "01001011",14427 => "11100111",14428 => "11010000",14429 => "11101101",14430 => "10010011",14431 => "10100010",14432 => "11100101",14433 => "11110010",14434 => "11110001",14435 => "10011100",14436 => "10000110",14437 => "10100000",14438 => "01110001",14439 => "11000001",14440 => "10110111",14441 => "11100000",14442 => "11001111",14443 => "00111111",14444 => "10001101",14445 => "11011100",14446 => "11100011",14447 => "10001011",14448 => "01111101",14449 => "11001011",14450 => "00010001",14451 => "00101001",14452 => "01000111",14453 => "00010000",14454 => "01100110",14455 => "11111011",14456 => "00111001",14457 => "10001010",14458 => "10001000",14459 => "10101010",14460 => "11101110",14461 => "10011000",14462 => "00100110",14463 => "00001110",14464 => "01010001",14465 => "01001101",14466 => "10100101",14467 => "10010001",14468 => "00101100",14469 => "10110001",14470 => "01001010",14471 => "00101001",14472 => "00101110",14473 => "10000010",14474 => "10011000",14475 => "00001010",14476 => "00101010",14477 => "01010110",14478 => "00110111",14479 => "11101001",14480 => "10100000",14481 => "00011010",14482 => "01101010",14483 => "10001111",14484 => "10010110",14485 => "01011011",14486 => "11111010",14487 => "00010010",14488 => "01000110",14489 => "10001001",14490 => "10100110",14491 => "00100001",14492 => "01000011",14493 => "00111101",14494 => "11111000",14495 => "10011101",14496 => "01100011",14497 => "01110101",14498 => "11101001",14499 => "01101000",14500 => "00010011",14501 => "01111101",14502 => "01001010",14503 => "00001001",14504 => "01110001",14505 => "01111110",14506 => "00001010",14507 => "00011010",14508 => "10110010",14509 => "11011011",14510 => "01110110",14511 => "10101000",14512 => "11110011",14513 => "10100111",14514 => "11100000",14515 => "11101001",14516 => "11011111",14517 => "10000110",14518 => "10100101",14519 => "00001110",14520 => "01100001",14521 => "10110011",14522 => "00100111",14523 => "11100010",14524 => "01111011",14525 => "00010011",14526 => "11110010",14527 => "00110010",14528 => "00111001",14529 => "10100000",14530 => "10101011",14531 => "11010001",14532 => "01001101",14533 => "01110100",14534 => "10111000",14535 => "01010111",14536 => "10101101",14537 => "00110000",14538 => "11101010",14539 => "10110010",14540 => "00001001",14541 => "00000011",14542 => "00100100",14543 => "11110000",14544 => "10101101",14545 => "10011010",14546 => "01001000",14547 => "11111110",14548 => "10001010",14549 => "11101010",14550 => "01001010",14551 => "00101011",14552 => "11111110",14553 => "10110111",14554 => "00000010",14555 => "11000010",14556 => "01110001",14557 => "11011001",14558 => "00001110",14559 => "00010010",14560 => "00011000",14561 => "00110111",14562 => "10110011",14563 => "00110111",14564 => "10001001",14565 => "01100011",14566 => "10110000",14567 => "11010101",14568 => "00111110",14569 => "10000011",14570 => "11001101",14571 => "01010111",14572 => "11011001",14573 => "01101001",14574 => "00101001",14575 => "11001100",14576 => "11100011",14577 => "11001010",14578 => "11011010",14579 => "01001011",14580 => "11011100",14581 => "10111011",14582 => "11111011",14583 => "11111101",14584 => "10101101",14585 => "10111010",14586 => "10001001",14587 => "11011000",14588 => "00010000",14589 => "00111100",14590 => "11000001",14591 => "11101011",14592 => "01010100",14593 => "00011100",14594 => "11101001",14595 => "11101011",14596 => "10101111",14597 => "01011110",14598 => "01010100",14599 => "00110000",14600 => "01001110",14601 => "01000000",14602 => "00010100",14603 => "11100110",14604 => "10111011",14605 => "10110011",14606 => "01001001",14607 => "10111110",14608 => "01010110",14609 => "01000000",14610 => "00011100",14611 => "01010001",14612 => "00111110",14613 => "00000010",14614 => "10110000",14615 => "11001110",14616 => "00100101",14617 => "10100100",14618 => "01100100",14619 => "10101111",14620 => "00011000",14621 => "11011010",14622 => "00011010",14623 => "10110000",14624 => "10101100",14625 => "10001001",14626 => "11100110",14627 => "00010010",14628 => "01101110",14629 => "00111110",14630 => "10111010",14631 => "11101110",14632 => "10010100",14633 => "11110110",14634 => "10010111",14635 => "00100010",14636 => "10010111",14637 => "10101010",14638 => "00101100",14639 => "01111111",14640 => "10000110",14641 => "10110011",14642 => "01110001",14643 => "01000101",14644 => "01111001",14645 => "00111010",14646 => "10111110",14647 => "10001100",14648 => "01000101",14649 => "01001100",14650 => "00000000",14651 => "11010111",14652 => "11100000",14653 => "00100011",14654 => "10001100",14655 => "01001000",14656 => "11100011",14657 => "11000101",14658 => "11001010",14659 => "00110010",14660 => "10011001",14661 => "00100010",14662 => "10100110",14663 => "01100101",14664 => "01001011",14665 => "00010010",14666 => "00110111",14667 => "11111000",14668 => "11000111",14669 => "01010011",14670 => "00101111",14671 => "00000011",14672 => "10011001",14673 => "00100101",14674 => "11001100",14675 => "10111000",14676 => "01110110",14677 => "00100000",14678 => "00100101",14679 => "01011111",14680 => "00000001",14681 => "01101010",14682 => "10010010",14683 => "01110010",14684 => "01010101",14685 => "10000110",14686 => "01000000",14687 => "11000101",14688 => "00001111",14689 => "00000100",14690 => "11100000",14691 => "10100000",14692 => "00011111",14693 => "11110001",14694 => "10100000",14695 => "00111000",14696 => "01011011",14697 => "10000000",14698 => "00111110",14699 => "01110011",14700 => "11101100",14701 => "10110011",14702 => "10001110",14703 => "10011000",14704 => "11011001",14705 => "00110110",14706 => "11000101",14707 => "00100110",14708 => "10011101",14709 => "00001010",14710 => "11011010",14711 => "10100111",14712 => "11110100",14713 => "11101100",14714 => "10110101",14715 => "00000111",14716 => "01110011",14717 => "10011100",14718 => "10111010",14719 => "11101011",14720 => "10101001",14721 => "01101011",14722 => "10011001",14723 => "11100100",14724 => "11110000",14725 => "01010000",14726 => "10110101",14727 => "10000111",14728 => "01011111",14729 => "01100001",14730 => "00110000",14731 => "01011111",14732 => "10001010",14733 => "00011100",14734 => "11001001",14735 => "00001110",14736 => "10110111",14737 => "00101100",14738 => "10111010",14739 => "11000010",14740 => "00111101",14741 => "10001101",14742 => "00110010",14743 => "11010010",14744 => "00110100",14745 => "01000011",14746 => "00001011",14747 => "11010011",14748 => "10100001",14749 => "00100000",14750 => "01011001",14751 => "01000100",14752 => "01011011",14753 => "00000011",14754 => "10000000",14755 => "10100110",14756 => "11011011",14757 => "11100100",14758 => "01011010",14759 => "10111111",14760 => "00010011",14761 => "00101110",14762 => "00111111",14763 => "00010110",14764 => "01010101",14765 => "01011000",14766 => "00011001",14767 => "11111010",14768 => "00000011",14769 => "11101000",14770 => "00010010",14771 => "01000001",14772 => "00110100",14773 => "00010101",14774 => "11000111",14775 => "01111010",14776 => "00000010",14777 => "11101110",14778 => "00100111",14779 => "11101100",14780 => "10111011",14781 => "01100001",14782 => "00101000",14783 => "11111000",14784 => "10010001",14785 => "10101011",14786 => "01101011",14787 => "00010100",14788 => "11010001",14789 => "01101001",14790 => "10011111",14791 => "01000111",14792 => "00000111",14793 => "11110011",14794 => "11111111",14795 => "00110010",14796 => "11101111",14797 => "00000111",14798 => "10111110",14799 => "11000000",14800 => "01010110",14801 => "11001000",14802 => "01110100",14803 => "10011001",14804 => "01110100",14805 => "10010111",14806 => "00101011",14807 => "11100111",14808 => "11111001",14809 => "11110111",14810 => "00100111",14811 => "11011101",14812 => "01110011",14813 => "11011001",14814 => "00110100",14815 => "11100001",14816 => "11100011",14817 => "00001000",14818 => "10010100",14819 => "01000001",14820 => "10001101",14821 => "00011100",14822 => "00001100",14823 => "01000100",14824 => "01100000",14825 => "11000111",14826 => "10000000",14827 => "11011111",14828 => "10010000",14829 => "01001001",14830 => "01100111",14831 => "00101001",14832 => "10100001",14833 => "00001001",14834 => "11110000",14835 => "10011000",14836 => "11001100",14837 => "01110110",14838 => "01001010",14839 => "00101010",14840 => "10001000",14841 => "10100011",14842 => "11011101",14843 => "10101111",14844 => "11000100",14845 => "01100001",14846 => "00100111",14847 => "11001000",14848 => "00010011",14849 => "01110000",14850 => "10011111",14851 => "11001010",14852 => "01101001",14853 => "01000110",14854 => "00111010",14855 => "00101111",14856 => "00001001",14857 => "11110110",14858 => "11011011",14859 => "00110001",14860 => "01110101",14861 => "10111111",14862 => "11001110",14863 => "11110100",14864 => "11101111",14865 => "11011000",14866 => "01100100",14867 => "11011001",14868 => "01110011",14869 => "11110001",14870 => "11000111",14871 => "00111010",14872 => "11101000",14873 => "10110010",14874 => "00001101",14875 => "10110100",14876 => "00111010",14877 => "01001010",14878 => "00010010",14879 => "01111111",14880 => "11011001",14881 => "10100011",14882 => "00001000",14883 => "01110111",14884 => "10010110",14885 => "11011101",14886 => "11100010",14887 => "10000101",14888 => "11111100",14889 => "00001110",14890 => "01010000",14891 => "00011111",14892 => "01011001",14893 => "10110100",14894 => "11100000",14895 => "01100011",14896 => "01101000",14897 => "00101011",14898 => "00011100",14899 => "00110010",14900 => "00111110",14901 => "10111010",14902 => "10111101",14903 => "00011100",14904 => "00011011",14905 => "10100011",14906 => "11010001",14907 => "10100100",14908 => "01111001",14909 => "01010101",14910 => "00010001",14911 => "00011011",14912 => "00111010",14913 => "10011101",14914 => "10010111",14915 => "00001000",14916 => "01100000",14917 => "00111001",14918 => "10011111",14919 => "11100110",14920 => "10001011",14921 => "01111100",14922 => "11001111",14923 => "11111011",14924 => "01110110",14925 => "00111011",14926 => "10011001",14927 => "11010100",14928 => "00001100",14929 => "01110000",14930 => "10110010",14931 => "11100000",14932 => "11000000",14933 => "01100001",14934 => "11101110",14935 => "01110000",14936 => "01111100",14937 => "01000100",14938 => "00110100",14939 => "00011111",14940 => "11100110",14941 => "00011011",14942 => "00101010",14943 => "11111101",14944 => "01111111",14945 => "01110101",14946 => "00011010",14947 => "01100100",14948 => "00110100",14949 => "11101101",14950 => "00010011",14951 => "10100000",14952 => "10111010",14953 => "11000001",14954 => "00101101",14955 => "01000000",14956 => "10100110",14957 => "10111101",14958 => "10010011",14959 => "11100101",14960 => "00010100",14961 => "01011010",14962 => "10000001",14963 => "11001101",14964 => "10110000",14965 => "10101001",14966 => "10011111",14967 => "00101110",14968 => "00101101",14969 => "01111100",14970 => "00011110",14971 => "10010000",14972 => "11011111",14973 => "01100011",14974 => "10010011",14975 => "00100000",14976 => "00001011",14977 => "01111111",14978 => "01100000",14979 => "00010110",14980 => "10010011",14981 => "00010010",14982 => "00111010",14983 => "10001111",14984 => "00100011",14985 => "01100011",14986 => "00010011",14987 => "11111000",14988 => "11011110",14989 => "11101011",14990 => "01001011",14991 => "10101011",14992 => "01001010",14993 => "01010100",14994 => "01110101",14995 => "10000101",14996 => "00100110",14997 => "11001010",14998 => "00100111",14999 => "01011010",15000 => "00111111",15001 => "00101100",15002 => "11011000",15003 => "01011110",15004 => "10100000",15005 => "01100100",15006 => "01011011",15007 => "10101001",15008 => "01101011",15009 => "11011101",15010 => "11100110",15011 => "01001001",15012 => "00101001",15013 => "11100000",15014 => "11110101",15015 => "11001001",15016 => "11001000",15017 => "00111100",15018 => "10111100",15019 => "10000000",15020 => "10101100",15021 => "10101001",15022 => "00001111",15023 => "00111100",15024 => "01000010",15025 => "00000101",15026 => "11010110",15027 => "00101011",15028 => "11011100",15029 => "10010011",15030 => "10010100",15031 => "01011011",15032 => "00111000",15033 => "10001010",15034 => "11010000",15035 => "01110111",15036 => "00101001",15037 => "00001110",15038 => "01011011",15039 => "01001100",15040 => "10101100",15041 => "10011110",15042 => "01100000",15043 => "01111010",15044 => "01001101",15045 => "11101000",15046 => "10101100",15047 => "01000001",15048 => "10011100",15049 => "00100110",15050 => "00011011",15051 => "11010100",15052 => "01010001",15053 => "00010011",15054 => "01101001",15055 => "11110011",15056 => "11011101",15057 => "01100111",15058 => "10110011",15059 => "11001110",15060 => "10111011",15061 => "00011001",15062 => "10111011",15063 => "01010101",15064 => "01101110",15065 => "10010110",15066 => "10011001",15067 => "10001011",15068 => "10010010",15069 => "11000111",15070 => "00000100",15071 => "11111100",15072 => "01001001",15073 => "01001010",15074 => "00001000",15075 => "00010110",15076 => "00010101",15077 => "00011010",15078 => "10100111",15079 => "01001111",15080 => "00000111",15081 => "11000100",15082 => "00010110",15083 => "00000010",15084 => "01111100",15085 => "01010111",15086 => "01100110",15087 => "01110101",15088 => "00111011",15089 => "11110001",15090 => "00111010",15091 => "11000010",15092 => "00110110",15093 => "01000110",15094 => "00101110",15095 => "00101101",15096 => "01011001",15097 => "01110001",15098 => "01111100",15099 => "11111100",15100 => "01011000",15101 => "01010100",15102 => "00010101",15103 => "10000001",15104 => "11100100",15105 => "00100110",15106 => "11101001",15107 => "10000000",15108 => "10110010",15109 => "10110000",15110 => "00110100",15111 => "11010110",15112 => "11101100",15113 => "01101000",15114 => "11111101",15115 => "01011001",15116 => "10010100",15117 => "11101010",15118 => "01010011",15119 => "11111010",15120 => "10101110",15121 => "01000011",15122 => "10010110",15123 => "10111010",15124 => "00000011",15125 => "01101100",15126 => "00001000",15127 => "00101011",15128 => "01010000",15129 => "00011100",15130 => "10000000",15131 => "10011111",15132 => "10000011",15133 => "00101010",15134 => "10100101",15135 => "01101001",15136 => "11101001",15137 => "10100110",15138 => "10111001",15139 => "10010101",15140 => "11111011",15141 => "00100101",15142 => "11101001",15143 => "11011100",15144 => "00000110",15145 => "01011000",15146 => "10010000",15147 => "11010000",15148 => "00111100",15149 => "01001111",15150 => "11111000",15151 => "00011101",15152 => "11101011",15153 => "10111011",15154 => "01100111",15155 => "00111000",15156 => "01000110",15157 => "10001010",15158 => "11110110",15159 => "10110010",15160 => "11000011",15161 => "00101010",15162 => "10100001",15163 => "01111110",15164 => "10110111",15165 => "10111001",15166 => "11011101",15167 => "11111011",15168 => "01001010",15169 => "10010101",15170 => "00001011",15171 => "01100101",15172 => "00101111",15173 => "00101110",15174 => "10100101",15175 => "00011001",15176 => "10010001",15177 => "10010101",15178 => "11001110",15179 => "10011000",15180 => "01111010",15181 => "10000011",15182 => "01100100",15183 => "01010100",15184 => "10001100",15185 => "00001100",15186 => "10011010",15187 => "11011111",15188 => "11000010",15189 => "00010100",15190 => "10100100",15191 => "11101010",15192 => "10100111",15193 => "01101111",15194 => "00111110",15195 => "01000000",15196 => "10101001",15197 => "01100110",15198 => "00011000",15199 => "01001100",15200 => "00001111",15201 => "11100001",15202 => "10111000",15203 => "11100001",15204 => "00010110",15205 => "00101111",15206 => "00101110",15207 => "10010100",15208 => "01101111",15209 => "00101110",15210 => "11000110",15211 => "11010111",15212 => "11111010",15213 => "10001001",15214 => "10011110",15215 => "10000111",15216 => "00110110",15217 => "11010001",15218 => "10111000",15219 => "01101001",15220 => "01111000",15221 => "10010101",15222 => "11111101",15223 => "01101001",15224 => "01000101",15225 => "11110011",15226 => "00101010",15227 => "11001110",15228 => "10100010",15229 => "10101001",15230 => "00001000",15231 => "11101101",15232 => "10111011",15233 => "10100010",15234 => "01101010",15235 => "10111000",15236 => "00010110",15237 => "11010101",15238 => "11010011",15239 => "11100010",15240 => "10101111",15241 => "01100010",15242 => "01111110",15243 => "00101111",15244 => "10100101",15245 => "00011100",15246 => "00001001",15247 => "00011110",15248 => "00111110",15249 => "00010000",15250 => "01111111",15251 => "00011111",15252 => "01111110",15253 => "10011000",15254 => "00111001",15255 => "00110001",15256 => "00110000",15257 => "01101011",15258 => "01101010",15259 => "00010111",15260 => "11010100",15261 => "01010101",15262 => "10100001",15263 => "10001000",15264 => "11111101",15265 => "00001111",15266 => "00101010",15267 => "01100110",15268 => "01001111",15269 => "10110011",15270 => "11000010",15271 => "00101001",15272 => "00000010",15273 => "00011000",15274 => "11001010",15275 => "10011001",15276 => "00100010",15277 => "01000111",15278 => "00110100",15279 => "11110010",15280 => "10011100",15281 => "11001011",15282 => "10110111",15283 => "11001010",15284 => "01010000",15285 => "00110110",15286 => "01100111",15287 => "01111001",15288 => "11110100",15289 => "10100011",15290 => "00000111",15291 => "11011110",15292 => "10100000",15293 => "11111001",15294 => "10010111",15295 => "00110000",15296 => "01011001",15297 => "01001100",15298 => "11001100",15299 => "11000111",15300 => "10011010",15301 => "01110100",15302 => "01100111",15303 => "00111011",15304 => "11001001",15305 => "10110101",15306 => "01000011",15307 => "10101111",15308 => "01110011",15309 => "01111010",15310 => "01111100",15311 => "01010011",15312 => "10010010",15313 => "11001000",15314 => "01010000",15315 => "11011011",15316 => "00111101",15317 => "01001010",15318 => "10101010",15319 => "01101000",15320 => "01110111",15321 => "10110000",15322 => "00000001",15323 => "10000010",15324 => "01101100",15325 => "11100110",15326 => "10011101",15327 => "11001110",15328 => "01110110",15329 => "01000001",15330 => "10000010",15331 => "10010010",15332 => "10001011",15333 => "11110000",15334 => "10000000",15335 => "01011111",15336 => "00000101",15337 => "00000110",15338 => "11100010",15339 => "11000000",15340 => "00001111",15341 => "00011001",15342 => "00001100",15343 => "11001100",15344 => "11100110",15345 => "01100100",15346 => "10100010",15347 => "11100100",15348 => "11001111",15349 => "10100010",15350 => "00100000",15351 => "01010100",15352 => "10101110",15353 => "01101011",15354 => "11101001",15355 => "01100110",15356 => "10001000",15357 => "10101010",15358 => "00010110",15359 => "00010111",15360 => "10000010",15361 => "11111011",15362 => "01010111",15363 => "10100000",15364 => "10011000",15365 => "10001000",15366 => "10000100",15367 => "00000110",15368 => "10110011",15369 => "10010101",15370 => "11100001",15371 => "10001000",15372 => "01011111",15373 => "00011110",15374 => "10101010",15375 => "01110011",15376 => "00111001",15377 => "00100100",15378 => "10011101",15379 => "01000111",15380 => "11000011",15381 => "00010101",15382 => "01010110",15383 => "00000001",15384 => "00110100",15385 => "00101010",15386 => "11011110",15387 => "11001110",15388 => "10111011",15389 => "00111110",15390 => "00000110",15391 => "11000010",15392 => "01011110",15393 => "01111111",15394 => "11101001",15395 => "11000100",15396 => "01000111",15397 => "10110101",15398 => "11111011",15399 => "10100100",15400 => "11110001",15401 => "11100101",15402 => "11110100",15403 => "01010010",15404 => "00110100",15405 => "11101001",15406 => "11001110",15407 => "00101111",15408 => "11000000",15409 => "00001001",15410 => "00110001",15411 => "01011101",15412 => "01000000",15413 => "00001100",15414 => "00101000",15415 => "10001011",15416 => "10100010",15417 => "10010100",15418 => "01110010",15419 => "10111000",15420 => "00011010",15421 => "00010000",15422 => "01110110",15423 => "01010000",15424 => "01000010",15425 => "10001110",15426 => "10110011",15427 => "11111100",15428 => "00000101",15429 => "11100001",15430 => "10100100",15431 => "00110111",15432 => "11001011",15433 => "10100110",15434 => "11101010",15435 => "10110111",15436 => "10010000",15437 => "00100001",15438 => "10101010",15439 => "01011001",15440 => "10110001",15441 => "11111110",15442 => "10001100",15443 => "01110011",15444 => "11100011",15445 => "10011100",15446 => "00100001",15447 => "11000011",15448 => "01010010",15449 => "11110111",15450 => "00100110",15451 => "11101110",15452 => "11111000",15453 => "11001101",15454 => "11001011",15455 => "11101010",15456 => "00110011",15457 => "01101000",15458 => "01011011",15459 => "00111000",15460 => "11001011",15461 => "01101010",15462 => "00001011",15463 => "10010000",15464 => "10100101",15465 => "10101001",15466 => "10100000",15467 => "01000010",15468 => "00110011",15469 => "10010000",15470 => "01111011",15471 => "01100110",15472 => "10001001",15473 => "11011011",15474 => "10100101",15475 => "11010000",15476 => "11111001",15477 => "00001111",15478 => "00111100",15479 => "01101001",15480 => "01100001",15481 => "11010110",15482 => "11000101",15483 => "01011010",15484 => "11000011",15485 => "00001110",15486 => "10001011",15487 => "00011100",15488 => "00010110",15489 => "00111001",15490 => "01100000",15491 => "10110110",15492 => "00000110",15493 => "01101101",15494 => "11100101",15495 => "00100011",15496 => "10111011",15497 => "00010111",15498 => "01110001",15499 => "11101010",15500 => "11010111",15501 => "10100110",15502 => "11010000",15503 => "11100100",15504 => "10110110",15505 => "11001001",15506 => "11100101",15507 => "10111101",15508 => "00000101",15509 => "00111110",15510 => "10101011",15511 => "01001011",15512 => "00010000",15513 => "11100110",15514 => "11000011",15515 => "01110110",15516 => "00001100",15517 => "00110011",15518 => "10110001",15519 => "10010101",15520 => "00000001",15521 => "00110010",15522 => "00101110",15523 => "11101011",15524 => "00011101",15525 => "10010100",15526 => "10100011",15527 => "10000000",15528 => "11001110",15529 => "01011100",15530 => "11001111",15531 => "01000001",15532 => "11000110",15533 => "11010100",15534 => "11110101",15535 => "01001011",15536 => "01111111",15537 => "00101111",15538 => "01011101",15539 => "11110000",15540 => "00111010",15541 => "10100010",15542 => "11101001",15543 => "11111111",15544 => "01011101",15545 => "00101101",15546 => "01111111",15547 => "00010100",15548 => "10110111",15549 => "01100100",15550 => "01110100",15551 => "00010100",15552 => "00000110",15553 => "10010110",15554 => "01010001",15555 => "00110010",15556 => "00100011",15557 => "01010111",15558 => "01000010",15559 => "10000011",15560 => "00011111",15561 => "10100011",15562 => "00110011",15563 => "10011101",15564 => "00111000",15565 => "11101010",15566 => "01110111",15567 => "11011001",15568 => "10101111",15569 => "11010000",15570 => "00110000",15571 => "11100100",15572 => "00110000",15573 => "01001110",15574 => "11111000",15575 => "00010000",15576 => "01111101",15577 => "00101001",15578 => "10000100",15579 => "01110000",15580 => "00001011",15581 => "00010010",15582 => "01011011",15583 => "11101111",15584 => "10110100",15585 => "10011111",15586 => "10000010",15587 => "00001000",15588 => "01010001",15589 => "11000010",15590 => "01100010",15591 => "00010001",15592 => "00100110",15593 => "11101110",15594 => "01101111",15595 => "01101100",15596 => "11000000",15597 => "01111110",15598 => "11110110",15599 => "11010110",15600 => "01001011",15601 => "10011001",15602 => "01101011",15603 => "00111110",15604 => "01111101",15605 => "01100000",15606 => "00110110",15607 => "00011011",15608 => "10000101",15609 => "10110001",15610 => "11010110",15611 => "01100100",15612 => "01110010",15613 => "10101110",15614 => "00111000",15615 => "00000001",15616 => "11000011",15617 => "01101110",15618 => "10000110",15619 => "01000100",15620 => "01100000",15621 => "00100000",15622 => "01101101",15623 => "01000101",15624 => "10001000",15625 => "01011001",15626 => "11010001",15627 => "10101111",15628 => "00001111",15629 => "00001000",15630 => "00101011",15631 => "01110111",15632 => "01011000",15633 => "10001001",15634 => "10010011",15635 => "10011000",15636 => "11111011",15637 => "10111110",15638 => "10100111",15639 => "01100100",15640 => "11100101",15641 => "01110110",15642 => "01100011",15643 => "00101001",15644 => "00110101",15645 => "01010111",15646 => "11001110",15647 => "00100010",15648 => "10110101",15649 => "11110101",15650 => "10110010",15651 => "00000000",15652 => "01111011",15653 => "10101110",15654 => "01001100",15655 => "10101001",15656 => "10101101",15657 => "10001011",15658 => "01111111",15659 => "01101101",15660 => "00100101",15661 => "00111010",15662 => "01111111",15663 => "01101010",15664 => "10010011",15665 => "00110000",15666 => "11110000",15667 => "00110010",15668 => "00011011",15669 => "11110111",15670 => "10001011",15671 => "10111001",15672 => "10111001",15673 => "01001000",15674 => "01101100",15675 => "11101011",15676 => "01101001",15677 => "00011101",15678 => "11001111",15679 => "11010100",15680 => "01011011",15681 => "11111000",15682 => "11011011",15683 => "10000010",15684 => "01111000",15685 => "00110101",15686 => "00000010",15687 => "00110100",15688 => "00010100",15689 => "01100110",15690 => "10101010",15691 => "10100011",15692 => "10110100",15693 => "10101100",15694 => "01000010",15695 => "00001100",15696 => "11111111",15697 => "10010111",15698 => "01110001",15699 => "10101001",15700 => "11101001",15701 => "01000001",15702 => "01110101",15703 => "11101000",15704 => "00110100",15705 => "10011101",15706 => "10111100",15707 => "11010101",15708 => "11101111",15709 => "01001010",15710 => "01100111",15711 => "11010010",15712 => "10111001",15713 => "00111111",15714 => "10000011",15715 => "10100100",15716 => "01101010",15717 => "01100001",15718 => "10000100",15719 => "01010110",15720 => "10111010",15721 => "11011010",15722 => "11101011",15723 => "10101011",15724 => "00011111",15725 => "10101000",15726 => "01100101",15727 => "10010001",15728 => "00010011",15729 => "10100010",15730 => "00110111",15731 => "00010110",15732 => "10110010",15733 => "10110110",15734 => "10110100",15735 => "00001110",15736 => "10111011",15737 => "11110100",15738 => "10100110",15739 => "01011011",15740 => "11110111",15741 => "11100101",15742 => "11000111",15743 => "11010000",15744 => "11110111",15745 => "10111110",15746 => "00100111",15747 => "10000111",15748 => "10000111",15749 => "00111010",15750 => "11011111",15751 => "10010110",15752 => "10101101",15753 => "00001001",15754 => "01100110",15755 => "01011001",15756 => "11011100",15757 => "11101110",15758 => "11000101",15759 => "01101101",15760 => "01011110",15761 => "01100011",15762 => "10011000",15763 => "11100010",15764 => "01001011",15765 => "10000111",15766 => "01011010",15767 => "00011111",15768 => "01100001",15769 => "11110011",15770 => "10100111",15771 => "10100100",15772 => "00100011",15773 => "11000000",15774 => "01101001",15775 => "01111110",15776 => "11001111",15777 => "00000011",15778 => "11110000",15779 => "10010111",15780 => "10111001",15781 => "11101000",15782 => "00000110",15783 => "01100100",15784 => "00111110",15785 => "10100010",15786 => "11111010",15787 => "00100011",15788 => "11001110",15789 => "01000000",15790 => "00101100",15791 => "01101111",15792 => "01000101",15793 => "00000111",15794 => "10001000",15795 => "11111110",15796 => "11011100",15797 => "11011000",15798 => "11010111",15799 => "10001000",15800 => "00001010",15801 => "01011001",15802 => "11010000",15803 => "01010000",15804 => "10001100",15805 => "11010100",15806 => "01100011",15807 => "00101101",15808 => "11110110",15809 => "01011110",15810 => "01000011",15811 => "01011001",15812 => "10110001",15813 => "10101000",15814 => "01000110",15815 => "01011101",15816 => "11000110",15817 => "10100010",15818 => "00001001",15819 => "11011001",15820 => "01010000",15821 => "00010000",15822 => "01111010",15823 => "11001101",15824 => "01100011",15825 => "10011010",15826 => "01011100",15827 => "10101100",15828 => "11101111",15829 => "11100100",15830 => "00000010",15831 => "00111111",15832 => "00000110",15833 => "10110111",15834 => "00001001",15835 => "00100110",15836 => "01010001",15837 => "01001111",15838 => "01000101",15839 => "01010101",15840 => "10101110",15841 => "01111110",15842 => "01110110",15843 => "10110111",15844 => "10010001",15845 => "11001101",15846 => "01001000",15847 => "11110100",15848 => "11010101",15849 => "11000011",15850 => "11011000",15851 => "00011001",15852 => "00010101",15853 => "00011000",15854 => "10011111",15855 => "10011000",15856 => "11111101",15857 => "11111111",15858 => "11110011",15859 => "00110100",15860 => "10111001",15861 => "10110010",15862 => "00111011",15863 => "01100101",15864 => "01011100",15865 => "01000001",15866 => "00001101",15867 => "00100010",15868 => "11000001",15869 => "00010111",15870 => "10011001",15871 => "10001010",15872 => "11011101",15873 => "11111010",15874 => "11101011",15875 => "10011101",15876 => "10001010",15877 => "01101111",15878 => "00000011",15879 => "10111111",15880 => "10100011",15881 => "10101101",15882 => "01011110",15883 => "10110010",15884 => "11101101",15885 => "01010101",15886 => "10111100",15887 => "11101101",15888 => "11111101",15889 => "00111110",15890 => "00000110",15891 => "10111101",15892 => "11100001",15893 => "11101110",15894 => "11000111",15895 => "00101011",15896 => "11011111",15897 => "01111010",15898 => "00100000",15899 => "10111011",15900 => "11110111",15901 => "01101100",15902 => "00011011",15903 => "10010111",15904 => "10111011",15905 => "00011111",15906 => "00101011",15907 => "01000100",15908 => "00011101",15909 => "00011100",15910 => "11111110",15911 => "11001100",15912 => "10110111",15913 => "11100000",15914 => "01110011",15915 => "01010111",15916 => "10000011",15917 => "10111011",15918 => "11001100",15919 => "10100001",15920 => "01111000",15921 => "10010001",15922 => "00011101",15923 => "11010101",15924 => "00011111",15925 => "00110100",15926 => "00100110",15927 => "10010110",15928 => "00100000",15929 => "11101101",15930 => "00010010",15931 => "00000011",15932 => "01011110",15933 => "01111110",15934 => "11100101",15935 => "01000000",15936 => "00111101",15937 => "01110101",15938 => "01000101",15939 => "00111000",15940 => "01011100",15941 => "11011011",15942 => "01101101",15943 => "10101000",15944 => "00010010",15945 => "01101001",15946 => "11000111",15947 => "00001000",15948 => "00111001",15949 => "11111110",15950 => "10101110",15951 => "11110001",15952 => "00110100",15953 => "11110001",15954 => "00000011",15955 => "11111001",15956 => "10100101",15957 => "00000010",15958 => "11000000",15959 => "01010001",15960 => "11011101",15961 => "00110011",15962 => "10000010",15963 => "10010010",15964 => "01001111",15965 => "11110110",15966 => "00101101",15967 => "10111111",15968 => "00100011",15969 => "10001101",15970 => "00101010",15971 => "00011001",15972 => "11111000",15973 => "10000100",15974 => "01001010",15975 => "10101100",15976 => "01001001",15977 => "11101001",15978 => "11101100",15979 => "01111001",15980 => "11011001",15981 => "11100101",15982 => "11101100",15983 => "11000011",15984 => "11000001",15985 => "01110100",15986 => "11010001",15987 => "01110100",15988 => "00110010",15989 => "00100100",15990 => "10101111",15991 => "11101100",15992 => "11101011",15993 => "10000011",15994 => "01000100",15995 => "10000100",15996 => "11101011",15997 => "01011001",15998 => "10010010",15999 => "01100000",16000 => "01001000",16001 => "11100111",16002 => "11111110",16003 => "10110011",16004 => "01101111",16005 => "00101001",16006 => "11001101",16007 => "10001011",16008 => "01001100",16009 => "11000000",16010 => "01001100",16011 => "11101110",16012 => "10000010",16013 => "10011011",16014 => "10111111",16015 => "11111110",16016 => "00011110",16017 => "10111010",16018 => "00010010",16019 => "10010000",16020 => "10001100",16021 => "00000010",16022 => "00110010",16023 => "01000101",16024 => "11000110",16025 => "00100000",16026 => "11011110",16027 => "11110101",16028 => "01011101",16029 => "01001101",16030 => "10011110",16031 => "01001110",16032 => "10010011",16033 => "01010010",16034 => "01101100",16035 => "11001101",16036 => "10001010",16037 => "11000100",16038 => "11001000",16039 => "00000010",16040 => "10001101",16041 => "00100011",16042 => "01000010",16043 => "10111100",16044 => "11110011",16045 => "11001010",16046 => "11011000",16047 => "01101011",16048 => "01101010",16049 => "10100100",16050 => "10100001",16051 => "01101110",16052 => "11010111",16053 => "11000111",16054 => "00010101",16055 => "01100101",16056 => "00111100",16057 => "11001011",16058 => "00111100",16059 => "01011110",16060 => "11101101",16061 => "10010010",16062 => "00100000",16063 => "10100101",16064 => "10110110",16065 => "11011111",16066 => "01100010",16067 => "10110011",16068 => "00100111",16069 => "01011101",16070 => "10111001",16071 => "00101001",16072 => "00011111",16073 => "11011010",16074 => "10011100",16075 => "11110010",16076 => "00001101",16077 => "10001011",16078 => "11100101",16079 => "01010111",16080 => "11010100",16081 => "10101010",16082 => "01110001",16083 => "00001101",16084 => "01010111",16085 => "10011100",16086 => "00110010",16087 => "00011110",16088 => "11111110",16089 => "01110010",16090 => "00010101",16091 => "11010001",16092 => "00000111",16093 => "10001010",16094 => "00101011",16095 => "00010100",16096 => "10111110",16097 => "00001001",16098 => "00101100",16099 => "10110100",16100 => "00101000",16101 => "00000100",16102 => "11011111",16103 => "11110011",16104 => "10100100",16105 => "11100101",16106 => "01011111",16107 => "00001111",16108 => "00001111",16109 => "01011011",16110 => "00111010",16111 => "00100011",16112 => "00011011",16113 => "01001011",16114 => "10001011",16115 => "00001101",16116 => "10011000",16117 => "11101000",16118 => "01110001",16119 => "11100001",16120 => "11011001",16121 => "00110111",16122 => "11000011",16123 => "11010010",16124 => "00100010",16125 => "10011010",16126 => "00111010",16127 => "00110101",16128 => "01011110",16129 => "10000100",16130 => "11101001",16131 => "00110011",16132 => "01111010",16133 => "10010010",16134 => "01000100",16135 => "01111111",16136 => "00111100",16137 => "00101111",16138 => "10001011",16139 => "10000101",16140 => "01101010",16141 => "11111001",16142 => "10100110",16143 => "11100110",16144 => "00011011",16145 => "01000011",16146 => "00101111",16147 => "00100011",16148 => "10101010",16149 => "10000010",16150 => "11100011",16151 => "10110000",16152 => "11000000",16153 => "01101110",16154 => "11001001",16155 => "11111101",16156 => "10010111",16157 => "01111110",16158 => "10110010",16159 => "00100000",16160 => "00101010",16161 => "11010001",16162 => "00011100",16163 => "01101011",16164 => "00111111",16165 => "00001110",16166 => "10000110",16167 => "01011011",16168 => "10001000",16169 => "11100111",16170 => "11011110",16171 => "10101110",16172 => "11010110",16173 => "00111010",16174 => "11000111",16175 => "10000101",16176 => "11011100",16177 => "10101000",16178 => "10111100",16179 => "11101011",16180 => "11000111",16181 => "11101111",16182 => "01011101",16183 => "01000110",16184 => "00000010",16185 => "00111001",16186 => "11111111",16187 => "00101010",16188 => "10010101",16189 => "00010101",16190 => "00110011",16191 => "00100001",16192 => "11011100",16193 => "11010001",16194 => "00100011",16195 => "10010000",16196 => "00101110",16197 => "10010111",16198 => "00010011",16199 => "10000111",16200 => "11000011",16201 => "10101111",16202 => "11111111",16203 => "11100011",16204 => "10010100",16205 => "01110001",16206 => "00111100",16207 => "00111010",16208 => "10011011",16209 => "01011101",16210 => "11011100",16211 => "01011110",16212 => "01011000",16213 => "11011001",16214 => "00111000",16215 => "00000000",16216 => "01101011",16217 => "11001110",16218 => "01100110",16219 => "10010101",16220 => "01001101",16221 => "01110110",16222 => "11001001",16223 => "01101011",16224 => "01011111",16225 => "10011110",16226 => "11001000",16227 => "11101001",16228 => "11100101",16229 => "00111010",16230 => "10001101",16231 => "00110010",16232 => "10101101",16233 => "11101010",16234 => "11001000",16235 => "00101110",16236 => "01001010",16237 => "11100100",16238 => "10110100",16239 => "11010001",16240 => "10101000",16241 => "00100111",16242 => "01101111",16243 => "01000000",16244 => "01100111",16245 => "10110000",16246 => "00011101",16247 => "10111100",16248 => "11011010",16249 => "11101101",16250 => "00011000",16251 => "00001110",16252 => "10011111",16253 => "11101000",16254 => "00101100",16255 => "10001011",16256 => "00011000",16257 => "10111110",16258 => "00010101",16259 => "00101110",16260 => "10011101",16261 => "00100111",16262 => "10110110",16263 => "10000001",16264 => "11010101",16265 => "01111101",16266 => "11111001",16267 => "11000100",16268 => "11100100",16269 => "11100100",16270 => "10100000",16271 => "11111010",16272 => "01101000",16273 => "10010110",16274 => "00010101",16275 => "01011011",16276 => "10111101",16277 => "10110010",16278 => "01100100",16279 => "11111001",16280 => "11100011",16281 => "01111110",16282 => "10100011",16283 => "01100111",16284 => "11111111",16285 => "00001011",16286 => "01100000",16287 => "01101100",16288 => "10101000",16289 => "11101110",16290 => "01111001",16291 => "10111011",16292 => "11011000",16293 => "01110101",16294 => "01011010",16295 => "11100011",16296 => "11110100",16297 => "11010101",16298 => "11000011",16299 => "10011001",16300 => "10101111",16301 => "01111011",16302 => "00101110",16303 => "00000000",16304 => "10011001",16305 => "11010111",16306 => "01101101",16307 => "11111101",16308 => "00011001",16309 => "10110010",16310 => "11110010",16311 => "11111001",16312 => "10101100",16313 => "01010000",16314 => "11101101",16315 => "10010010",16316 => "11010101",16317 => "11100101",16318 => "11100111",16319 => "11000110",16320 => "11011110",16321 => "10110110",16322 => "11010100",16323 => "10000011",16324 => "01101101",16325 => "10100011",16326 => "11100010",16327 => "11100011",16328 => "10100011",16329 => "11110011",16330 => "10101001",16331 => "00111111",16332 => "11000110",16333 => "00101100",16334 => "10001000",16335 => "10010001",16336 => "01101111",16337 => "10110000",16338 => "10101110",16339 => "10110110",16340 => "11111100",16341 => "01110000",16342 => "01110111",16343 => "01000101",16344 => "11010000",16345 => "00100001",16346 => "01111101",16347 => "00010001",16348 => "00101111",16349 => "00110101",16350 => "01010000",16351 => "10100010",16352 => "01110010",16353 => "11000100",16354 => "01010110",16355 => "00011100",16356 => "11111110",16357 => "00010010",16358 => "11010010",16359 => "11001111",16360 => "01111110",16361 => "11010110",16362 => "11000110",16363 => "10111000",16364 => "00101111",16365 => "11101100",16366 => "01111011",16367 => "10100000",16368 => "11001010",16369 => "00101010",16370 => "11010100",16371 => "00010010",16372 => "01100010",16373 => "00011111",16374 => "00001000",16375 => "11001101",16376 => "01101110",16377 => "11010111",16378 => "11110111",16379 => "00010100",16380 => "10011000",16381 => "01011001",16382 => "10110011",16383 => "10111110",16384 => "11100000",16385 => "00000110",16386 => "01100011",16387 => "00011000",16388 => "00011000",16389 => "11101101",16390 => "10001100",16391 => "00101111",16392 => "11111001",16393 => "10110100",16394 => "10010100",16395 => "11111010",16396 => "11011001",16397 => "11101101",16398 => "10001000",16399 => "00111100",16400 => "00010010",16401 => "00011100",16402 => "01000110",16403 => "10100011",16404 => "00101010",16405 => "10101100",16406 => "01001100",16407 => "10111101",16408 => "11000110",16409 => "10011100",16410 => "10110101",16411 => "10110010",16412 => "10100101",16413 => "00100100",16414 => "01111011",16415 => "11100100",16416 => "00011000",16417 => "01001010",16418 => "10110011",16419 => "10001001",16420 => "00111111",16421 => "10010000",16422 => "01111001",16423 => "01101110",16424 => "00000110",16425 => "10111111",16426 => "11110001",16427 => "01101011",16428 => "00000001",16429 => "10011010",16430 => "00011101",16431 => "10010001",16432 => "11001101",16433 => "10010111",16434 => "00001101",16435 => "11001101",16436 => "11010000",16437 => "11001101",16438 => "00111000",16439 => "01010011",16440 => "11110111",16441 => "00100011",16442 => "10000001",16443 => "10011100",16444 => "01101000",16445 => "01010010",16446 => "10110000",16447 => "11010101",16448 => "11010101",16449 => "11000000",16450 => "01001001",16451 => "10000000",16452 => "10100001",16453 => "11110001",16454 => "01001110",16455 => "01000111",16456 => "11000100",16457 => "00100011",16458 => "01011110",16459 => "01001100",16460 => "11111001",16461 => "11010110",16462 => "10000001",16463 => "00000011",16464 => "00001001",16465 => "01101011",16466 => "10001011",16467 => "10000100",16468 => "00111100",16469 => "00010110",16470 => "01111000",16471 => "01111101",16472 => "10111101",16473 => "01110000",16474 => "00010100",16475 => "01010001",16476 => "11010111",16477 => "11100001",16478 => "00011001",16479 => "01011100",16480 => "00011001",16481 => "10011011",16482 => "11100101",16483 => "00001110",16484 => "10101100",16485 => "00100110",16486 => "11111111",16487 => "01101011",16488 => "10101101",16489 => "11011101",16490 => "00100001",16491 => "11001011",16492 => "00110111",16493 => "01110101",16494 => "01100010",16495 => "10000101",16496 => "01101011",16497 => "01000001",16498 => "00100101",16499 => "01110110",16500 => "11110011",16501 => "10010001",16502 => "01010101",16503 => "11100110",16504 => "11111111",16505 => "11100111",16506 => "10011100",16507 => "11010000",16508 => "11100001",16509 => "10010101",16510 => "10110111",16511 => "01100101",16512 => "10001101",16513 => "01010111",16514 => "01011111",16515 => "10101100",16516 => "01001001",16517 => "01101011",16518 => "00011011",16519 => "00000001",16520 => "00100010",16521 => "00000111",16522 => "01111111",16523 => "10011011",16524 => "10100100",16525 => "11000011",16526 => "00110101",16527 => "00011101",16528 => "10011110",16529 => "11100110",16530 => "01000100",16531 => "00011001",16532 => "01011101",16533 => "10011000",16534 => "00001110",16535 => "11001001",16536 => "10110101",16537 => "10101000",16538 => "01010100",16539 => "01001101",16540 => "01100101",16541 => "01011101",16542 => "01000011",16543 => "10110001",16544 => "00010100",16545 => "11101011",16546 => "10110010",16547 => "11100100",16548 => "00010100",16549 => "10110111",16550 => "10100100",16551 => "10111101",16552 => "10001000",16553 => "11011011",16554 => "11111000",16555 => "01110100",16556 => "00111011",16557 => "01111100",16558 => "11010101",16559 => "00011001",16560 => "10111001",16561 => "01111011",16562 => "11101110",16563 => "10110010",16564 => "00111101",16565 => "11101000",16566 => "00100010",16567 => "00101001",16568 => "11101111",16569 => "10011110",16570 => "10101001",16571 => "01001101",16572 => "10011010",16573 => "10100011",16574 => "01010000",16575 => "11011011",16576 => "10001001",16577 => "11011100",16578 => "10010101",16579 => "10000111",16580 => "10001100",16581 => "11011011",16582 => "00011010",16583 => "00000001",16584 => "10010110",16585 => "01111010",16586 => "11010011",16587 => "01101100",16588 => "01101101",16589 => "00111110",16590 => "01011010",16591 => "01011001",16592 => "11100010",16593 => "00001001",16594 => "10011110",16595 => "00011101",16596 => "01011100",16597 => "01110001",16598 => "01111011",16599 => "00011101",16600 => "11001000",16601 => "00101011",16602 => "10001001",16603 => "10000000",16604 => "10110111",16605 => "00010110",16606 => "10001011",16607 => "10100100",16608 => "00111010",16609 => "11001000",16610 => "11101100",16611 => "00011111",16612 => "11000100",16613 => "11110000",16614 => "10111100",16615 => "11111110",16616 => "01110011",16617 => "00010000",16618 => "10010011",16619 => "01001100",16620 => "01001101",16621 => "01011011",16622 => "00000011",16623 => "10011111",16624 => "11011011",16625 => "01000010",16626 => "11110011",16627 => "11101000",16628 => "01001001",16629 => "10101000",16630 => "00000011",16631 => "10110001",16632 => "01101000",16633 => "10100001",16634 => "11001010",16635 => "10110011",16636 => "01100000",16637 => "00101100",16638 => "01111011",16639 => "10100001",16640 => "01011001",16641 => "01000100",16642 => "00011001",16643 => "10011111",16644 => "00001111",16645 => "11000110",16646 => "10011010",16647 => "11000111",16648 => "10001011",16649 => "00011101",16650 => "01010000",16651 => "10001000",16652 => "11101010",16653 => "10011111",16654 => "11010010",16655 => "11010010",16656 => "11011010",16657 => "10111001",16658 => "10001011",16659 => "00010111",16660 => "10101010",16661 => "11101011",16662 => "10010110",16663 => "10010101",16664 => "00000011",16665 => "11110011",16666 => "11101001",16667 => "01101010",16668 => "11100101",16669 => "00000011",16670 => "11000000",16671 => "10011010",16672 => "11100010",16673 => "11110110",16674 => "11000101",16675 => "10010001",16676 => "01001011",16677 => "11100101",16678 => "11101001",16679 => "10011111",16680 => "11100101",16681 => "10100011",16682 => "01001111",16683 => "11011110",16684 => "01011011",16685 => "11000100",16686 => "11101000",16687 => "11010000",16688 => "00011110",16689 => "10100011",16690 => "10010001",16691 => "10011111",16692 => "01111101",16693 => "01110011",16694 => "11111001",16695 => "01111110",16696 => "11010011",16697 => "00011101",16698 => "00000101",16699 => "00111100",16700 => "00011101",16701 => "11111100",16702 => "01100000",16703 => "11111101",16704 => "00111110",16705 => "10001000",16706 => "10111001",16707 => "01100110",16708 => "10011010",16709 => "01010110",16710 => "10110001",16711 => "00011011",16712 => "11111110",16713 => "01001110",16714 => "00001100",16715 => "11100100",16716 => "10010100",16717 => "01111101",16718 => "01010001",16719 => "01001101",16720 => "01111010",16721 => "00111101",16722 => "00001110",16723 => "00110111",16724 => "01100011",16725 => "10010101",16726 => "10001000",16727 => "01101110",16728 => "11000011",16729 => "00111000",16730 => "00100010",16731 => "10100010",16732 => "10111011",16733 => "00110001",16734 => "11100000",16735 => "01101000",16736 => "10101110",16737 => "10101111",16738 => "10111110",16739 => "00010100",16740 => "10101110",16741 => "10100110",16742 => "00011100",16743 => "00110110",16744 => "10111100",16745 => "10011110",16746 => "00101100",16747 => "01101101",16748 => "10100111",16749 => "01011100",16750 => "11001011",16751 => "11111011",16752 => "00011001",16753 => "00101001",16754 => "10110010",16755 => "00010100",16756 => "00010000",16757 => "10010011",16758 => "11101100",16759 => "10001101",16760 => "01000011",16761 => "01010111",16762 => "00010000",16763 => "10111011",16764 => "01001101",16765 => "01110011",16766 => "10101000",16767 => "00110100",16768 => "00011011",16769 => "00100001",16770 => "10110000",16771 => "10000110",16772 => "11111011",16773 => "00110010",16774 => "01001000",16775 => "00010101",16776 => "11101000",16777 => "01100101",16778 => "11000110",16779 => "01101000",16780 => "11101000",16781 => "01000100",16782 => "00101101",16783 => "00100111",16784 => "01101101",16785 => "10000100",16786 => "01000100",16787 => "10110001",16788 => "10010101",16789 => "01110001",16790 => "11100110",16791 => "10010001",16792 => "01011101",16793 => "00110100",16794 => "11010101",16795 => "00100110",16796 => "01001100",16797 => "00000110",16798 => "01110010",16799 => "00101101",16800 => "01101001",16801 => "00101000",16802 => "11001111",16803 => "01110111",16804 => "00011011",16805 => "00010100",16806 => "10010111",16807 => "01100101",16808 => "11111000",16809 => "00011001",16810 => "00000101",16811 => "00100000",16812 => "01100000",16813 => "10000110",16814 => "00111011",16815 => "00111011",16816 => "01010011",16817 => "01111100",16818 => "00111110",16819 => "10110010",16820 => "10100010",16821 => "10001011",16822 => "11101011",16823 => "11000010",16824 => "10010010",16825 => "01110000",16826 => "00101110",16827 => "11001000",16828 => "00010001",16829 => "01110001",16830 => "01101101",16831 => "10000010",16832 => "01010100",16833 => "00011110",16834 => "11001110",16835 => "11000010",16836 => "10010110",16837 => "11110011",16838 => "11010110",16839 => "10010100",16840 => "10011100",16841 => "01000100",16842 => "01001001",16843 => "01101110",16844 => "11110001",16845 => "10011001",16846 => "11011100",16847 => "11100000",16848 => "10001011",16849 => "11110000",16850 => "00010111",16851 => "00010110",16852 => "10000101",16853 => "10011001",16854 => "00111000",16855 => "01000100",16856 => "01000110",16857 => "01111100",16858 => "11000010",16859 => "11000010",16860 => "00011111",16861 => "01101110",16862 => "10000010",16863 => "01010011",16864 => "11110000",16865 => "11110011",16866 => "10101000",16867 => "00101110",16868 => "00000101",16869 => "11000011",16870 => "00001100",16871 => "00111101",16872 => "00000100",16873 => "00001110",16874 => "10011100",16875 => "01010001",16876 => "11111110",16877 => "01111100",16878 => "10100000",16879 => "01101011",16880 => "11101010",16881 => "01100101",16882 => "11011110",16883 => "10100000",16884 => "10100010",16885 => "00010101",16886 => "11101010",16887 => "11010011",16888 => "01011011",16889 => "01010101",16890 => "01100011",16891 => "11000101",16892 => "10110000",16893 => "00000101",16894 => "11011011",16895 => "10000111",16896 => "01011010",16897 => "11010101",16898 => "10000000",16899 => "10101010",16900 => "10100100",16901 => "10100011",16902 => "01110100",16903 => "10011010",16904 => "10101100",16905 => "00110010",16906 => "01110011",16907 => "10011111",16908 => "00100000",16909 => "00011011",16910 => "00011011",16911 => "00100011",16912 => "11110001",16913 => "11000110",16914 => "01111111",16915 => "10110110",16916 => "10100100",16917 => "11001000",16918 => "00000100",16919 => "11001000",16920 => "10011100",16921 => "10111110",16922 => "11101001",16923 => "00100101",16924 => "11110011",16925 => "00101001",16926 => "01011010",16927 => "00010010",16928 => "00000001",16929 => "10001100",16930 => "10111111",16931 => "11100111",16932 => "10110100",16933 => "10000110",16934 => "01010100",16935 => "00011001",16936 => "11001100",16937 => "01111101",16938 => "10010010",16939 => "11101001",16940 => "00110101",16941 => "11011010",16942 => "11010011",16943 => "11111110",16944 => "01111000",16945 => "00100011",16946 => "10001111",16947 => "01100101",16948 => "10001111",16949 => "00011100",16950 => "11010011",16951 => "00010100",16952 => "00010110",16953 => "01011001",16954 => "00100000",16955 => "01001001",16956 => "00111110",16957 => "10101010",16958 => "01111101",16959 => "11010110",16960 => "11100000",16961 => "11010000",16962 => "01100111",16963 => "11101011",16964 => "00000000",16965 => "10010011",16966 => "10001000",16967 => "00010011",16968 => "00101001",16969 => "10011100",16970 => "00111101",16971 => "10110011",16972 => "00111010",16973 => "00111000",16974 => "01001011",16975 => "00100000",16976 => "01000110",16977 => "11101111",16978 => "00010110",16979 => "00000000",16980 => "00100000",16981 => "00100111",16982 => "10100110",16983 => "11100011",16984 => "11010010",16985 => "00011010",16986 => "10110011",16987 => "10001011",16988 => "00110110",16989 => "10110111",16990 => "11101110",16991 => "00101011",16992 => "01000011",16993 => "11000000",16994 => "00001011",16995 => "10001011",16996 => "00101111",16997 => "00100011",16998 => "00101111",16999 => "00111100",17000 => "00011110",17001 => "00000110",17002 => "00010000",17003 => "11100010",17004 => "00000101",17005 => "11010100",17006 => "11010101",17007 => "01100001",17008 => "00001011",17009 => "10000001",17010 => "11110110",17011 => "11110110",17012 => "11111011",17013 => "00101001",17014 => "00101100",17015 => "01100011",17016 => "11010100",17017 => "01011110",17018 => "01111010",17019 => "11010110",17020 => "10110011",17021 => "00001110",17022 => "10100111",17023 => "01011100",17024 => "01011011",17025 => "00110000",17026 => "01010000",17027 => "11001100",17028 => "00110111",17029 => "11111011",17030 => "10001110",17031 => "00110011",17032 => "11101000",17033 => "01101001",17034 => "00101101",17035 => "00100111",17036 => "10000110",17037 => "01000111",17038 => "10000111",17039 => "11101101",17040 => "00110010",17041 => "10000010",17042 => "01100000",17043 => "11010000",17044 => "01110110",17045 => "00101100",17046 => "11100111",17047 => "11111000",17048 => "00001011",17049 => "11001001",17050 => "11110111",17051 => "10101100",17052 => "00110011",17053 => "01001101",17054 => "00010110",17055 => "10111111",17056 => "10011101",17057 => "10100001",17058 => "00000000",17059 => "01110010",17060 => "01010110",17061 => "11111011",17062 => "01111010",17063 => "00000110",17064 => "11011101",17065 => "01101010",17066 => "00111100",17067 => "01011111",17068 => "01101011",17069 => "01000001",17070 => "01010000",17071 => "00010100",17072 => "00101111",17073 => "00010001",17074 => "11110101",17075 => "00111110",17076 => "01010010",17077 => "11001011",17078 => "01011110",17079 => "11111101",17080 => "10101001",17081 => "10010100",17082 => "01111010",17083 => "01101010",17084 => "10001100",17085 => "01111111",17086 => "01010000",17087 => "10000000",17088 => "00000101",17089 => "11110101",17090 => "00011110",17091 => "00001001",17092 => "11011111",17093 => "00101101",17094 => "01010001",17095 => "01011011",17096 => "01111000",17097 => "01111011",17098 => "10111111",17099 => "11110110",17100 => "00110110",17101 => "11101000",17102 => "00010101",17103 => "00000111",17104 => "01101100",17105 => "00001110",17106 => "01000110",17107 => "01010010",17108 => "00101000",17109 => "01010001",17110 => "00111110",17111 => "01011001",17112 => "11101001",17113 => "10000111",17114 => "00011010",17115 => "11100111",17116 => "11110011",17117 => "01011111",17118 => "00110111",17119 => "00110111",17120 => "11100101",17121 => "01010011",17122 => "11010001",17123 => "10101000",17124 => "10010001",17125 => "11011110",17126 => "00001110",17127 => "10101110",17128 => "01011010",17129 => "11001001",17130 => "00000101",17131 => "00111100",17132 => "10010101",17133 => "10101000",17134 => "11101111",17135 => "10001100",17136 => "10011111",17137 => "10010110",17138 => "11000011",17139 => "10101011",17140 => "00000001",17141 => "00101001",17142 => "00101111",17143 => "10110110",17144 => "10100000",17145 => "00100000",17146 => "11101010",17147 => "00000010",17148 => "00110110",17149 => "00011010",17150 => "01011010",17151 => "11010101",17152 => "10101100",17153 => "11000100",17154 => "10000100",17155 => "11100000",17156 => "11101011",17157 => "10111000",17158 => "10100011",17159 => "01000011",17160 => "00101001",17161 => "00010000",17162 => "00101000",17163 => "01001101",17164 => "01110110",17165 => "11001111",17166 => "00101000",17167 => "10111011",17168 => "10000110",17169 => "11100110",17170 => "01100110",17171 => "01100101",17172 => "00100111",17173 => "10000111",17174 => "10110111",17175 => "01111010",17176 => "00011111",17177 => "01010111",17178 => "00100000",17179 => "01100011",17180 => "10000000",17181 => "10011110",17182 => "10101001",17183 => "11000000",17184 => "01010110",17185 => "01101111",17186 => "11100000",17187 => "00000011",17188 => "00101000",17189 => "00011110",17190 => "00110111",17191 => "00100001",17192 => "10100110",17193 => "01011111",17194 => "01101010",17195 => "00101101",17196 => "11010111",17197 => "11011011",17198 => "11010010",17199 => "11001110",17200 => "00000101",17201 => "11100111",17202 => "01010101",17203 => "10011000",17204 => "11101010",17205 => "10110101",17206 => "01000111",17207 => "01110111",17208 => "11110011",17209 => "00100011",17210 => "11101110",17211 => "10101011",17212 => "11000100",17213 => "11100101",17214 => "10011010",17215 => "10001111",17216 => "00100011",17217 => "11000010",17218 => "01000100",17219 => "00011001",17220 => "10111000",17221 => "11110000",17222 => "00110101",17223 => "01111101",17224 => "11110010",17225 => "00011101",17226 => "00110010",17227 => "01101101",17228 => "11100100",17229 => "00000101",17230 => "11011111",17231 => "01100010",17232 => "00101100",17233 => "11000001",17234 => "10110111",17235 => "11111110",17236 => "11011011",17237 => "11011110",17238 => "11110001",17239 => "01100110",17240 => "00000000",17241 => "00110010",17242 => "10010100",17243 => "01010110",17244 => "11101100",17245 => "01110011",17246 => "11011111",17247 => "11001010",17248 => "01111110",17249 => "00100001",17250 => "10001001",17251 => "10100110",17252 => "10111110",17253 => "10100111",17254 => "10110001",17255 => "11011110",17256 => "11010001",17257 => "00001011",17258 => "11110011",17259 => "01110100",17260 => "11101011",17261 => "10111101",17262 => "01010111",17263 => "01111110",17264 => "00001000",17265 => "00010110",17266 => "11010110",17267 => "00010110",17268 => "00101001",17269 => "00000000",17270 => "00011110",17271 => "10010100",17272 => "01110010",17273 => "01000101",17274 => "01111110",17275 => "00010101",17276 => "01100100",17277 => "00001010",17278 => "11100011",17279 => "01011101",17280 => "10011000",17281 => "11101000",17282 => "10011011",17283 => "00001001",17284 => "00011111",17285 => "01111101",17286 => "11011110",17287 => "00110001",17288 => "10100101",17289 => "00011011",17290 => "11001011",17291 => "11101010",17292 => "01011000",17293 => "10000000",17294 => "01001000",17295 => "11100011",17296 => "10001100",17297 => "01001101",17298 => "01101111",17299 => "01011100",17300 => "11110011",17301 => "11000111",17302 => "00110000",17303 => "00011001",17304 => "01000011",17305 => "01111110",17306 => "00101101",17307 => "01011001",17308 => "00011011",17309 => "10010010",17310 => "11010010",17311 => "01111101",17312 => "10100111",17313 => "01001111",17314 => "01101001",17315 => "00101101",17316 => "11101111",17317 => "10010100",17318 => "11011011",17319 => "10110001",17320 => "10101101",17321 => "00010110",17322 => "01001101",17323 => "11100010",17324 => "11010110",17325 => "01110011",17326 => "11011011",17327 => "10011010",17328 => "11011111",17329 => "11000101",17330 => "11100101",17331 => "11101111",17332 => "11010000",17333 => "10011101",17334 => "00010000",17335 => "00010110",17336 => "10011110",17337 => "11000100",17338 => "11011110",17339 => "00100110",17340 => "10101001",17341 => "10001010",17342 => "00011110",17343 => "01010100",17344 => "11001011",17345 => "11000101",17346 => "10111101",17347 => "00100110",17348 => "11000110",17349 => "00000011",17350 => "01001000",17351 => "10111011",17352 => "01110111",17353 => "11110101",17354 => "11110011",17355 => "01110011",17356 => "11000011",17357 => "10000110",17358 => "00111110",17359 => "11110001",17360 => "11011110",17361 => "01000100",17362 => "01001100",17363 => "10101010",17364 => "11010110",17365 => "10000001",17366 => "11111001",17367 => "00111110",17368 => "00011101",17369 => "00010100",17370 => "10011101",17371 => "00110001",17372 => "10001010",17373 => "00001011",17374 => "00100101",17375 => "11100011",17376 => "01000001",17377 => "10101011",17378 => "00001011",17379 => "10000000",17380 => "10000001",17381 => "11101010",17382 => "11101011",17383 => "10000111",17384 => "01010101",17385 => "00111110",17386 => "00101010",17387 => "00010111",17388 => "11000110",17389 => "10001101",17390 => "10011001",17391 => "00001111",17392 => "00000101",17393 => "01011110",17394 => "01001010",17395 => "11100010",17396 => "10110000",17397 => "01100110",17398 => "01100101",17399 => "01001100",17400 => "01100100",17401 => "11110011",17402 => "00110011",17403 => "11110000",17404 => "00101001",17405 => "00110000",17406 => "00100010",17407 => "10101101",17408 => "11111001",17409 => "01010001",17410 => "01100011",17411 => "11101001",17412 => "10010000",17413 => "11101010",17414 => "10010111",17415 => "11111001",17416 => "10000100",17417 => "01010001",17418 => "00001101",17419 => "01100111",17420 => "01011111",17421 => "11011110",17422 => "00110111",17423 => "01010111",17424 => "01000001",17425 => "11100001",17426 => "00010110",17427 => "10110110",17428 => "10011111",17429 => "01111100",17430 => "00110001",17431 => "11001011",17432 => "10101110",17433 => "11110000",17434 => "01001111",17435 => "11010100",17436 => "01000100",17437 => "11001111",17438 => "10001010",17439 => "11010010",17440 => "00111010",17441 => "11011011",17442 => "01001100",17443 => "00100100",17444 => "00110011",17445 => "00011011",17446 => "01110011",17447 => "01011001",17448 => "01011101",17449 => "10110110",17450 => "00011000",17451 => "10111000",17452 => "11001111",17453 => "10101100",17454 => "11110011",17455 => "01001101",17456 => "11011111",17457 => "00010100",17458 => "11000011",17459 => "01110101",17460 => "01110000",17461 => "00000110",17462 => "01101010",17463 => "11111000",17464 => "11101111",17465 => "11111010",17466 => "00000100",17467 => "01111000",17468 => "01101100",17469 => "00010111",17470 => "10101000",17471 => "10100111",17472 => "11111000",17473 => "00000100",17474 => "10111100",17475 => "01101011",17476 => "01110101",17477 => "00111001",17478 => "11100111",17479 => "11011011",17480 => "00010011",17481 => "10100101",17482 => "01111011",17483 => "00000111",17484 => "01110100",17485 => "01110011",17486 => "01101111",17487 => "10000101",17488 => "00011000",17489 => "11100100",17490 => "00010001",17491 => "11110001",17492 => "10010011",17493 => "01101101",17494 => "01011011",17495 => "11100000",17496 => "11010100",17497 => "11111000",17498 => "01101100",17499 => "11001000",17500 => "01010111",17501 => "11101010",17502 => "00001001",17503 => "11000000",17504 => "10011111",17505 => "01011010",17506 => "10100011",17507 => "00101101",17508 => "01101001",17509 => "10100001",17510 => "11010011",17511 => "00001100",17512 => "11110101",17513 => "01111010",17514 => "11010000",17515 => "11100000",17516 => "00010101",17517 => "01101010",17518 => "00100000",17519 => "11111011",17520 => "01110100",17521 => "11110101",17522 => "11010000",17523 => "11110111",17524 => "00000111",17525 => "00100010",17526 => "10101101",17527 => "10110111",17528 => "10111111",17529 => "10001010",17530 => "00100101",17531 => "10101110",17532 => "00001110",17533 => "00110010",17534 => "00000100",17535 => "00101011",17536 => "10110101",17537 => "10101110",17538 => "01101100",17539 => "11000011",17540 => "10011111",17541 => "11000000",17542 => "10001011",17543 => "10110010",17544 => "00000111",17545 => "11010000",17546 => "00111000",17547 => "10101011",17548 => "10100011",17549 => "11000001",17550 => "00111100",17551 => "01000011",17552 => "01101010",17553 => "11001111",17554 => "00101011",17555 => "01000000",17556 => "11111010",17557 => "00010010",17558 => "01101111",17559 => "00101000",17560 => "01001111",17561 => "10000111",17562 => "10110010",17563 => "00010001",17564 => "10111011",17565 => "00000011",17566 => "10000110",17567 => "11111001",17568 => "00010100",17569 => "01001100",17570 => "10000110",17571 => "01111100",17572 => "10111011",17573 => "11001010",17574 => "01101101",17575 => "01101110",17576 => "11011101",17577 => "11110111",17578 => "10110000",17579 => "00001001",17580 => "11011110",17581 => "11010010",17582 => "10000110",17583 => "01100001",17584 => "11001001",17585 => "11010110",17586 => "10001001",17587 => "00101001",17588 => "00111100",17589 => "11110100",17590 => "00000001",17591 => "00111011",17592 => "10000001",17593 => "01011001",17594 => "00111101",17595 => "10110001",17596 => "11101100",17597 => "11011110",17598 => "00001001",17599 => "00011100",17600 => "11111100",17601 => "00010111",17602 => "00010110",17603 => "01111010",17604 => "01010000",17605 => "11001100",17606 => "11101101",17607 => "11010011",17608 => "00011011",17609 => "11110000",17610 => "10011000",17611 => "01000101",17612 => "11100100",17613 => "01001010",17614 => "00100010",17615 => "01111000",17616 => "00011000",17617 => "11010101",17618 => "00001111",17619 => "10000010",17620 => "11111010",17621 => "01111110",17622 => "01111110",17623 => "00000101",17624 => "00101111",17625 => "01110000",17626 => "01110101",17627 => "11101100",17628 => "11011011",17629 => "10101111",17630 => "01110011",17631 => "11011100",17632 => "10000100",17633 => "11010000",17634 => "10111010",17635 => "11100011",17636 => "00100001",17637 => "10100101",17638 => "11110101",17639 => "01111101",17640 => "11100101",17641 => "00100001",17642 => "00001101",17643 => "00111011",17644 => "11101010",17645 => "10100101",17646 => "00100000",17647 => "00111100",17648 => "10001000",17649 => "01100010",17650 => "11000111",17651 => "00010100",17652 => "11110001",17653 => "10001001",17654 => "01000011",17655 => "10111011",17656 => "01010110",17657 => "01111011",17658 => "01000000",17659 => "11011110",17660 => "01000110",17661 => "01100001",17662 => "01100111",17663 => "00101111",17664 => "01110000",17665 => "11001011",17666 => "10010111",17667 => "10001011",17668 => "00001101",17669 => "00001001",17670 => "11010011",17671 => "00011110",17672 => "10011001",17673 => "10010111",17674 => "10001000",17675 => "00101110",17676 => "01100101",17677 => "10101011",17678 => "11010100",17679 => "00110100",17680 => "00011111",17681 => "00111100",17682 => "11000101",17683 => "10000010",17684 => "00011010",17685 => "01010010",17686 => "11111101",17687 => "11101101",17688 => "01010101",17689 => "01011010",17690 => "10010000",17691 => "01000000",17692 => "11010101",17693 => "11001001",17694 => "01111011",17695 => "11011000",17696 => "11101001",17697 => "10110101",17698 => "10110110",17699 => "11000001",17700 => "11001000",17701 => "00100101",17702 => "10110011",17703 => "00000100",17704 => "01110010",17705 => "00011101",17706 => "01111101",17707 => "11001100",17708 => "01001010",17709 => "11111011",17710 => "11011101",17711 => "00111101",17712 => "10010101",17713 => "00011110",17714 => "01110011",17715 => "01000100",17716 => "01000011",17717 => "01000111",17718 => "01111101",17719 => "01111101",17720 => "01000101",17721 => "00110011",17722 => "00101000",17723 => "10010110",17724 => "10101101",17725 => "11000100",17726 => "00110110",17727 => "01001011",17728 => "01111100",17729 => "10100011",17730 => "10100101",17731 => "01001100",17732 => "00101100",17733 => "10001000",17734 => "00001100",17735 => "00001100",17736 => "10101101",17737 => "01100111",17738 => "11010101",17739 => "10101100",17740 => "00001010",17741 => "01011110",17742 => "00100011",17743 => "10010011",17744 => "01010010",17745 => "11000111",17746 => "10111000",17747 => "00110000",17748 => "00001110",17749 => "01110010",17750 => "00111100",17751 => "11111001",17752 => "00110111",17753 => "11110010",17754 => "01001011",17755 => "00011100",17756 => "00000010",17757 => "00111111",17758 => "01110110",17759 => "01011011",17760 => "10101110",17761 => "10110111",17762 => "00010100",17763 => "10001010",17764 => "11011000",17765 => "01010101",17766 => "00011001",17767 => "01010101",17768 => "01011010",17769 => "11001111",17770 => "00011000",17771 => "01111101",17772 => "00101010",17773 => "11100010",17774 => "11111101",17775 => "11111101",17776 => "10010101",17777 => "01011011",17778 => "00010000",17779 => "11010000",17780 => "10011010",17781 => "00110001",17782 => "10001100",17783 => "11001010",17784 => "01001110",17785 => "01110101",17786 => "00010111",17787 => "10100100",17788 => "10000000",17789 => "00100100",17790 => "01011011",17791 => "10110110",17792 => "00101111",17793 => "11101110",17794 => "00101110",17795 => "01100100",17796 => "10110010",17797 => "10000000",17798 => "00011000",17799 => "00101011",17800 => "00010100",17801 => "10010111",17802 => "11001000",17803 => "10011001",17804 => "10111111",17805 => "10000100",17806 => "00110100",17807 => "01000100",17808 => "00100111",17809 => "10000000",17810 => "10001011",17811 => "10111110",17812 => "10011010",17813 => "01100010",17814 => "00110011",17815 => "01110101",17816 => "00000000",17817 => "10011011",17818 => "11011010",17819 => "11011111",17820 => "00011011",17821 => "00011111",17822 => "01111110",17823 => "01101000",17824 => "00111100",17825 => "01001100",17826 => "00011011",17827 => "11110101",17828 => "01110010",17829 => "00010110",17830 => "00111010",17831 => "00011110",17832 => "11100011",17833 => "11110011",17834 => "01001110",17835 => "01000110",17836 => "11010100",17837 => "00000000",17838 => "10010110",17839 => "01100101",17840 => "00000011",17841 => "01111111",17842 => "11110100",17843 => "11101111",17844 => "10000000",17845 => "00100000",17846 => "01101000",17847 => "01100101",17848 => "10110100",17849 => "01100110",17850 => "11001101",17851 => "11010101",17852 => "10101100",17853 => "01011000",17854 => "10100000",17855 => "00100101",17856 => "11100110",17857 => "10111101",17858 => "10000110",17859 => "01101101",17860 => "11010110",17861 => "11111111",17862 => "00101110",17863 => "11100110",17864 => "00011100",17865 => "10010000",17866 => "00001000",17867 => "00010000",17868 => "00000111",17869 => "10110101",17870 => "10010110",17871 => "00010110",17872 => "11011101",17873 => "11110101",17874 => "00000110",17875 => "10111111",17876 => "11010010",17877 => "10011110",17878 => "11011001",17879 => "11011001",17880 => "11100000",17881 => "10011001",17882 => "10011010",17883 => "01100111",17884 => "00110000",17885 => "01100110",17886 => "01110110",17887 => "00110001",17888 => "01100011",17889 => "10001110",17890 => "10100010",17891 => "10011010",17892 => "10110101",17893 => "01111100",17894 => "10011111",17895 => "11000010",17896 => "00100101",17897 => "11010001",17898 => "01000111",17899 => "00101101",17900 => "10110110",17901 => "11011010",17902 => "01101110",17903 => "01100001",17904 => "00011011",17905 => "11101111",17906 => "11001111",17907 => "10111011",17908 => "10111010",17909 => "01111010",17910 => "10011000",17911 => "11110101",17912 => "10110011",17913 => "10111011",17914 => "11110110",17915 => "10100101",17916 => "11100100",17917 => "01001111",17918 => "00010001",17919 => "11110000",17920 => "10011100",17921 => "10000111",17922 => "00011111",17923 => "00010010",17924 => "00010011",17925 => "10010101",17926 => "11011011",17927 => "00001001",17928 => "11110110",17929 => "11111000",17930 => "01010011",17931 => "01011101",17932 => "01101010",17933 => "11011010",17934 => "11001110",17935 => "11101111",17936 => "10111110",17937 => "01110111",17938 => "01101001",17939 => "11010011",17940 => "10011101",17941 => "10111110",17942 => "10011110",17943 => "00101010",17944 => "01111110",17945 => "01010011",17946 => "01001011",17947 => "10011100",17948 => "10110000",17949 => "00000010",17950 => "01010101",17951 => "11010110",17952 => "01100110",17953 => "11010011",17954 => "01010001",17955 => "00100011",17956 => "10111110",17957 => "11001001",17958 => "11010101",17959 => "01110010",17960 => "01111111",17961 => "00011000",17962 => "01011001",17963 => "00110011",17964 => "01100101",17965 => "11001000",17966 => "01111101",17967 => "10010010",17968 => "10010000",17969 => "00101001",17970 => "10010011",17971 => "00110110",17972 => "01011000",17973 => "00110111",17974 => "11011011",17975 => "10110001",17976 => "01110010",17977 => "00000100",17978 => "01000111",17979 => "00001101",17980 => "10110011",17981 => "00110010",17982 => "00110110",17983 => "00001011",17984 => "10000000",17985 => "00010001",17986 => "10111010",17987 => "01111000",17988 => "01111000",17989 => "01110001",17990 => "00000001",17991 => "10101001",17992 => "01011111",17993 => "11011100",17994 => "01111000",17995 => "00000111",17996 => "00010000",17997 => "01000111",17998 => "00100101",17999 => "01100100",18000 => "10000011",18001 => "10111001",18002 => "11010100",18003 => "10010011",18004 => "11111110",18005 => "11011110",18006 => "11110010",18007 => "00101100",18008 => "10110111",18009 => "10100110",18010 => "10011001",18011 => "10001101",18012 => "00011101",18013 => "00000101",18014 => "11110110",18015 => "01001101",18016 => "01110000",18017 => "00001100",18018 => "11101100",18019 => "01110010",18020 => "01011110",18021 => "10010000",18022 => "11101001",18023 => "10111000",18024 => "01010100",18025 => "00110101",18026 => "01001111",18027 => "01101110",18028 => "10000001",18029 => "01101010",18030 => "10000001",18031 => "11011010",18032 => "10101100",18033 => "10110001",18034 => "01111111",18035 => "01100101",18036 => "01100011",18037 => "11111011",18038 => "00110011",18039 => "11101110",18040 => "00000101",18041 => "11000001",18042 => "01101001",18043 => "10111000",18044 => "10101101",18045 => "11110111",18046 => "10100011",18047 => "01101100",18048 => "10010001",18049 => "00011111",18050 => "00101101",18051 => "01101011",18052 => "00001010",18053 => "00110011",18054 => "10100100",18055 => "11111011",18056 => "10000100",18057 => "10101010",18058 => "01000000",18059 => "00110101",18060 => "01000011",18061 => "01111010",18062 => "01110001",18063 => "10101010",18064 => "00100100",18065 => "00111011",18066 => "11001110",18067 => "11111110",18068 => "11101110",18069 => "11010101",18070 => "00011001",18071 => "00001011",18072 => "00110101",18073 => "01110110",18074 => "01011010",18075 => "11100011",18076 => "00001110",18077 => "00011000",18078 => "10010001",18079 => "00101000",18080 => "00011101",18081 => "11000001",18082 => "01001110",18083 => "10110010",18084 => "10111100",18085 => "11010000",18086 => "00011111",18087 => "11000100",18088 => "01001000",18089 => "00010111",18090 => "10010110",18091 => "10000100",18092 => "00000000",18093 => "01001001",18094 => "01101101",18095 => "11000011",18096 => "11001010",18097 => "11111000",18098 => "11101110",18099 => "10111001",18100 => "11001000",18101 => "10000011",18102 => "01011011",18103 => "10000101",18104 => "10000010",18105 => "11010110",18106 => "11100010",18107 => "11001110",18108 => "01111001",18109 => "10011111",18110 => "00100110",18111 => "00111010",18112 => "11000000",18113 => "00001111",18114 => "01111010",18115 => "00011010",18116 => "11001011",18117 => "01001000",18118 => "10000001",18119 => "01110001",18120 => "00011100",18121 => "01110011",18122 => "11110110",18123 => "00100100",18124 => "10111101",18125 => "01010111",18126 => "01010001",18127 => "10111100",18128 => "01111011",18129 => "01110001",18130 => "11011110",18131 => "01110001",18132 => "00111101",18133 => "10111100",18134 => "00100100",18135 => "10001011",18136 => "00000100",18137 => "11101100",18138 => "10100101",18139 => "11011000",18140 => "11111101",18141 => "00010010",18142 => "00101111",18143 => "01111101",18144 => "00011100",18145 => "11011010",18146 => "01111110",18147 => "01001111",18148 => "10011111",18149 => "11010110",18150 => "01010000",18151 => "11001000",18152 => "11000010",18153 => "11001111",18154 => "11101000",18155 => "11110011",18156 => "11011001",18157 => "11010110",18158 => "11100001",18159 => "11100110",18160 => "00110010",18161 => "00011001",18162 => "01000000",18163 => "11011101",18164 => "00011010",18165 => "11001011",18166 => "00100100",18167 => "11010111",18168 => "11111010",18169 => "11100011",18170 => "11001110",18171 => "00110111",18172 => "00101010",18173 => "10010111",18174 => "11001101",18175 => "11110010",18176 => "11000101",18177 => "00001101",18178 => "01110101",18179 => "01111010",18180 => "00110110",18181 => "10011001",18182 => "11000010",18183 => "11100111",18184 => "11011001",18185 => "10110001",18186 => "10101110",18187 => "00000001",18188 => "01101011",18189 => "11010001",18190 => "11010011",18191 => "00000011",18192 => "00011100",18193 => "00110010",18194 => "00101110",18195 => "00000110",18196 => "11101001",18197 => "10001001",18198 => "01100100",18199 => "01111001",18200 => "00111111",18201 => "01000101",18202 => "11110100",18203 => "11111000",18204 => "01110001",18205 => "01101110",18206 => "01011101",18207 => "01001101",18208 => "10000000",18209 => "00011100",18210 => "11001100",18211 => "00110001",18212 => "01110011",18213 => "00011010",18214 => "10001001",18215 => "01011001",18216 => "11101110",18217 => "00000010",18218 => "00011100",18219 => "01010001",18220 => "11000110",18221 => "11001111",18222 => "00100010",18223 => "01001011",18224 => "00011001",18225 => "11111110",18226 => "10110000",18227 => "11100100",18228 => "10000010",18229 => "00100100",18230 => "10101011",18231 => "10010000",18232 => "01100100",18233 => "10110001",18234 => "00101010",18235 => "01010100",18236 => "11100110",18237 => "11110111",18238 => "01010110",18239 => "10111011",18240 => "01101000",18241 => "10010100",18242 => "11100001",18243 => "11100010",18244 => "01000110",18245 => "11110010",18246 => "11011001",18247 => "10101000",18248 => "11110110",18249 => "11110010",18250 => "10000101",18251 => "00010001",18252 => "11110110",18253 => "10100010",18254 => "10010011",18255 => "01111011",18256 => "11110010",18257 => "00101010",18258 => "10001100",18259 => "00100101",18260 => "10100100",18261 => "01000100",18262 => "00010001",18263 => "10010100",18264 => "00100001",18265 => "11110111",18266 => "00010010",18267 => "11111010",18268 => "01001010",18269 => "01110000",18270 => "11101101",18271 => "10111111",18272 => "11100000",18273 => "00001100",18274 => "01001011",18275 => "00010000",18276 => "01100011",18277 => "01111010",18278 => "10011010",18279 => "00001111",18280 => "10111001",18281 => "00011110",18282 => "00100001",18283 => "10111110",18284 => "10110000",18285 => "01011111",18286 => "00011011",18287 => "11010100",18288 => "01011110",18289 => "11100110",18290 => "01110110",18291 => "10000111",18292 => "10010001",18293 => "11001000",18294 => "11100001",18295 => "11011001",18296 => "11010100",18297 => "01101100",18298 => "10101110",18299 => "00111011",18300 => "01001100",18301 => "10101000",18302 => "11011100",18303 => "10111101",18304 => "01110010",18305 => "00000011",18306 => "11101000",18307 => "10111101",18308 => "00010000",18309 => "01100011",18310 => "01010111",18311 => "10000000",18312 => "11001000",18313 => "00111011",18314 => "10011111",18315 => "11101101",18316 => "00110101",18317 => "11001011",18318 => "11011101",18319 => "11100110",18320 => "01111100",18321 => "11010100",18322 => "11000011",18323 => "01111001",18324 => "00011101",18325 => "01101100",18326 => "00011000",18327 => "00101001",18328 => "00100101",18329 => "00111001",18330 => "00101001",18331 => "11001111",18332 => "01101111",18333 => "00000111",18334 => "01000001",18335 => "11110011",18336 => "01001110",18337 => "01000101",18338 => "11001100",18339 => "00111001",18340 => "10001000",18341 => "10000010",18342 => "01011000",18343 => "00010001",18344 => "00001010",18345 => "10010110",18346 => "00011101",18347 => "00101100",18348 => "01000001",18349 => "01101011",18350 => "01000001",18351 => "10111000",18352 => "01101010",18353 => "00000011",18354 => "11010000",18355 => "01111001",18356 => "01011010",18357 => "11010010",18358 => "01010010",18359 => "00011110",18360 => "10111000",18361 => "11011110",18362 => "10000101",18363 => "00110101",18364 => "10100100",18365 => "11000101",18366 => "00011010",18367 => "10000110",18368 => "01000111",18369 => "10011000",18370 => "00001110",18371 => "10100000",18372 => "10101010",18373 => "00111000",18374 => "00010011",18375 => "01010111",18376 => "10010010",18377 => "10100111",18378 => "00111010",18379 => "11100101",18380 => "00011101",18381 => "11111001",18382 => "01111111",18383 => "10100111",18384 => "10010000",18385 => "10110110",18386 => "11101111",18387 => "10011100",18388 => "11100010",18389 => "00101010",18390 => "00010111",18391 => "11100111",18392 => "01101111",18393 => "01001111",18394 => "00011001",18395 => "10001000",18396 => "11110110",18397 => "00111110",18398 => "01111110",18399 => "11101000",18400 => "10000001",18401 => "10000000",18402 => "01000010",18403 => "10111110",18404 => "11101010",18405 => "01101101",18406 => "00111000",18407 => "11000110",18408 => "01010101",18409 => "01010000",18410 => "01100010",18411 => "11010001",18412 => "10111111",18413 => "00100100",18414 => "01110100",18415 => "01000111",18416 => "10101100",18417 => "01110100",18418 => "01011100",18419 => "01101001",18420 => "10111101",18421 => "10000010",18422 => "11111101",18423 => "11111000",18424 => "01111111",18425 => "00100110",18426 => "11101111",18427 => "10010110",18428 => "10011000",18429 => "10001000",18430 => "10001111",18431 => "10111111",18432 => "01000100",18433 => "10111010",18434 => "00001100",18435 => "01010101",18436 => "10000001",18437 => "01011000",18438 => "11101111",18439 => "11001010",18440 => "00100010",18441 => "00001010",18442 => "00001100",18443 => "11100010",18444 => "11011011",18445 => "01110000",18446 => "11110011",18447 => "10101001",18448 => "01010110",18449 => "10000011",18450 => "00100100",18451 => "01111111",18452 => "10011110",18453 => "11001101",18454 => "10010001",18455 => "10010000",18456 => "01100110",18457 => "00000110",18458 => "01101110",18459 => "00100000",18460 => "01101001",18461 => "10011000",18462 => "00111100",18463 => "10111000",18464 => "00011000",18465 => "10101101",18466 => "11100101",18467 => "10111110",18468 => "00011011",18469 => "00110111",18470 => "11110111",18471 => "00100001",18472 => "00110111",18473 => "10111011",18474 => "01011000",18475 => "01110001",18476 => "11100001",18477 => "01001000",18478 => "01001101",18479 => "11001100",18480 => "11000011",18481 => "01011110",18482 => "01010101",18483 => "01000000",18484 => "11010110",18485 => "11110101",18486 => "00001101",18487 => "00101000",18488 => "01001100",18489 => "11010110",18490 => "01101001",18491 => "10011101",18492 => "01010100",18493 => "00101101",18494 => "10100100",18495 => "10001110",18496 => "00000000",18497 => "01111011",18498 => "10011011",18499 => "10100010",18500 => "11000111",18501 => "11011101",18502 => "00100011",18503 => "10010100",18504 => "00101101",18505 => "10011010",18506 => "10000110",18507 => "01111011",18508 => "10110111",18509 => "11000000",18510 => "00000000",18511 => "11010110",18512 => "00111110",18513 => "00010111",18514 => "10100001",18515 => "11001100",18516 => "01110011",18517 => "11000000",18518 => "01000010",18519 => "01100001",18520 => "11011010",18521 => "11111001",18522 => "10000110",18523 => "01110111",18524 => "00110001",18525 => "01111001",18526 => "01110111",18527 => "01010111",18528 => "11011100",18529 => "10110011",18530 => "11110011",18531 => "10001111",18532 => "00110111",18533 => "00100000",18534 => "00111100",18535 => "10011101",18536 => "10001000",18537 => "00101110",18538 => "10001000",18539 => "01100001",18540 => "10100001",18541 => "11100110",18542 => "01010000",18543 => "01110101",18544 => "00101111",18545 => "11111111",18546 => "10010101",18547 => "00000101",18548 => "10110111",18549 => "00100101",18550 => "11100001",18551 => "00101110",18552 => "00011010",18553 => "01101001",18554 => "10000010",18555 => "11010000",18556 => "10111000",18557 => "11101001",18558 => "11010110",18559 => "11100000",18560 => "10100100",18561 => "01101010",18562 => "00010110",18563 => "00110001",18564 => "10000001",18565 => "00000100",18566 => "01110101",18567 => "11111000",18568 => "10111111",18569 => "00011010",18570 => "01011000",18571 => "00101010",18572 => "00111100",18573 => "10111110",18574 => "00010000",18575 => "10010001",18576 => "10000001",18577 => "10101000",18578 => "11111101",18579 => "10000110",18580 => "00100111",18581 => "11101001",18582 => "11010100",18583 => "10100011",18584 => "01000000",18585 => "11100000",18586 => "10101100",18587 => "11110101",18588 => "10011101",18589 => "01001111",18590 => "11110001",18591 => "11001011",18592 => "01111111",18593 => "00011101",18594 => "01111001",18595 => "00111000",18596 => "10110010",18597 => "00010100",18598 => "00100111",18599 => "10000000",18600 => "10001110",18601 => "01000111",18602 => "11001111",18603 => "00101011",18604 => "10100101",18605 => "00110000",18606 => "00100100",18607 => "00111111",18608 => "11010100",18609 => "11000101",18610 => "00100101",18611 => "01011100",18612 => "10111010",18613 => "11011001",18614 => "00010110",18615 => "11001011",18616 => "11011110",18617 => "01111010",18618 => "10001001",18619 => "11001101",18620 => "10101011",18621 => "01000011",18622 => "10000010",18623 => "01001000",18624 => "11011100",18625 => "10001111",18626 => "01100111",18627 => "10111110",18628 => "00000011",18629 => "11100010",18630 => "10111100",18631 => "10001111",18632 => "00011100",18633 => "10110000",18634 => "11111011",18635 => "00111001",18636 => "01000001",18637 => "11010110",18638 => "00110101",18639 => "11011001",18640 => "00010001",18641 => "00111100",18642 => "11101001",18643 => "01001000",18644 => "10001111",18645 => "11100110",18646 => "10011010",18647 => "10001000",18648 => "01100110",18649 => "11111100",18650 => "10000111",18651 => "11011110",18652 => "11100001",18653 => "11001010",18654 => "10110100",18655 => "10011010",18656 => "10100101",18657 => "10010100",18658 => "00111000",18659 => "01111001",18660 => "10111000",18661 => "00111001",18662 => "11111010",18663 => "00111101",18664 => "11110010",18665 => "11000101",18666 => "01001110",18667 => "00110010",18668 => "11011000",18669 => "10111011",18670 => "11010001",18671 => "01011000",18672 => "00000101",18673 => "10111100",18674 => "11001001",18675 => "00001111",18676 => "10011001",18677 => "00111110",18678 => "10100001",18679 => "11010001",18680 => "11001110",18681 => "11101011",18682 => "01000110",18683 => "10101101",18684 => "10011111",18685 => "00000010",18686 => "01001100",18687 => "00000001",18688 => "01110000",18689 => "10010001",18690 => "10000110",18691 => "01000101",18692 => "00111001",18693 => "11010010",18694 => "10010101",18695 => "00110001",18696 => "10101010",18697 => "01100000",18698 => "01001110",18699 => "01010001",18700 => "11110110",18701 => "01010100",18702 => "11111111",18703 => "00010100",18704 => "01010011",18705 => "01111111",18706 => "01011100",18707 => "11100110",18708 => "10100000",18709 => "00100011",18710 => "11110011",18711 => "01111101",18712 => "10011111",18713 => "10011010",18714 => "00000001",18715 => "11110011",18716 => "00101110",18717 => "10100011",18718 => "01010010",18719 => "01011010",18720 => "00110101",18721 => "00100110",18722 => "01110101",18723 => "01101011",18724 => "10010100",18725 => "01001110",18726 => "11110100",18727 => "01011100",18728 => "00111100",18729 => "01001101",18730 => "01010010",18731 => "10000011",18732 => "00000111",18733 => "10110010",18734 => "01011001",18735 => "00001111",18736 => "11101110",18737 => "11110000",18738 => "11001001",18739 => "11100101",18740 => "11110101",18741 => "11000111",18742 => "01110011",18743 => "00110100",18744 => "10101010",18745 => "11100001",18746 => "10101011",18747 => "00111011",18748 => "10000100",18749 => "01110101",18750 => "01001111",18751 => "11011010",18752 => "00010100",18753 => "00000011",18754 => "01111001",18755 => "01010101",18756 => "10101111",18757 => "01010111",18758 => "00011101",18759 => "11000111",18760 => "00011000",18761 => "11100000",18762 => "01010000",18763 => "10111011",18764 => "10111000",18765 => "01110111",18766 => "10101100",18767 => "01101000",18768 => "11011000",18769 => "01010011",18770 => "11001001",18771 => "11110100",18772 => "01011000",18773 => "10011000",18774 => "01001101",18775 => "10101101",18776 => "11011000",18777 => "01110011",18778 => "11101111",18779 => "10011110",18780 => "10010110",18781 => "11101110",18782 => "10110011",18783 => "10000111",18784 => "10101000",18785 => "10101000",18786 => "00101111",18787 => "01010111",18788 => "11011101",18789 => "10010100",18790 => "00110110",18791 => "10100001",18792 => "00111100",18793 => "01110011",18794 => "01010000",18795 => "01011001",18796 => "10111000",18797 => "10100100",18798 => "00110111",18799 => "00010010",18800 => "01101000",18801 => "00001010",18802 => "01011101",18803 => "00101001",18804 => "01001101",18805 => "01001101",18806 => "00110111",18807 => "11101000",18808 => "10010001",18809 => "11001110",18810 => "11010111",18811 => "00001001",18812 => "11001101",18813 => "11111011",18814 => "00101010",18815 => "01010000",18816 => "01001001",18817 => "01000001",18818 => "00000100",18819 => "01111110",18820 => "11111011",18821 => "00010110",18822 => "00011010",18823 => "11100011",18824 => "11111111",18825 => "10101100",18826 => "11010001",18827 => "11111100",18828 => "00110001",18829 => "00111101",18830 => "01001101",18831 => "00011000",18832 => "01001101",18833 => "00110001",18834 => "00000000",18835 => "00001100",18836 => "11000011",18837 => "10011001",18838 => "10011011",18839 => "11101101",18840 => "01100011",18841 => "00111101",18842 => "10100101",18843 => "11111010",18844 => "11110100",18845 => "10111001",18846 => "10111100",18847 => "11000001",18848 => "10001101",18849 => "10001111",18850 => "01100011",18851 => "11111100",18852 => "11011001",18853 => "10111111",18854 => "01010100",18855 => "00010101",18856 => "10001010",18857 => "00011010",18858 => "10000111",18859 => "11111101",18860 => "10111111",18861 => "00111110",18862 => "10101000",18863 => "10110010",18864 => "10101100",18865 => "00010010",18866 => "01111100",18867 => "00001100",18868 => "11101101",18869 => "11001001",18870 => "00110100",18871 => "11010101",18872 => "11101001",18873 => "10001111",18874 => "10001000",18875 => "10111000",18876 => "10111010",18877 => "11100111",18878 => "11101110",18879 => "11101011",18880 => "10000011",18881 => "10100110",18882 => "00000011",18883 => "11110110",18884 => "10010001",18885 => "01111110",18886 => "00010001",18887 => "11111011",18888 => "10010111",18889 => "11010101",18890 => "01000011",18891 => "01000100",18892 => "10001000",18893 => "00111101",18894 => "00010001",18895 => "00100111",18896 => "00011110",18897 => "00110111",18898 => "00101101",18899 => "01000001",18900 => "01011100",18901 => "10111011",18902 => "00111101",18903 => "11110100",18904 => "01110011",18905 => "01110101",18906 => "10011001",18907 => "11010111",18908 => "00111110",18909 => "10110110",18910 => "01100101",18911 => "11110110",18912 => "10010100",18913 => "01111100",18914 => "11110011",18915 => "01001001",18916 => "10001100",18917 => "10011000",18918 => "11110000",18919 => "11011101",18920 => "10111001",18921 => "00011101",18922 => "11110110",18923 => "11010101",18924 => "10010100",18925 => "00001000",18926 => "11011011",18927 => "01111011",18928 => "11011011",18929 => "01101010",18930 => "10111001",18931 => "00100010",18932 => "11100001",18933 => "10010111",18934 => "11110011",18935 => "00011100",18936 => "10111001",18937 => "10111110",18938 => "01011100",18939 => "01101001",18940 => "00111100",18941 => "11111111",18942 => "01101110",18943 => "00110011",18944 => "01100000",18945 => "00001000",18946 => "00001111",18947 => "11101100",18948 => "01100100",18949 => "10010000",18950 => "10101110",18951 => "00010111",18952 => "10100101",18953 => "10100011",18954 => "10010101",18955 => "11010010",18956 => "00000010",18957 => "11111001",18958 => "11011100",18959 => "11000001",18960 => "01101101",18961 => "10110010",18962 => "00001001",18963 => "01001011",18964 => "01111101",18965 => "10010100",18966 => "10111001",18967 => "10110010",18968 => "11001010",18969 => "01011000",18970 => "11011000",18971 => "01110001",18972 => "01101011",18973 => "10111000",18974 => "10101100",18975 => "11100101",18976 => "00000110",18977 => "00000010",18978 => "00110000",18979 => "01000111",18980 => "00000111",18981 => "01011100",18982 => "00111111",18983 => "00101111",18984 => "10000110",18985 => "10000011",18986 => "11111110",18987 => "10000110",18988 => "10010001",18989 => "11101011",18990 => "11110100",18991 => "11100101",18992 => "00110000",18993 => "01000111",18994 => "00110100",18995 => "10100110",18996 => "10000111",18997 => "01100010",18998 => "10111110",18999 => "01100101",19000 => "01001000",19001 => "10110010",19002 => "10010001",19003 => "01100011",19004 => "11110011",19005 => "11101001",19006 => "10110011",19007 => "01001101",19008 => "01000100",19009 => "00111011",19010 => "01101110",19011 => "01100011",19012 => "00100110",19013 => "01011001",19014 => "01111001",19015 => "01001000",19016 => "00001011",19017 => "11011100",19018 => "11101110",19019 => "11101101",19020 => "00011010",19021 => "11111000",19022 => "01101010",19023 => "10111000",19024 => "10011001",19025 => "11110000",19026 => "10100110",19027 => "11111110",19028 => "01101101",19029 => "10000000",19030 => "11010101",19031 => "11111010",19032 => "00010000",19033 => "11100001",19034 => "01100010",19035 => "01001011",19036 => "11101110",19037 => "11011111",19038 => "00011110",19039 => "01001110",19040 => "01011101",19041 => "01100100",19042 => "00000000",19043 => "00001000",19044 => "01101111",19045 => "01001100",19046 => "01000111",19047 => "00111000",19048 => "10011010",19049 => "00001001",19050 => "00100011",19051 => "00001001",19052 => "10010001",19053 => "00100100",19054 => "01100011",19055 => "10001001",19056 => "00110010",19057 => "11110010",19058 => "00010110",19059 => "00100010",19060 => "10011001",19061 => "00111000",19062 => "00110001",19063 => "11110010",19064 => "01111001",19065 => "11111100",19066 => "10011100",19067 => "00110001",19068 => "01001011",19069 => "01011110",19070 => "01011110",19071 => "00001110",19072 => "00011010",19073 => "11110101",19074 => "01001011",19075 => "10001100",19076 => "10010100",19077 => "00010011",19078 => "00110111",19079 => "11111011",19080 => "10011110",19081 => "10100011",19082 => "10011011",19083 => "10000011",19084 => "10010011",19085 => "00000010",19086 => "00000000",19087 => "01010000",19088 => "01110011",19089 => "00011101",19090 => "01011100",19091 => "10000011",19092 => "01011110",19093 => "10011100",19094 => "01101101",19095 => "01111001",19096 => "10101011",19097 => "00101110",19098 => "00011001",19099 => "11000110",19100 => "01111110",19101 => "10001110",19102 => "10011001",19103 => "01101111",19104 => "01011100",19105 => "10000110",19106 => "10010000",19107 => "10000111",19108 => "11111011",19109 => "00110110",19110 => "01011111",19111 => "01111011",19112 => "10100011",19113 => "10100001",19114 => "01100110",19115 => "00000110",19116 => "10000100",19117 => "11000100",19118 => "00010001",19119 => "10011010",19120 => "00010101",19121 => "00001010",19122 => "10101000",19123 => "01111110",19124 => "01100101",19125 => "00011100",19126 => "10110011",19127 => "11011001",19128 => "11111010",19129 => "00000111",19130 => "11000010",19131 => "11110010",19132 => "00100111",19133 => "01011010",19134 => "10111100",19135 => "01000001",19136 => "11110000",19137 => "01011000",19138 => "00001110",19139 => "11000110",19140 => "00111011",19141 => "10001111",19142 => "10000111",19143 => "01001101",19144 => "10111101",19145 => "01110011",19146 => "00000101",19147 => "01101100",19148 => "00101101",19149 => "00111000",19150 => "01100000",19151 => "11010000",19152 => "01101101",19153 => "11101000",19154 => "11101101",19155 => "00110011",19156 => "11011100",19157 => "10001101",19158 => "10010100",19159 => "01001110",19160 => "11111000",19161 => "01000111",19162 => "10101010",19163 => "00111111",19164 => "11000100",19165 => "00011001",19166 => "00001011",19167 => "01111100",19168 => "01011000",19169 => "01100000",19170 => "00100010",19171 => "11000011",19172 => "00100111",19173 => "01001000",19174 => "11011100",19175 => "00010011",19176 => "11011000",19177 => "00001000",19178 => "11100111",19179 => "00011100",19180 => "10001011",19181 => "00101100",19182 => "00010110",19183 => "01100110",19184 => "00100110",19185 => "11111000",19186 => "11010101",19187 => "10101011",19188 => "11111111",19189 => "11110111",19190 => "10100111",19191 => "01010000",19192 => "01111100",19193 => "11111001",19194 => "00110000",19195 => "10111101",19196 => "10110100",19197 => "10011110",19198 => "10001111",19199 => "11110001",19200 => "00010010",19201 => "00101001",19202 => "10010010",19203 => "01010010",19204 => "00001000",19205 => "00001001",19206 => "00001111",19207 => "01110000",19208 => "01000101",19209 => "01000001",19210 => "00111110",19211 => "01011001",19212 => "01001011",19213 => "01000000",19214 => "11110001",19215 => "10100110",19216 => "00101111",19217 => "01000100",19218 => "00011110",19219 => "10010010",19220 => "11001011",19221 => "10111011",19222 => "10111001",19223 => "00100000",19224 => "10000011",19225 => "00101100",19226 => "01111010",19227 => "01011111",19228 => "11101100",19229 => "11000011",19230 => "10110101",19231 => "10011101",19232 => "01011000",19233 => "00111100",19234 => "10000110",19235 => "01101110",19236 => "11001001",19237 => "11001100",19238 => "11000101",19239 => "00101000",19240 => "00110101",19241 => "11011111",19242 => "10100111",19243 => "11001101",19244 => "00010101",19245 => "11110101",19246 => "01101110",19247 => "01000101",19248 => "11100100",19249 => "00011011",19250 => "11010000",19251 => "11000001",19252 => "00100000",19253 => "11111110",19254 => "01100010",19255 => "10000010",19256 => "01000010",19257 => "00101100",19258 => "11101011",19259 => "01000111",19260 => "11101101",19261 => "01001100",19262 => "01101101",19263 => "10000111",19264 => "00111110",19265 => "00101111",19266 => "00011010",19267 => "10000000",19268 => "10100110",19269 => "11001011",19270 => "10111010",19271 => "00000110",19272 => "11100001",19273 => "00001100",19274 => "00111000",19275 => "01000111",19276 => "10100010",19277 => "01011101",19278 => "00111111",19279 => "00000010",19280 => "11110010",19281 => "11001100",19282 => "01011011",19283 => "00000101",19284 => "11010100",19285 => "00010001",19286 => "01100011",19287 => "10101000",19288 => "01001110",19289 => "11111011",19290 => "11100100",19291 => "01100011",19292 => "10110101",19293 => "10100010",19294 => "11001001",19295 => "01011100",19296 => "10010011",19297 => "11000000",19298 => "01010100",19299 => "01000111",19300 => "11101100",19301 => "10000101",19302 => "11111111",19303 => "01101101",19304 => "11010110",19305 => "00011110",19306 => "11110110",19307 => "00000000",19308 => "01101000",19309 => "01011010",19310 => "10100011",19311 => "00010011",19312 => "11001011",19313 => "00001001",19314 => "10100010",19315 => "01011000",19316 => "10001010",19317 => "01111000",19318 => "11000011",19319 => "10110001",19320 => "10110100",19321 => "10111100",19322 => "00101111",19323 => "01100000",19324 => "01000001",19325 => "11001001",19326 => "10010100",19327 => "01111111",19328 => "01011001",19329 => "10100111",19330 => "10010111",19331 => "11100100",19332 => "01110110",19333 => "00011010",19334 => "00010001",19335 => "00110110",19336 => "11011011",19337 => "10000001",19338 => "11010010",19339 => "10101000",19340 => "01111100",19341 => "10000101",19342 => "10110011",19343 => "11100000",19344 => "11110100",19345 => "01110000",19346 => "01000001",19347 => "11111111",19348 => "11010101",19349 => "10101011",19350 => "10001011",19351 => "11101110",19352 => "01001011",19353 => "10010000",19354 => "00010001",19355 => "10111101",19356 => "00110100",19357 => "10011111",19358 => "10100010",19359 => "00000001",19360 => "01101111",19361 => "00001001",19362 => "10000001",19363 => "10111000",19364 => "10010011",19365 => "11001111",19366 => "01101000",19367 => "00110110",19368 => "10100101",19369 => "00010011",19370 => "11111000",19371 => "11110001",19372 => "11001111",19373 => "01100000",19374 => "11111011",19375 => "01111100",19376 => "10001101",19377 => "10001000",19378 => "00100001",19379 => "10010111",19380 => "11100110",19381 => "10010010",19382 => "00111101",19383 => "10000101",19384 => "00011010",19385 => "00010100",19386 => "10110010",19387 => "10001001",19388 => "11111011",19389 => "11001101",19390 => "01100100",19391 => "11001101",19392 => "10100111",19393 => "11100001",19394 => "01011101",19395 => "11000110",19396 => "10110001",19397 => "11011010",19398 => "10101001",19399 => "11001100",19400 => "00011010",19401 => "11101110",19402 => "01000010",19403 => "11111000",19404 => "11100000",19405 => "00010101",19406 => "01111010",19407 => "01010111",19408 => "10001100",19409 => "11010000",19410 => "00001110",19411 => "10001001",19412 => "00111010",19413 => "11011000",19414 => "01000011",19415 => "01101011",19416 => "00000100",19417 => "00011010",19418 => "10011001",19419 => "11100111",19420 => "11111110",19421 => "00101111",19422 => "10111110",19423 => "00010101",19424 => "00101110",19425 => "11001001",19426 => "00000000",19427 => "10000100",19428 => "11111101",19429 => "00001000",19430 => "11001110",19431 => "00001101",19432 => "01111110",19433 => "00001101",19434 => "10001000",19435 => "01011010",19436 => "01100100",19437 => "01111000",19438 => "10000010",19439 => "00000001",19440 => "11010110",19441 => "11100111",19442 => "10001100",19443 => "11101011",19444 => "01001100",19445 => "11101100",19446 => "11111101",19447 => "00100011",19448 => "01111101",19449 => "10010001",19450 => "11111011",19451 => "10101000",19452 => "00001110",19453 => "01110100",19454 => "01111000",19455 => "00001110",19456 => "11101100",19457 => "01010011",19458 => "00101111",19459 => "10001010",19460 => "11110110",19461 => "00011111",19462 => "01110010",19463 => "01110111",19464 => "11011111",19465 => "01101001",19466 => "00110001",19467 => "01100110",19468 => "01010100",19469 => "01011111",19470 => "10110110",19471 => "11011100",19472 => "00010111",19473 => "10010010",19474 => "10100010",19475 => "11101100",19476 => "11011111",19477 => "01101010",19478 => "10111110",19479 => "11110110",19480 => "11001011",19481 => "00000100",19482 => "10101001",19483 => "11111111",19484 => "00110111",19485 => "00011011",19486 => "01010111",19487 => "11000100",19488 => "01111110",19489 => "10011000",19490 => "01011100",19491 => "01101000",19492 => "10000000",19493 => "10001011",19494 => "01111011",19495 => "01111010",19496 => "01111000",19497 => "11100110",19498 => "01100001",19499 => "11101000",19500 => "00011000",19501 => "00111010",19502 => "11111010",19503 => "10100001",19504 => "10101100",19505 => "11010010",19506 => "01000110",19507 => "11101001",19508 => "00010010",19509 => "11011000",19510 => "01001100",19511 => "10111010",19512 => "01011010",19513 => "11010100",19514 => "11110100",19515 => "11100000",19516 => "11100010",19517 => "00110101",19518 => "11011011",19519 => "01100011",19520 => "11110010",19521 => "01011000",19522 => "01001111",19523 => "01001010",19524 => "11010010",19525 => "11010011",19526 => "11110110",19527 => "00011000",19528 => "10100100",19529 => "00001110",19530 => "01110001",19531 => "10100000",19532 => "00000001",19533 => "10000010",19534 => "10100101",19535 => "01111011",19536 => "10011100",19537 => "01011000",19538 => "00100111",19539 => "10100100",19540 => "11110100",19541 => "00101000",19542 => "10111101",19543 => "01110100",19544 => "10001011",19545 => "10110100",19546 => "00111011",19547 => "01011101",19548 => "11101011",19549 => "10000111",19550 => "00010000",19551 => "01110001",19552 => "11010001",19553 => "11011000",19554 => "11111000",19555 => "00101001",19556 => "01100000",19557 => "01100101",19558 => "11011110",19559 => "01000000",19560 => "01101001",19561 => "01011111",19562 => "11010101",19563 => "00001101",19564 => "00000110",19565 => "00111111",19566 => "00110000",19567 => "00000101",19568 => "01101100",19569 => "00100110",19570 => "10100111",19571 => "10101100",19572 => "10010010",19573 => "00001011",19574 => "10010011",19575 => "01110001",19576 => "11011101",19577 => "11110001",19578 => "00000011",19579 => "10101000",19580 => "01110001",19581 => "11111000",19582 => "00111011",19583 => "11101101",19584 => "00000000",19585 => "01010011",19586 => "11101011",19587 => "00101010",19588 => "10010110",19589 => "11100000",19590 => "10111000",19591 => "11000110",19592 => "00110010",19593 => "10000011",19594 => "01010100",19595 => "10001001",19596 => "01000100",19597 => "10000100",19598 => "10000010",19599 => "01001100",19600 => "01011110",19601 => "11111000",19602 => "01110011",19603 => "00010101",19604 => "00100110",19605 => "10001101",19606 => "11010101",19607 => "00001110",19608 => "11001110",19609 => "11101100",19610 => "11100011",19611 => "01001100",19612 => "10000001",19613 => "11000010",19614 => "10100000",19615 => "01001110",19616 => "01111101",19617 => "00011100",19618 => "10110000",19619 => "01000101",19620 => "11100101",19621 => "10101010",19622 => "01110111",19623 => "01101100",19624 => "00010110",19625 => "11010110",19626 => "10000011",19627 => "11110100",19628 => "11001011",19629 => "01011110",19630 => "10100101",19631 => "00010110",19632 => "10001001",19633 => "00110011",19634 => "10111111",19635 => "11101110",19636 => "00100000",19637 => "11010100",19638 => "01100111",19639 => "00110001",19640 => "11111100",19641 => "11110011",19642 => "01100111",19643 => "00110110",19644 => "00011110",19645 => "00111010",19646 => "10110111",19647 => "01001110",19648 => "10111100",19649 => "10100010",19650 => "10011001",19651 => "00001000",19652 => "11010111",19653 => "01111001",19654 => "11000011",19655 => "11000111",19656 => "00000110",19657 => "00100011",19658 => "11000001",19659 => "11000101",19660 => "11101110",19661 => "11101100",19662 => "00100010",19663 => "10000100",19664 => "11001010",19665 => "10010010",19666 => "01001001",19667 => "10110110",19668 => "11010100",19669 => "00110011",19670 => "00100001",19671 => "01001100",19672 => "00110100",19673 => "10001100",19674 => "01011100",19675 => "11000011",19676 => "11110011",19677 => "00101010",19678 => "10010011",19679 => "10111011",19680 => "10111101",19681 => "00111001",19682 => "11000111",19683 => "00010000",19684 => "00011110",19685 => "00000111",19686 => "00010100",19687 => "00100010",19688 => "10110011",19689 => "10001011",19690 => "00110010",19691 => "10000011",19692 => "01111001",19693 => "00101011",19694 => "00110011",19695 => "01011111",19696 => "01010101",19697 => "01101001",19698 => "00110110",19699 => "01101100",19700 => "01110100",19701 => "11001010",19702 => "10100001",19703 => "00100001",19704 => "01001101",19705 => "01010110",19706 => "10101111",19707 => "01110100",19708 => "00010001",19709 => "10111110",19710 => "10001101",19711 => "01001100",19712 => "00011111",19713 => "00010100",19714 => "11000010",19715 => "01101001",19716 => "01010101",19717 => "00000100",19718 => "11010001",19719 => "10000100",19720 => "11111110",19721 => "01111000",19722 => "10110010",19723 => "10001101",19724 => "11100100",19725 => "11101001",19726 => "11011110",19727 => "11101100",19728 => "11001010",19729 => "01010111",19730 => "10111110",19731 => "01000001",19732 => "01010010",19733 => "01000001",19734 => "10001100",19735 => "01001110",19736 => "00000101",19737 => "11000100",19738 => "00101010",19739 => "10010010",19740 => "11110100",19741 => "00101010",19742 => "10111111",19743 => "00010010",19744 => "11000101",19745 => "11110011",19746 => "10100111",19747 => "00111000",19748 => "11111101",19749 => "00100100",19750 => "00000000",19751 => "00000100",19752 => "01000111",19753 => "10110111",19754 => "10100101",19755 => "00111001",19756 => "11101110",19757 => "00000101",19758 => "11111100",19759 => "11001011",19760 => "00100100",19761 => "10101100",19762 => "11010100",19763 => "10111110",19764 => "00011110",19765 => "10101100",19766 => "11100110",19767 => "11001010",19768 => "00000100",19769 => "10101010",19770 => "01010010",19771 => "11001101",19772 => "11000101",19773 => "01111010",19774 => "11010011",19775 => "11101000",19776 => "00111000",19777 => "01001000",19778 => "00010101",19779 => "11110110",19780 => "11110010",19781 => "10100000",19782 => "11100110",19783 => "00110011",19784 => "00110001",19785 => "11111100",19786 => "00100001",19787 => "11000101",19788 => "10010010",19789 => "01111101",19790 => "11011000",19791 => "11010000",19792 => "11110001",19793 => "10000011",19794 => "11001001",19795 => "11110110",19796 => "10001101",19797 => "11110100",19798 => "00010010",19799 => "01001011",19800 => "11110101",19801 => "10101101",19802 => "01101110",19803 => "01001000",19804 => "01001101",19805 => "11010001",19806 => "00000001",19807 => "10000000",19808 => "00011111",19809 => "00110000",19810 => "01000011",19811 => "10001010",19812 => "01011110",19813 => "10100001",19814 => "01001100",19815 => "00010010",19816 => "10001111",19817 => "01101110",19818 => "10001001",19819 => "10110011",19820 => "10000000",19821 => "00100100",19822 => "10010100",19823 => "11001101",19824 => "00000111",19825 => "00011111",19826 => "10101001",19827 => "01101010",19828 => "00100000",19829 => "01001001",19830 => "01110001",19831 => "00000100",19832 => "01100011",19833 => "11110000",19834 => "00010011",19835 => "10110001",19836 => "11100100",19837 => "01100101",19838 => "00010010",19839 => "10011110",19840 => "11010101",19841 => "01110111",19842 => "10110110",19843 => "10100000",19844 => "01011111",19845 => "00100101",19846 => "01010101",19847 => "10100010",19848 => "01010011",19849 => "10011110",19850 => "11001001",19851 => "01110111",19852 => "11101110",19853 => "11010000",19854 => "11001000",19855 => "10111000",19856 => "11010001",19857 => "11101100",19858 => "10010111",19859 => "01000110",19860 => "01100101",19861 => "00100011",19862 => "10000100",19863 => "10010000",19864 => "11001111",19865 => "10100101",19866 => "11001100",19867 => "00001000",19868 => "01100101",19869 => "01101100",19870 => "01101110",19871 => "11000110",19872 => "01110000",19873 => "10001000",19874 => "11010001",19875 => "11100001",19876 => "00101110",19877 => "01111101",19878 => "01111100",19879 => "11010010",19880 => "01000111",19881 => "10000101",19882 => "00010011",19883 => "11101111",19884 => "00110110",19885 => "01010100",19886 => "00000010",19887 => "00101100",19888 => "10110001",19889 => "11110011",19890 => "10001111",19891 => "01010000",19892 => "00110010",19893 => "01001110",19894 => "01000001",19895 => "00101011",19896 => "10010000",19897 => "01110110",19898 => "11001010",19899 => "11111110",19900 => "01010100",19901 => "10110000",19902 => "11011100",19903 => "10101111",19904 => "11011010",19905 => "01001000",19906 => "00010011",19907 => "00010100",19908 => "10010110",19909 => "01000001",19910 => "01101100",19911 => "10000001",19912 => "10100101",19913 => "01010110",19914 => "00000100",19915 => "11010110",19916 => "00111010",19917 => "00011011",19918 => "00001011",19919 => "00011011",19920 => "10110100",19921 => "11100010",19922 => "11110011",19923 => "01110001",19924 => "00011010",19925 => "00000011",19926 => "11010001",19927 => "11011010",19928 => "00010001",19929 => "11100011",19930 => "00011011",19931 => "01010000",19932 => "11101001",19933 => "00000001",19934 => "10010000",19935 => "10011011",19936 => "11110000",19937 => "11110100",19938 => "11100000",19939 => "10010110",19940 => "11001111",19941 => "01011010",19942 => "01100001",19943 => "01100101",19944 => "10110011",19945 => "10010000",19946 => "00100001",19947 => "11010110",19948 => "00000001",19949 => "00110111",19950 => "10011000",19951 => "00001000",19952 => "11010100",19953 => "00001100",19954 => "00111010",19955 => "00100011",19956 => "11111011",19957 => "01011101",19958 => "01100001",19959 => "10100001",19960 => "01001000",19961 => "11010111",19962 => "11011011",19963 => "11101101",19964 => "11010111",19965 => "10111010",19966 => "01010010",19967 => "00111000",19968 => "01000000",19969 => "00111100",19970 => "10010110",19971 => "00011011",19972 => "00111100",19973 => "11101001",19974 => "11000011",19975 => "10111001",19976 => "00000100",19977 => "10010011",19978 => "10011001",19979 => "11001001",19980 => "11101010",19981 => "10000101",19982 => "01100011",19983 => "00100010",19984 => "11110111",19985 => "10111101",19986 => "01010111",19987 => "00000010",19988 => "11111000",19989 => "01100011",19990 => "01110000",19991 => "01111011",19992 => "01000001",19993 => "11001101",19994 => "01100100",19995 => "01011110",19996 => "10100100",19997 => "11101101",19998 => "11010101",19999 => "00010110",20000 => "11101001",20001 => "00000000",20002 => "01011000",20003 => "01010111",20004 => "00101001",20005 => "11000001",20006 => "01000001",20007 => "10101101",20008 => "10111111",20009 => "10000011",20010 => "10010100",20011 => "11000101",20012 => "10101010",20013 => "00000001",20014 => "01000001",20015 => "00000010",20016 => "11110110",20017 => "00101001",20018 => "10101011",20019 => "00111111",20020 => "00100001",20021 => "11001111",20022 => "11100001",20023 => "00011000",20024 => "10101000",20025 => "01110101",20026 => "11110000",20027 => "01011011",20028 => "10001000",20029 => "01011100",20030 => "10101010",20031 => "01010111",20032 => "11101001",20033 => "11000000",20034 => "11110110",20035 => "11100111",20036 => "01100100",20037 => "01100111",20038 => "11100000",20039 => "00110100",20040 => "10001011",20041 => "01101100",20042 => "11101111",20043 => "01010011",20044 => "01010101",20045 => "11011101",20046 => "10111001",20047 => "01001111",20048 => "00011011",20049 => "11011000",20050 => "11001101",20051 => "11000100",20052 => "11111110",20053 => "00011100",20054 => "00111100",20055 => "00011001",20056 => "10111011",20057 => "00101010",20058 => "01000111",20059 => "11010111",20060 => "00010010",20061 => "01111101",20062 => "11110101",20063 => "10101010",20064 => "01111000",20065 => "11011111",20066 => "00100111",20067 => "00010000",20068 => "11101000",20069 => "11101110",20070 => "01111011",20071 => "10000100",20072 => "10010001",20073 => "11110101",20074 => "00101100",20075 => "00000000",20076 => "00101101",20077 => "01001110",20078 => "01001110",20079 => "00011000",20080 => "00111001",20081 => "11001011",20082 => "01011000",20083 => "10111110",20084 => "01111111",20085 => "10000111",20086 => "01101000",20087 => "10000100",20088 => "00100111",20089 => "11111100",20090 => "00100100",20091 => "11011111",20092 => "01101000",20093 => "00011100",20094 => "01000111",20095 => "01000111",20096 => "11111100",20097 => "11110001",20098 => "01101101",20099 => "00010101",20100 => "01000010",20101 => "11000101",20102 => "10001111",20103 => "00011110",20104 => "11110001",20105 => "11100110",20106 => "00111111",20107 => "10000101",20108 => "01011110",20109 => "10010111",20110 => "10101101",20111 => "00011010",20112 => "10101011",20113 => "11110111",20114 => "11111110",20115 => "00011010",20116 => "00111001",20117 => "11000100",20118 => "01111101",20119 => "10001100",20120 => "10011000",20121 => "11011000",20122 => "10111011",20123 => "11101010",20124 => "11010001",20125 => "01001111",20126 => "11000100",20127 => "01011010",20128 => "00000010",20129 => "10000001",20130 => "01110100",20131 => "10000100",20132 => "10010010",20133 => "01101011",20134 => "01001111",20135 => "11001000",20136 => "01110110",20137 => "11110110",20138 => "01101001",20139 => "01000101",20140 => "00100101",20141 => "10010011",20142 => "01100010",20143 => "01001001",20144 => "00001101",20145 => "01101110",20146 => "00101001",20147 => "10011001",20148 => "00011111",20149 => "00111101",20150 => "00011101",20151 => "11000010",20152 => "00001100",20153 => "11100110",20154 => "01100101",20155 => "10011110",20156 => "11100010",20157 => "01001100",20158 => "11111101",20159 => "00101101",20160 => "10110100",20161 => "01000010",20162 => "10101011",20163 => "10000010",20164 => "00010111",20165 => "01101010",20166 => "00101111",20167 => "10010111",20168 => "10010000",20169 => "01000110",20170 => "10110111",20171 => "00111010",20172 => "11100100",20173 => "11010001",20174 => "10011110",20175 => "11110100",20176 => "11111000",20177 => "00010011",20178 => "10000110",20179 => "00110011",20180 => "10001000",20181 => "00110000",20182 => "10011001",20183 => "11101000",20184 => "10010110",20185 => "00011101",20186 => "00010101",20187 => "00111000",20188 => "00010001",20189 => "11010000",20190 => "01011110",20191 => "01110100",20192 => "00101100",20193 => "10001110",20194 => "00100100",20195 => "00100010",20196 => "10001101",20197 => "00010001",20198 => "00000000",20199 => "01011011",20200 => "11110100",20201 => "01101011",20202 => "01000111",20203 => "10011100",20204 => "10110101",20205 => "00110101",20206 => "01100000",20207 => "11110000",20208 => "01001010",20209 => "10111000",20210 => "01100010",20211 => "00010100",20212 => "00000100",20213 => "11011010",20214 => "00100000",20215 => "01111101",20216 => "11110001",20217 => "10000100",20218 => "00100110",20219 => "10110100",20220 => "10100110",20221 => "00110101",20222 => "00110110",20223 => "10111110",20224 => "10101110",20225 => "10010111",20226 => "10010100",20227 => "01101000",20228 => "00100010",20229 => "00100001",20230 => "00001110",20231 => "00101100",20232 => "00000111",20233 => "10001100",20234 => "01011011",20235 => "01100001",20236 => "11110001",20237 => "00000010",20238 => "01100101",20239 => "10010111",20240 => "10110100",20241 => "11100011",20242 => "11000010",20243 => "11011100",20244 => "10100001",20245 => "10100011",20246 => "10111000",20247 => "00011000",20248 => "01101101",20249 => "01111111",20250 => "10100100",20251 => "01000110",20252 => "00111110",20253 => "11110111",20254 => "10110011",20255 => "00110010",20256 => "00001001",20257 => "00111010",20258 => "11100000",20259 => "11110011",20260 => "01000110",20261 => "00110011",20262 => "11101011",20263 => "10111110",20264 => "11100001",20265 => "01000010",20266 => "10001101",20267 => "00111000",20268 => "11010111",20269 => "00000010",20270 => "11111111",20271 => "01110001",20272 => "00001101",20273 => "00001101",20274 => "11111111",20275 => "10000011",20276 => "01101001",20277 => "00000001",20278 => "11001111",20279 => "01001100",20280 => "11110100",20281 => "10001011",20282 => "01010100",20283 => "01001101",20284 => "10110011",20285 => "00111100",20286 => "10110101",20287 => "00111111",20288 => "10001001",20289 => "10000001",20290 => "10100111",20291 => "11010000",20292 => "01011000",20293 => "10110001",20294 => "10111011",20295 => "10001111",20296 => "11001111",20297 => "10111010",20298 => "01110110",20299 => "10011010",20300 => "00111100",20301 => "11001000",20302 => "00110100",20303 => "01101111",20304 => "00101010",20305 => "11010110",20306 => "10011010",20307 => "01001110",20308 => "00100110",20309 => "11101000",20310 => "01101100",20311 => "00011011",20312 => "10000100",20313 => "00101100",20314 => "11100110",20315 => "01101111",20316 => "01011100",20317 => "10011110",20318 => "10111000",20319 => "00011011",20320 => "01010000",20321 => "01000000",20322 => "01010111",20323 => "01100100",20324 => "10011001",20325 => "11011111",20326 => "10100010",20327 => "01001100",20328 => "11111111",20329 => "01001001",20330 => "10111111",20331 => "10111001",20332 => "00101100",20333 => "00101010",20334 => "11010001",20335 => "10111001",20336 => "10111010",20337 => "00000010",20338 => "11000100",20339 => "10101100",20340 => "11111111",20341 => "01111111",20342 => "11101001",20343 => "00000111",20344 => "11101110",20345 => "01001100",20346 => "01101110",20347 => "10110110",20348 => "11000100",20349 => "01000010",20350 => "11000111",20351 => "00111100",20352 => "01001000",20353 => "11000110",20354 => "01010111",20355 => "00101010",20356 => "10111011",20357 => "00001100",20358 => "11010010",20359 => "00110101",20360 => "11100011",20361 => "01001000",20362 => "00001101",20363 => "00010001",20364 => "10101101",20365 => "00110110",20366 => "11100101",20367 => "01010001",20368 => "10100110",20369 => "11011101",20370 => "00010110",20371 => "11100110",20372 => "01001010",20373 => "00111011",20374 => "01110010",20375 => "01001000",20376 => "01011111",20377 => "11110101",20378 => "10100010",20379 => "11001000",20380 => "00010110",20381 => "01011111",20382 => "10010011",20383 => "00000100",20384 => "00111110",20385 => "11111101",20386 => "11111011",20387 => "00001111",20388 => "10100101",20389 => "00010011",20390 => "10101110",20391 => "11001000",20392 => "10001000",20393 => "11010100",20394 => "01101111",20395 => "11001011",20396 => "01110010",20397 => "01000011",20398 => "01101100",20399 => "01001010",20400 => "00010011",20401 => "00111101",20402 => "10001110",20403 => "11111011",20404 => "10100111",20405 => "10001100",20406 => "10101111",20407 => "11011100",20408 => "10100000",20409 => "11011011",20410 => "00010010",20411 => "01111100",20412 => "11101110",20413 => "10000101",20414 => "11010110",20415 => "11001000",20416 => "10010100",20417 => "01101011",20418 => "01010101",20419 => "10110110",20420 => "00100011",20421 => "01110000",20422 => "11111101",20423 => "11010110",20424 => "00011101",20425 => "01010101",20426 => "11000110",20427 => "01100100",20428 => "11000111",20429 => "10100110",20430 => "00110010",20431 => "00010011",20432 => "10101010",20433 => "01010011",20434 => "11010111",20435 => "10001000",20436 => "11100110",20437 => "00011110",20438 => "11011010",20439 => "01111110",20440 => "10110100",20441 => "10001000",20442 => "11000011",20443 => "01100101",20444 => "01000111",20445 => "01110101",20446 => "10011001",20447 => "00110000",20448 => "11110100",20449 => "10011011",20450 => "00101110",20451 => "00000011",20452 => "10001101",20453 => "00101111",20454 => "01111000",20455 => "00101111",20456 => "01100011",20457 => "11010101",20458 => "10000000",20459 => "10001110",20460 => "10000110",20461 => "10001010",20462 => "00111110",20463 => "11000101",20464 => "01111001",20465 => "00111101",20466 => "00000000",20467 => "11100010",20468 => "11101110",20469 => "11110100",20470 => "00111101",20471 => "10101100",20472 => "10001010",20473 => "01101101",20474 => "00011011",20475 => "11111110",20476 => "01001101",20477 => "10101011",20478 => "11100010",20479 => "00000011",20480 => "11101000",20481 => "11110001",20482 => "11101000",20483 => "11001001",20484 => "10011010",20485 => "01000110",20486 => "01001010",20487 => "11110000",20488 => "00011101",20489 => "10010110",20490 => "11001110",20491 => "11011100",20492 => "01110011",20493 => "01101110",20494 => "10011100",20495 => "11001110",20496 => "11111101",20497 => "11100001",20498 => "00101101",20499 => "01000000",20500 => "01110101",20501 => "11001000",20502 => "00101111",20503 => "00100100",20504 => "01010100",20505 => "11100110",20506 => "11001010",20507 => "10000111",20508 => "11001101",20509 => "11011110",20510 => "10110111",20511 => "11000011",20512 => "00010110",20513 => "00011010",20514 => "10111101",20515 => "10110011",20516 => "10110100",20517 => "00001110",20518 => "00001000",20519 => "10000101",20520 => "10011101",20521 => "10110011",20522 => "11110010",20523 => "00100100",20524 => "11101010",20525 => "00110000",20526 => "01001111",20527 => "01010101",20528 => "00100010",20529 => "00010110",20530 => "10011111",20531 => "00000010",20532 => "01101110",20533 => "00011101",20534 => "00010010",20535 => "11011101",20536 => "00001111",20537 => "00010000",20538 => "00100111",20539 => "10101010",20540 => "01100100",20541 => "11010000",20542 => "01111000",20543 => "01001110",20544 => "00101011",20545 => "10010011",20546 => "10001111",20547 => "00011011",20548 => "11100111",20549 => "11000100",20550 => "01101010",20551 => "00101000",20552 => "10100000",20553 => "01110011",20554 => "01111101",20555 => "10001000",20556 => "00010101",20557 => "00001110",20558 => "11100100",20559 => "01000011",20560 => "00111011",20561 => "10101011",20562 => "11010011",20563 => "00010110",20564 => "01110100",20565 => "11001011",20566 => "00000101",20567 => "00110110",20568 => "00000010",20569 => "01000001",20570 => "00100011",20571 => "10010001",20572 => "10111000",20573 => "10011011",20574 => "10101111",20575 => "00011111",20576 => "00000111",20577 => "10010110",20578 => "00100011",20579 => "11001000",20580 => "10010101",20581 => "11001000",20582 => "00110010",20583 => "11011110",20584 => "00111101",20585 => "01100001",20586 => "10100010",20587 => "11001000",20588 => "11001110",20589 => "01100010",20590 => "11011101",20591 => "11110001",20592 => "01110100",20593 => "01001101",20594 => "10000101",20595 => "11010000",20596 => "01111101",20597 => "11100100",20598 => "10000010",20599 => "11101001",20600 => "01001110",20601 => "01111000",20602 => "11001101",20603 => "01011100",20604 => "11101010",20605 => "01000111",20606 => "11101000",20607 => "00111100",20608 => "00001111",20609 => "11110011",20610 => "00001001",20611 => "11111001",20612 => "10100010",20613 => "11000010",20614 => "01000100",20615 => "10110111",20616 => "10011000",20617 => "00011010",20618 => "10110010",20619 => "00100100",20620 => "01101010",20621 => "10000000",20622 => "00110001",20623 => "10001101",20624 => "11101111",20625 => "00011000",20626 => "10000001",20627 => "10100010",20628 => "10011110",20629 => "01001010",20630 => "11000001",20631 => "11100101",20632 => "01001001",20633 => "10000010",20634 => "00110010",20635 => "10010100",20636 => "11001100",20637 => "01001000",20638 => "10010001",20639 => "01111000",20640 => "00100001",20641 => "00011110",20642 => "10000001",20643 => "00111010",20644 => "00010001",20645 => "01000000",20646 => "01101010",20647 => "10001000",20648 => "00100001",20649 => "11001000",20650 => "00000100",20651 => "10010110",20652 => "00100111",20653 => "01001001",20654 => "11101101",20655 => "00111100",20656 => "01101100",20657 => "01011100",20658 => "00101000",20659 => "11101011",20660 => "01110001",20661 => "01001001",20662 => "11010001",20663 => "01011011",20664 => "10110001",20665 => "01010011",20666 => "00111111",20667 => "01000011",20668 => "10000010",20669 => "11000010",20670 => "11110000",20671 => "10010010",20672 => "01110011",20673 => "01111011",20674 => "00010001",20675 => "10110010",20676 => "11100011",20677 => "10001010",20678 => "00001011",20679 => "01101101",20680 => "01110001",20681 => "01111100",20682 => "10101011",20683 => "11111111",20684 => "00010100",20685 => "00011101",20686 => "11110010",20687 => "10111111",20688 => "00110001",20689 => "00001111",20690 => "01100100",20691 => "01011111",20692 => "00111010",20693 => "00100100",20694 => "01101100",20695 => "00011011",20696 => "00100000",20697 => "01001011",20698 => "01011101",20699 => "01111100",20700 => "11001001",20701 => "01011100",20702 => "11011001",20703 => "01111111",20704 => "10000000",20705 => "10111010",20706 => "00011110",20707 => "10110001",20708 => "10001010",20709 => "11010010",20710 => "01000101",20711 => "11110010",20712 => "00001100",20713 => "01100010",20714 => "10010000",20715 => "11111111",20716 => "10111000",20717 => "01101000",20718 => "01000111",20719 => "01010110",20720 => "10000010",20721 => "01011110",20722 => "11011111",20723 => "00010101",20724 => "10100000",20725 => "01001101",20726 => "00110111",20727 => "00111110",20728 => "10011100",20729 => "10010110",20730 => "00100011",20731 => "10111011",20732 => "11101110",20733 => "00001100",20734 => "11011110",20735 => "11110010",20736 => "10011010",20737 => "10110101",20738 => "11010110",20739 => "00100111",20740 => "10000011",20741 => "11010111",20742 => "10100011",20743 => "10101010",20744 => "01011010",20745 => "11111110",20746 => "00010001",20747 => "00111001",20748 => "01101010",20749 => "10001010",20750 => "10110111",20751 => "10111011",20752 => "00101010",20753 => "00111011",20754 => "10000000",20755 => "01111001",20756 => "00001101",20757 => "00000111",20758 => "11111001",20759 => "00010011",20760 => "01110111",20761 => "11001010",20762 => "00000111",20763 => "00010111",20764 => "10101001",20765 => "11110001",20766 => "11001001",20767 => "10111000",20768 => "10010011",20769 => "11101111",20770 => "00111001",20771 => "01101010",20772 => "11011110",20773 => "01011101",20774 => "00001011",20775 => "10101011",20776 => "11010001",20777 => "10101011",20778 => "00001100",20779 => "10110010",20780 => "01010101",20781 => "01101110",20782 => "11010100",20783 => "11011100",20784 => "00111110",20785 => "00100110",20786 => "10010110",20787 => "01100100",20788 => "10111000",20789 => "11000101",20790 => "11001011",20791 => "01101110",20792 => "00110101",20793 => "00001100",20794 => "11111010",20795 => "01000011",20796 => "00111010",20797 => "10111010",20798 => "01110010",20799 => "10110101",20800 => "11011111",20801 => "11100101",20802 => "01111110",20803 => "01111100",20804 => "01001001",20805 => "10100010",20806 => "11001000",20807 => "00111110",20808 => "00100101",20809 => "00001001",20810 => "00001100",20811 => "11000101",20812 => "01011011",20813 => "11111011",20814 => "11000010",20815 => "00001111",20816 => "00011110",20817 => "01011110",20818 => "11101011",20819 => "00000111",20820 => "10010001",20821 => "10111100",20822 => "10101110",20823 => "00101011",20824 => "00001000",20825 => "01100100",20826 => "11001010",20827 => "10001000",20828 => "01011111",20829 => "00110010",20830 => "01011001",20831 => "10110111",20832 => "10000010",20833 => "00001001",20834 => "01000011",20835 => "10110000",20836 => "00101000",20837 => "00010111",20838 => "00010011",20839 => "00000010",20840 => "11001000",20841 => "11011111",20842 => "11110101",20843 => "00001010",20844 => "10000100",20845 => "10111100",20846 => "01101000",20847 => "00110110",20848 => "10001111",20849 => "10001011",20850 => "11110001",20851 => "00100110",20852 => "11110001",20853 => "10001111",20854 => "01111110",20855 => "10001011",20856 => "11111110",20857 => "11010011",20858 => "01110011",20859 => "00101111",20860 => "01111110",20861 => "10101000",20862 => "00110100",20863 => "11001011",20864 => "00110110",20865 => "00100110",20866 => "00111110",20867 => "00101001",20868 => "11011011",20869 => "00111011",20870 => "01110110",20871 => "00100110",20872 => "10000000",20873 => "01011101",20874 => "11101100",20875 => "10000100",20876 => "11011111",20877 => "01000101",20878 => "00110100",20879 => "10010011",20880 => "00101101",20881 => "00110000",20882 => "11000000",20883 => "11001001",20884 => "01011000",20885 => "01101111",20886 => "10110101",20887 => "00110110",20888 => "01101110",20889 => "11001010",20890 => "10001101",20891 => "01011100",20892 => "10111101",20893 => "00101010",20894 => "11100010",20895 => "10110011",20896 => "01111110",20897 => "10100110",20898 => "00000111",20899 => "11000000",20900 => "10000111",20901 => "01110110",20902 => "00000101",20903 => "10100011",20904 => "01111101",20905 => "10110101",20906 => "00101100",20907 => "01110001",20908 => "11001111",20909 => "11101100",20910 => "00011101",20911 => "00001111",20912 => "10000110",20913 => "11110001",20914 => "11110010",20915 => "11000011",20916 => "11100110",20917 => "10010010",20918 => "01001101",20919 => "10100110",20920 => "10101100",20921 => "11001111",20922 => "01100111",20923 => "10011101",20924 => "01100101",20925 => "00100000",20926 => "00101011",20927 => "00010101",20928 => "10010001",20929 => "00101011",20930 => "10101010",20931 => "11001100",20932 => "01101111",20933 => "01010101",20934 => "00001000",20935 => "01100101",20936 => "10001100",20937 => "00000011",20938 => "01100101",20939 => "11001010",20940 => "11100000",20941 => "00000110",20942 => "01101110",20943 => "00100101",20944 => "10001111",20945 => "01110100",20946 => "00000100",20947 => "00110111",20948 => "11100110",20949 => "11111011",20950 => "01100011",20951 => "00111010",20952 => "00001010",20953 => "10101010",20954 => "10101101",20955 => "00000111",20956 => "11101010",20957 => "10111011",20958 => "00001011",20959 => "11011111",20960 => "11001101",20961 => "00000110",20962 => "00111111",20963 => "00010011",20964 => "11000010",20965 => "11000100",20966 => "10100110",20967 => "10111011",20968 => "00101011",20969 => "10000100",20970 => "11010110",20971 => "01100001",20972 => "10001110",20973 => "00101101",20974 => "11111011",20975 => "00010010",20976 => "11110111",20977 => "10000101",20978 => "01000011",20979 => "01001010",20980 => "11001111",20981 => "11001000",20982 => "10101111",20983 => "10111110",20984 => "00110000",20985 => "10011001",20986 => "10010011",20987 => "11110111",20988 => "10111011",20989 => "00111111",20990 => "00111101",20991 => "01110100",20992 => "10011011",20993 => "00100101",20994 => "10010101",20995 => "01011001",20996 => "01110110",20997 => "10111000",20998 => "00001000",20999 => "00110111",21000 => "11100001",21001 => "11111011",21002 => "10101110",21003 => "00100011",21004 => "10101010",21005 => "00000000",21006 => "10011011",21007 => "10100000",21008 => "10000100",21009 => "11010111",21010 => "01100010",21011 => "10101111",21012 => "00111100",21013 => "10010011",21014 => "11110010",21015 => "01101101",21016 => "11001001",21017 => "01111001",21018 => "10111001",21019 => "00010001",21020 => "00011000",21021 => "10001111",21022 => "00010011",21023 => "11010111",21024 => "00010111",21025 => "00010000",21026 => "00100110",21027 => "11011010",21028 => "00110110",21029 => "11111010",21030 => "01011010",21031 => "00111110",21032 => "00110001",21033 => "01010001",21034 => "00110010",21035 => "10011111",21036 => "11010011",21037 => "10010011",21038 => "10101110",21039 => "00001001",21040 => "11101101",21041 => "11100000",21042 => "01111000",21043 => "01000001",21044 => "01010110",21045 => "11101011",21046 => "00101101",21047 => "00000010",21048 => "01100000",21049 => "00111101",21050 => "01110011",21051 => "10010001",21052 => "10101011",21053 => "10010101",21054 => "00010111",21055 => "11011001",21056 => "00110111",21057 => "01110001",21058 => "00000010",21059 => "11110100",21060 => "10001101",21061 => "10100011",21062 => "11011110",21063 => "00000110",21064 => "11010110",21065 => "10000011",21066 => "10100001",21067 => "11011010",21068 => "00101100",21069 => "11110010",21070 => "10010111",21071 => "11111101",21072 => "10111011",21073 => "10010110",21074 => "11000001",21075 => "10101110",21076 => "11110101",21077 => "00010000",21078 => "10001001",21079 => "00111000",21080 => "01100110",21081 => "00110011",21082 => "10001101",21083 => "00101010",21084 => "00001100",21085 => "01101111",21086 => "10110110",21087 => "01101010",21088 => "11111011",21089 => "01100001",21090 => "10100110",21091 => "10110111",21092 => "10100001",21093 => "00001110",21094 => "10100101",21095 => "01101011",21096 => "11110100",21097 => "01101000",21098 => "10011111",21099 => "10011001",21100 => "00111010",21101 => "01100010",21102 => "11100000",21103 => "01011110",21104 => "01100100",21105 => "01001101",21106 => "11011111",21107 => "11101111",21108 => "10000100",21109 => "01000111",21110 => "00001111",21111 => "00110111",21112 => "01101010",21113 => "10111111",21114 => "11111110",21115 => "10101000",21116 => "01001010",21117 => "01001000",21118 => "11010010",21119 => "01101001",21120 => "01110101",21121 => "01010101",21122 => "10000101",21123 => "10011100",21124 => "11110100",21125 => "00010010",21126 => "10110101",21127 => "01101101",21128 => "01110000",21129 => "10100111",21130 => "11010101",21131 => "01011111",21132 => "11100000",21133 => "00010001",21134 => "00110000",21135 => "10010010",21136 => "01110001",21137 => "00010100",21138 => "11001111",21139 => "01011001",21140 => "00111100",21141 => "10100010",21142 => "11000001",21143 => "10101001",21144 => "01001000",21145 => "00100000",21146 => "10001100",21147 => "11110101",21148 => "11001110",21149 => "10011101",21150 => "01001101",21151 => "10110001",21152 => "01110001",21153 => "10110111",21154 => "11001001",21155 => "10001101",21156 => "10011000",21157 => "11011001",21158 => "11011000",21159 => "10001100",21160 => "00001011",21161 => "11100101",21162 => "00101100",21163 => "10010111",21164 => "10110010",21165 => "11111011",21166 => "00001000",21167 => "10100001",21168 => "10101101",21169 => "10110110",21170 => "10000101",21171 => "01000011",21172 => "11001001",21173 => "11100100",21174 => "11000001",21175 => "10001100",21176 => "01000101",21177 => "00101010",21178 => "00110110",21179 => "01000000",21180 => "00010101",21181 => "00100101",21182 => "01111111",21183 => "10001010",21184 => "11101101",21185 => "01100010",21186 => "10000110",21187 => "11001101",21188 => "11110111",21189 => "11001000",21190 => "01011101",21191 => "00010011",21192 => "00110011",21193 => "01011100",21194 => "11111010",21195 => "01101001",21196 => "10110101",21197 => "00101100",21198 => "10010110",21199 => "10110100",21200 => "00111101",21201 => "00110000",21202 => "01100111",21203 => "00000011",21204 => "11100111",21205 => "00100010",21206 => "00110101",21207 => "00110101",21208 => "11111000",21209 => "11100000",21210 => "00000100",21211 => "11110101",21212 => "11100100",21213 => "01101101",21214 => "11100010",21215 => "11000001",21216 => "10111011",21217 => "01100110",21218 => "11101111",21219 => "01010000",21220 => "11101010",21221 => "10111011",21222 => "10011111",21223 => "01110010",21224 => "01100100",21225 => "10110001",21226 => "01000101",21227 => "10010000",21228 => "10010111",21229 => "10010111",21230 => "10110101",21231 => "10011100",21232 => "01001101",21233 => "11100101",21234 => "10001100",21235 => "01001111",21236 => "01010100",21237 => "00101111",21238 => "10001101",21239 => "11000000",21240 => "10000001",21241 => "11000000",21242 => "00110010",21243 => "10011111",21244 => "01001111",21245 => "00101111",21246 => "01001100",21247 => "11001111",21248 => "10011010",21249 => "11101100",21250 => "01110110",21251 => "00001111",21252 => "01110001",21253 => "01000001",21254 => "01000100",21255 => "00011101",21256 => "10101110",21257 => "00000001",21258 => "10111010",21259 => "10111100",21260 => "00000001",21261 => "00010011",21262 => "01111101",21263 => "01011011",21264 => "00101111",21265 => "10000010",21266 => "10101000",21267 => "01101111",21268 => "11111101",21269 => "00110001",21270 => "10100001",21271 => "10010001",21272 => "01011001",21273 => "11111101",21274 => "01011010",21275 => "01101010",21276 => "00100110",21277 => "01000100",21278 => "01000101",21279 => "00001010",21280 => "01111111",21281 => "00110010",21282 => "11100000",21283 => "00111000",21284 => "01100001",21285 => "11110110",21286 => "11010001",21287 => "00010001",21288 => "10100010",21289 => "00011110",21290 => "00100111",21291 => "01101101",21292 => "10101101",21293 => "11101000",21294 => "01110001",21295 => "10110010",21296 => "01001101",21297 => "00010010",21298 => "11011100",21299 => "11001000",21300 => "11010000",21301 => "11010011",21302 => "11011110",21303 => "00110100",21304 => "11100001",21305 => "01111010",21306 => "00111000",21307 => "11110000",21308 => "01000110",21309 => "01111000",21310 => "11010111",21311 => "10011110",21312 => "01011000",21313 => "01100100",21314 => "10101001",21315 => "11000100",21316 => "00010011",21317 => "00001001",21318 => "01110001",21319 => "01000001",21320 => "10010001",21321 => "00010111",21322 => "01001011",21323 => "01100100",21324 => "00001000",21325 => "10000001",21326 => "01111110",21327 => "00110010",21328 => "01010101",21329 => "00011110",21330 => "01000011",21331 => "00111000",21332 => "01111111",21333 => "01011010",21334 => "00110000",21335 => "00001111",21336 => "01101100",21337 => "01101000",21338 => "00100011",21339 => "11000000",21340 => "11001101",21341 => "01011110",21342 => "10011011",21343 => "11000010",21344 => "11001000",21345 => "01011001",21346 => "10000000",21347 => "10100111",21348 => "01000010",21349 => "10101001",21350 => "00010001",21351 => "11100100",21352 => "00110100",21353 => "11010101",21354 => "01100011",21355 => "00011110",21356 => "00010011",21357 => "01010010",21358 => "11000011",21359 => "11000110",21360 => "11011100",21361 => "10000111",21362 => "00000110",21363 => "10010101",21364 => "11000100",21365 => "00011010",21366 => "00000011",21367 => "00100010",21368 => "11101000",21369 => "11101001",21370 => "11110000",21371 => "00000000",21372 => "00011011",21373 => "01100110",21374 => "10100000",21375 => "11100000",21376 => "11010100",21377 => "00000011",21378 => "11000011",21379 => "00110100",21380 => "10101111",21381 => "11100001",21382 => "01110000",21383 => "11000100",21384 => "10001100",21385 => "01000011",21386 => "01110010",21387 => "10001000",21388 => "11110100",21389 => "10100111",21390 => "11011100",21391 => "11001101",21392 => "11010111",21393 => "10011110",21394 => "11100011",21395 => "01000110",21396 => "10000010",21397 => "01011110",21398 => "11110100",21399 => "11010011",21400 => "00011110",21401 => "11100100",21402 => "00011100",21403 => "10100000",21404 => "01100011",21405 => "01101011",21406 => "10000001",21407 => "11001001",21408 => "00110001",21409 => "10011110",21410 => "00000001",21411 => "01011100",21412 => "10011001",21413 => "00110011",21414 => "00111101",21415 => "11000111",21416 => "11000011",21417 => "00111000",21418 => "00111010",21419 => "01111101",21420 => "10110110",21421 => "01011011",21422 => "11100000",21423 => "00101101",21424 => "10101011",21425 => "10111011",21426 => "10100100",21427 => "00110100",21428 => "01101011",21429 => "10110110",21430 => "00110010",21431 => "11101111",21432 => "00001101",21433 => "10001100",21434 => "10011101",21435 => "11110000",21436 => "01001111",21437 => "01011011",21438 => "11101110",21439 => "11100111",21440 => "01100101",21441 => "11000011",21442 => "01010010",21443 => "11101001",21444 => "10010100",21445 => "01010010",21446 => "01100000",21447 => "11101100",21448 => "10001111",21449 => "01010000",21450 => "00001100",21451 => "00111110",21452 => "11100101",21453 => "11111011",21454 => "10111110",21455 => "10101010",21456 => "11010011",21457 => "10010011",21458 => "01010010",21459 => "10010101",21460 => "11110000",21461 => "01101101",21462 => "11101010",21463 => "11110111",21464 => "01111111",21465 => "00001010",21466 => "01111011",21467 => "00110011",21468 => "01010100",21469 => "01110000",21470 => "10110011",21471 => "10101001",21472 => "00101100",21473 => "01111000",21474 => "00010010",21475 => "01011010",21476 => "11011100",21477 => "11101100",21478 => "10100000",21479 => "00011100",21480 => "00111100",21481 => "11010010",21482 => "01110010",21483 => "11110111",21484 => "00110100",21485 => "01010100",21486 => "00001001",21487 => "00010010",21488 => "01101010",21489 => "01100010",21490 => "00101000",21491 => "01001011",21492 => "11000010",21493 => "10000011",21494 => "00010001",21495 => "10111111",21496 => "10100110",21497 => "11101001",21498 => "11101110",21499 => "11101010",21500 => "10000101",21501 => "01101001",21502 => "10000010",21503 => "00011000",21504 => "00101010",21505 => "11101000",21506 => "01010011",21507 => "00011000",21508 => "00111100",21509 => "01000010",21510 => "10011111",21511 => "00011001",21512 => "01011100",21513 => "10101011",21514 => "10011010",21515 => "00010011",21516 => "00011100",21517 => "11000000",21518 => "11000011",21519 => "01010100",21520 => "11101000",21521 => "10011000",21522 => "00010110",21523 => "00111000",21524 => "01101001",21525 => "11101011",21526 => "11101000",21527 => "00101011",21528 => "10101001",21529 => "01010100",21530 => "01011010",21531 => "00101001",21532 => "11110001",21533 => "10001010",21534 => "11010101",21535 => "11000001",21536 => "10000100",21537 => "01000101",21538 => "11110101",21539 => "01100000",21540 => "10011000",21541 => "00110000",21542 => "00001001",21543 => "01110101",21544 => "10010001",21545 => "10111100",21546 => "11110011",21547 => "00110010",21548 => "10000111",21549 => "00110010",21550 => "01110101",21551 => "10000011",21552 => "00001111",21553 => "00100011",21554 => "11111000",21555 => "01000001",21556 => "10100001",21557 => "10000011",21558 => "10000000",21559 => "01010001",21560 => "00111110",21561 => "11100011",21562 => "11001011",21563 => "11100111",21564 => "11101110",21565 => "00011011",21566 => "00101010",21567 => "01100000",21568 => "10101011",21569 => "11100000",21570 => "11010111",21571 => "00101011",21572 => "10110011",21573 => "11001001",21574 => "00100000",21575 => "00011000",21576 => "01010110",21577 => "00110100",21578 => "01001110",21579 => "10000001",21580 => "01101001",21581 => "11100100",21582 => "11001011",21583 => "10111010",21584 => "01111000",21585 => "10010000",21586 => "11100110",21587 => "10011001",21588 => "10010001",21589 => "10001100",21590 => "01101011",21591 => "01001000",21592 => "11110000",21593 => "10010111",21594 => "11101011",21595 => "00100110",21596 => "10100000",21597 => "00101000",21598 => "00100001",21599 => "10010111",21600 => "11010001",21601 => "01110001",21602 => "01010000",21603 => "00110101",21604 => "10001000",21605 => "11010011",21606 => "00101100",21607 => "01010000",21608 => "11111100",21609 => "10001110",21610 => "10001010",21611 => "01001101",21612 => "00111100",21613 => "00011011",21614 => "01111111",21615 => "01110111",21616 => "10010010",21617 => "00011101",21618 => "00101010",21619 => "10111111",21620 => "00011010",21621 => "00001101",21622 => "00010010",21623 => "00101001",21624 => "01000001",21625 => "10001001",21626 => "11000011",21627 => "00001110",21628 => "10110111",21629 => "10101010",21630 => "11000001",21631 => "00001001",21632 => "11100100",21633 => "01010101",21634 => "00000111",21635 => "01011100",21636 => "10001100",21637 => "10011110",21638 => "10111101",21639 => "11000100",21640 => "10011111",21641 => "00001100",21642 => "11111000",21643 => "10101110",21644 => "00100110",21645 => "10011110",21646 => "11000100",21647 => "11010110",21648 => "01111100",21649 => "00011110",21650 => "00000001",21651 => "01010001",21652 => "10100100",21653 => "11000000",21654 => "11001110",21655 => "10101101",21656 => "00110001",21657 => "11000001",21658 => "11001010",21659 => "00111000",21660 => "10111101",21661 => "01111101",21662 => "01001011",21663 => "10111011",21664 => "11101010",21665 => "00100001",21666 => "00010001",21667 => "01010100",21668 => "00011011",21669 => "00001110",21670 => "10101001",21671 => "01110111",21672 => "00100101",21673 => "10111110",21674 => "01010001",21675 => "11101111",21676 => "00111011",21677 => "01011001",21678 => "01100011",21679 => "11000100",21680 => "11011110",21681 => "10000011",21682 => "00011100",21683 => "01101011",21684 => "01101110",21685 => "11100001",21686 => "11111000",21687 => "10010100",21688 => "01110110",21689 => "00110101",21690 => "01110000",21691 => "11100101",21692 => "01101000",21693 => "10111101",21694 => "10010100",21695 => "11011000",21696 => "11100101",21697 => "01001111",21698 => "01110101",21699 => "11101101",21700 => "11111101",21701 => "11011001",21702 => "11010101",21703 => "01110001",21704 => "01000000",21705 => "11011101",21706 => "00011011",21707 => "01111100",21708 => "11110111",21709 => "01101000",21710 => "10111110",21711 => "11010100",21712 => "11111001",21713 => "01111100",21714 => "10010010",21715 => "00011110",21716 => "10101011",21717 => "00000010",21718 => "01011111",21719 => "00111001",21720 => "00110111",21721 => "11000110",21722 => "01001011",21723 => "11101011",21724 => "11001110",21725 => "11011111",21726 => "11000010",21727 => "11111100",21728 => "00010001",21729 => "00001001",21730 => "11001001",21731 => "01100001",21732 => "11000100",21733 => "00110001",21734 => "11000100",21735 => "11110001",21736 => "11100110",21737 => "11001101",21738 => "11010100",21739 => "01000101",21740 => "00110010",21741 => "01111111",21742 => "00101011",21743 => "11011101",21744 => "11001101",21745 => "10010011",21746 => "00110000",21747 => "10110000",21748 => "10110111",21749 => "10101001",21750 => "11110111",21751 => "00000111",21752 => "00101110",21753 => "11110001",21754 => "00000101",21755 => "11111011",21756 => "00001111",21757 => "00101110",21758 => "11100101",21759 => "10111111",21760 => "01011101",21761 => "01000011",21762 => "11001101",21763 => "00101110",21764 => "11110001",21765 => "10100100",21766 => "00110010",21767 => "10111100",21768 => "00111101",21769 => "10110011",21770 => "00100110",21771 => "01100101",21772 => "01101010",21773 => "11111110",21774 => "11001000",21775 => "00000001",21776 => "00110011",21777 => "11011011",21778 => "01000111",21779 => "10110111",21780 => "01100011",21781 => "01110001",21782 => "00011011",21783 => "10101011",21784 => "01011101",21785 => "10100110",21786 => "11101011",21787 => "01100110",21788 => "01011010",21789 => "01000000",21790 => "10111111",21791 => "00111100",21792 => "01000000",21793 => "00111100",21794 => "10101011",21795 => "01001100",21796 => "10011000",21797 => "11111111",21798 => "11001000",21799 => "11001110",21800 => "10100100",21801 => "10001000",21802 => "10100010",21803 => "00001111",21804 => "10111010",21805 => "00011010",21806 => "11001101",21807 => "01111110",21808 => "00000000",21809 => "01111110",21810 => "11010011",21811 => "10011111",21812 => "11000100",21813 => "11100000",21814 => "10000001",21815 => "11000100",21816 => "10110101",21817 => "00110011",21818 => "10101000",21819 => "10000111",21820 => "10001010",21821 => "11111100",21822 => "11011001",21823 => "10110011",21824 => "10011101",21825 => "00101101",21826 => "00111100",21827 => "01101000",21828 => "00001011",21829 => "10010110",21830 => "00011111",21831 => "00111101",21832 => "11111011",21833 => "01000010",21834 => "01100011",21835 => "10111111",21836 => "01001000",21837 => "11111000",21838 => "10010011",21839 => "11100011",21840 => "10001110",21841 => "01110011",21842 => "10010101",21843 => "01100101",21844 => "11110001",21845 => "01111111",21846 => "01000000",21847 => "01111010",21848 => "01010010",21849 => "11001000",21850 => "00100111",21851 => "10001000",21852 => "11101101",21853 => "00101111",21854 => "01001001",21855 => "10001100",21856 => "00000011",21857 => "00011111",21858 => "01111000",21859 => "11000101",21860 => "10100011",21861 => "00101110",21862 => "00010000",21863 => "10011011",21864 => "01011101",21865 => "01000001",21866 => "01111011",21867 => "01000011",21868 => "01111000",21869 => "10011101",21870 => "00010011",21871 => "01110010",21872 => "10100100",21873 => "01101100",21874 => "00001100",21875 => "10011100",21876 => "10101010",21877 => "01001001",21878 => "11110010",21879 => "10110101",21880 => "11101100",21881 => "00010000",21882 => "01011100",21883 => "00001011",21884 => "01101110",21885 => "01100010",21886 => "10011110",21887 => "01111010",21888 => "11010111",21889 => "01011101",21890 => "11110000",21891 => "01101000",21892 => "00010100",21893 => "01111010",21894 => "00111111",21895 => "01001011",21896 => "11001001",21897 => "00001001",21898 => "00000000",21899 => "01101110",21900 => "00101111",21901 => "01011100",21902 => "10011100",21903 => "01010101",21904 => "00110001",21905 => "00000110",21906 => "10100000",21907 => "11000100",21908 => "11000010",21909 => "00000101",21910 => "01100111",21911 => "10101110",21912 => "11001111",21913 => "01110000",21914 => "00111001",21915 => "10010111",21916 => "01000001",21917 => "00000111",21918 => "11101101",21919 => "01010000",21920 => "10000010",21921 => "10011111",21922 => "00101101",21923 => "11001011",21924 => "11010010",21925 => "10010100",21926 => "01001100",21927 => "10010101",21928 => "11010000",21929 => "01110100",21930 => "11111010",21931 => "11001101",21932 => "01111001",21933 => "10011111",21934 => "10000110",21935 => "11001101",21936 => "01001110",21937 => "10110111",21938 => "10100011",21939 => "11010101",21940 => "10111001",21941 => "00100101",21942 => "11000010",21943 => "00110110",21944 => "10000110",21945 => "10010010",21946 => "00110111",21947 => "10101101",21948 => "01101010",21949 => "00100100",21950 => "01110001",21951 => "01110110",21952 => "01110101",21953 => "10110111",21954 => "00001001",21955 => "01101110",21956 => "10001001",21957 => "01111011",21958 => "11011000",21959 => "00100100",21960 => "01111001",21961 => "01001011",21962 => "10100111",21963 => "00111011",21964 => "01100110",21965 => "11100011",21966 => "11110101",21967 => "00000000",21968 => "11110101",21969 => "11110111",21970 => "01011111",21971 => "00110000",21972 => "10000011",21973 => "11001100",21974 => "10011111",21975 => "00001001",21976 => "00001101",21977 => "10000101",21978 => "11111000",21979 => "11101011",21980 => "11101010",21981 => "01010100",21982 => "01001010",21983 => "11101110",21984 => "11010000",21985 => "11001011",21986 => "01110101",21987 => "00000001",21988 => "01110101",21989 => "11011110",21990 => "11100001",21991 => "11010111",21992 => "01110001",21993 => "00010011",21994 => "10101000",21995 => "01100010",21996 => "10000001",21997 => "11110001",21998 => "01101011",21999 => "01101001",22000 => "10010000",22001 => "00110000",22002 => "00010101",22003 => "00101011",22004 => "00100111",22005 => "10101000",22006 => "01101100",22007 => "00011001",22008 => "11100011",22009 => "11011100",22010 => "10000111",22011 => "01001111",22012 => "01101001",22013 => "00111101",22014 => "10000011",22015 => "10111010",22016 => "10100001",22017 => "11011100",22018 => "00001011",22019 => "00001101",22020 => "11100001",22021 => "10110010",22022 => "10001100",22023 => "00010101",22024 => "00111100",22025 => "01100001",22026 => "01111011",22027 => "00111011",22028 => "00110101",22029 => "00110100",22030 => "01011110",22031 => "10110011",22032 => "10101110",22033 => "10101001",22034 => "00000101",22035 => "11001000",22036 => "01000100",22037 => "11100010",22038 => "10101110",22039 => "01111000",22040 => "10110110",22041 => "11000000",22042 => "11100000",22043 => "00111110",22044 => "01101001",22045 => "00011010",22046 => "00011111",22047 => "11000101",22048 => "11100011",22049 => "11010010",22050 => "10101000",22051 => "01001101",22052 => "10101110",22053 => "00110010",22054 => "01100100",22055 => "11100100",22056 => "01010111",22057 => "10010011",22058 => "11100100",22059 => "10000000",22060 => "11011001",22061 => "10110001",22062 => "11111001",22063 => "11001011",22064 => "11111101",22065 => "11011100",22066 => "11101010",22067 => "00001111",22068 => "10000101",22069 => "10101110",22070 => "10100001",22071 => "00001100",22072 => "10101110",22073 => "11011001",22074 => "01000111",22075 => "01000010",22076 => "10011000",22077 => "11010100",22078 => "01100110",22079 => "11001100",22080 => "00100111",22081 => "10011110",22082 => "01000110",22083 => "00010000",22084 => "10001101",22085 => "10100100",22086 => "00110000",22087 => "11001011",22088 => "01110110",22089 => "00010101",22090 => "11111111",22091 => "00110110",22092 => "10100111",22093 => "00010010",22094 => "10110001",22095 => "00110001",22096 => "11111000",22097 => "10110100",22098 => "11101101",22099 => "01110110",22100 => "01100100",22101 => "01011001",22102 => "01111111",22103 => "00100110",22104 => "00001011",22105 => "10100100",22106 => "01010110",22107 => "11001110",22108 => "10111101",22109 => "10001010",22110 => "01000110",22111 => "01101100",22112 => "01101001",22113 => "11011011",22114 => "10000110",22115 => "11111111",22116 => "11000100",22117 => "11101011",22118 => "11011101",22119 => "10010000",22120 => "00000100",22121 => "00010010",22122 => "01110010",22123 => "11101010",22124 => "11101010",22125 => "00111011",22126 => "00111011",22127 => "11000101",22128 => "10001000",22129 => "01100000",22130 => "11101000",22131 => "01001000",22132 => "10010101",22133 => "01001011",22134 => "01100111",22135 => "11001110",22136 => "10100010",22137 => "00101111",22138 => "10000111",22139 => "11001010",22140 => "01100110",22141 => "01100011",22142 => "00110110",22143 => "10110110",22144 => "11010011",22145 => "10110100",22146 => "01101011",22147 => "11100111",22148 => "01111101",22149 => "10011010",22150 => "00010000",22151 => "10111001",22152 => "11011011",22153 => "01000010",22154 => "11111110",22155 => "01001001",22156 => "10111001",22157 => "01001000",22158 => "10110011",22159 => "11000000",22160 => "00101000",22161 => "11011110",22162 => "00101110",22163 => "11101111",22164 => "11001100",22165 => "10100000",22166 => "01011100",22167 => "11111010",22168 => "11000100",22169 => "10111100",22170 => "11101010",22171 => "01001101",22172 => "01000101",22173 => "10110001",22174 => "11010011",22175 => "00100010",22176 => "01011001",22177 => "01000011",22178 => "01110111",22179 => "10000101",22180 => "10010010",22181 => "11101111",22182 => "10110011",22183 => "10001111",22184 => "00001111",22185 => "11111000",22186 => "10110101",22187 => "10101000",22188 => "01011011",22189 => "11111111",22190 => "10011000",22191 => "01111100",22192 => "10011110",22193 => "01000110",22194 => "10011001",22195 => "01101000",22196 => "11000111",22197 => "01001001",22198 => "11000000",22199 => "10011000",22200 => "00101001",22201 => "01110011",22202 => "10000000",22203 => "11000110",22204 => "10011010",22205 => "01110100",22206 => "11110101",22207 => "10011110",22208 => "11000000",22209 => "10101110",22210 => "10110111",22211 => "10111010",22212 => "10110110",22213 => "11111010",22214 => "10001111",22215 => "00100111",22216 => "10010011",22217 => "01110100",22218 => "11011000",22219 => "11101011",22220 => "11111001",22221 => "01000101",22222 => "10101001",22223 => "11010011",22224 => "10111000",22225 => "00000001",22226 => "00110100",22227 => "11111001",22228 => "01010101",22229 => "10100010",22230 => "00010000",22231 => "10100111",22232 => "10001110",22233 => "01011011",22234 => "00101001",22235 => "11101101",22236 => "10110111",22237 => "00100100",22238 => "01001011",22239 => "10101000",22240 => "00000100",22241 => "10100001",22242 => "10101111",22243 => "11111101",22244 => "11111010",22245 => "01001011",22246 => "00101001",22247 => "10001011",22248 => "00110000",22249 => "11011100",22250 => "01011011",22251 => "10111001",22252 => "00000000",22253 => "00111010",22254 => "11101001",22255 => "10010101",22256 => "10101001",22257 => "11010011",22258 => "11110100",22259 => "01101010",22260 => "10111110",22261 => "00101111",22262 => "10001110",22263 => "10000100",22264 => "00101010",22265 => "11000010",22266 => "01111010",22267 => "11000001",22268 => "11111110",22269 => "01000010",22270 => "10110110",22271 => "01011001",22272 => "00000001",22273 => "11101010",22274 => "11010011",22275 => "10000010",22276 => "00001001",22277 => "11110001",22278 => "10110010",22279 => "00101101",22280 => "10110110",22281 => "00100101",22282 => "00100110",22283 => "11010111",22284 => "00101010",22285 => "01111001",22286 => "11100110",22287 => "11101100",22288 => "10010101",22289 => "00101110",22290 => "01000100",22291 => "10100111",22292 => "10011100",22293 => "01000110",22294 => "10110010",22295 => "10100101",22296 => "10110111",22297 => "00000010",22298 => "00010001",22299 => "10110110",22300 => "00010110",22301 => "00111000",22302 => "01011000",22303 => "10111101",22304 => "01000011",22305 => "00011101",22306 => "01101101",22307 => "10001010",22308 => "00000101",22309 => "01100001",22310 => "00100001",22311 => "11010101",22312 => "01100010",22313 => "00010110",22314 => "01011100",22315 => "11000111",22316 => "01111010",22317 => "00100111",22318 => "10100011",22319 => "10001110",22320 => "11110110",22321 => "01000100",22322 => "11100000",22323 => "10010101",22324 => "11000010",22325 => "00001100",22326 => "01111001",22327 => "10111010",22328 => "00000111",22329 => "00010011",22330 => "00111111",22331 => "11000100",22332 => "11110011",22333 => "00110111",22334 => "10010010",22335 => "00011100",22336 => "10011101",22337 => "01001001",22338 => "01111100",22339 => "11001110",22340 => "10100111",22341 => "11110011",22342 => "11101000",22343 => "10010111",22344 => "10111011",22345 => "10100111",22346 => "10110000",22347 => "10001011",22348 => "00010000",22349 => "10111010",22350 => "11000111",22351 => "11001001",22352 => "10100000",22353 => "00111010",22354 => "00101010",22355 => "11001101",22356 => "11110001",22357 => "10000001",22358 => "01000111",22359 => "10111000",22360 => "11111100",22361 => "10001011",22362 => "10110000",22363 => "11001101",22364 => "11010101",22365 => "00110011",22366 => "11100011",22367 => "10010010",22368 => "00110011",22369 => "10111110",22370 => "00011100",22371 => "11001101",22372 => "10110100",22373 => "00010010",22374 => "00011110",22375 => "00100001",22376 => "10100000",22377 => "10110111",22378 => "01111100",22379 => "00011011",22380 => "10110000",22381 => "11010110",22382 => "10001101",22383 => "10010110",22384 => "10100111",22385 => "10001001",22386 => "00111111",22387 => "00101010",22388 => "01101000",22389 => "01111100",22390 => "11110011",22391 => "00110111",22392 => "01100000",22393 => "11000111",22394 => "10111110",22395 => "00101110",22396 => "10001001",22397 => "00111010",22398 => "01001011",22399 => "11011000",22400 => "10110011",22401 => "00010111",22402 => "10110111",22403 => "00101011",22404 => "11100010",22405 => "10101011",22406 => "11110010",22407 => "00011100",22408 => "10111000",22409 => "00101001",22410 => "01010111",22411 => "11011100",22412 => "10101100",22413 => "01000110",22414 => "11101000",22415 => "00000101",22416 => "00011000",22417 => "11111101",22418 => "10111100",22419 => "10001011",22420 => "10000010",22421 => "00010110",22422 => "11010001",22423 => "01100011",22424 => "00001010",22425 => "01111111",22426 => "10000001",22427 => "00100011",22428 => "01100010",22429 => "00110100",22430 => "00100111",22431 => "11010010",22432 => "10010011",22433 => "10011010",22434 => "00011000",22435 => "10010111",22436 => "11110010",22437 => "11100001",22438 => "01001110",22439 => "10110000",22440 => "10000010",22441 => "11111011",22442 => "11001010",22443 => "10101100",22444 => "01010000",22445 => "00110111",22446 => "10110000",22447 => "11100011",22448 => "10000100",22449 => "11101101",22450 => "00110001",22451 => "10110000",22452 => "00110100",22453 => "01111001",22454 => "01000101",22455 => "11110000",22456 => "00101010",22457 => "10100100",22458 => "00010101",22459 => "11010110",22460 => "11111010",22461 => "10111100",22462 => "11000101",22463 => "11000110",22464 => "00011010",22465 => "10000010",22466 => "01101001",22467 => "00111011",22468 => "11001000",22469 => "01101011",22470 => "11000000",22471 => "01011000",22472 => "00000010",22473 => "11011001",22474 => "10111010",22475 => "00001101",22476 => "10100011",22477 => "01000100",22478 => "01000010",22479 => "10100011",22480 => "11100110",22481 => "11000010",22482 => "01001111",22483 => "00000100",22484 => "01101100",22485 => "01111011",22486 => "00001010",22487 => "11110010",22488 => "01010001",22489 => "10000010",22490 => "00111011",22491 => "10010100",22492 => "11111100",22493 => "11101010",22494 => "01101010",22495 => "10111000",22496 => "10001101",22497 => "10010101",22498 => "10010011",22499 => "11001001",22500 => "11110101",22501 => "00100111",22502 => "10000100",22503 => "11110100",22504 => "10001001",22505 => "10111101",22506 => "01010101",22507 => "10001011",22508 => "00100100",22509 => "10011111",22510 => "10011010",22511 => "00100111",22512 => "01110010",22513 => "00011001",22514 => "11000110",22515 => "10100110",22516 => "11110101",22517 => "01110101",22518 => "10111110",22519 => "01101100",22520 => "11110101",22521 => "01101111",22522 => "00011111",22523 => "10111010",22524 => "11101110",22525 => "01010110",22526 => "01101101",22527 => "01111001",22528 => "00011101",22529 => "10001100",22530 => "01110101",22531 => "00000111",22532 => "01000011",22533 => "01100101",22534 => "10010100",22535 => "11111110",22536 => "01100100",22537 => "11111110",22538 => "10101011",22539 => "00110011",22540 => "11101101",22541 => "01111011",22542 => "00000101",22543 => "01101010",22544 => "01000010",22545 => "00000011",22546 => "11000111",22547 => "11111010",22548 => "11101000",22549 => "00111001",22550 => "10100011",22551 => "11101101",22552 => "00001010",22553 => "01110000",22554 => "01011111",22555 => "10111110",22556 => "00000010",22557 => "01000001",22558 => "00111010",22559 => "00110100",22560 => "11000010",22561 => "10110110",22562 => "00011001",22563 => "01101111",22564 => "10010111",22565 => "00100100",22566 => "01011100",22567 => "11011101",22568 => "11111110",22569 => "10011111",22570 => "10100101",22571 => "01110001",22572 => "10001110",22573 => "00101100",22574 => "01001110",22575 => "01000111",22576 => "00001100",22577 => "10100101",22578 => "00010011",22579 => "10001011",22580 => "00010011",22581 => "00000101",22582 => "10101110",22583 => "11100111",22584 => "10010100",22585 => "10000100",22586 => "11000000",22587 => "01001010",22588 => "00011110",22589 => "10011011",22590 => "11011011",22591 => "01001011",22592 => "11001011",22593 => "10000111",22594 => "01011000",22595 => "00010100",22596 => "01110101",22597 => "00010011",22598 => "10100001",22599 => "00101101",22600 => "11001111",22601 => "11011111",22602 => "00111000",22603 => "11101100",22604 => "11101100",22605 => "00111100",22606 => "10110110",22607 => "10101000",22608 => "11101011",22609 => "10000011",22610 => "00100100",22611 => "01001010",22612 => "10100000",22613 => "01011011",22614 => "00110010",22615 => "11001010",22616 => "00000100",22617 => "11011001",22618 => "00111101",22619 => "10010111",22620 => "10110101",22621 => "01011110",22622 => "10011001",22623 => "11001011",22624 => "00010100",22625 => "10011010",22626 => "01111100",22627 => "01000111",22628 => "10011101",22629 => "11001001",22630 => "01100101",22631 => "10100110",22632 => "00110100",22633 => "11111100",22634 => "00001011",22635 => "11100111",22636 => "10101100",22637 => "10001010",22638 => "01101111",22639 => "11011010",22640 => "01010010",22641 => "10001010",22642 => "01111000",22643 => "11001101",22644 => "11110000",22645 => "10001100",22646 => "01111111",22647 => "10010110",22648 => "00111110",22649 => "01000011",22650 => "00000010",22651 => "00001000",22652 => "00101000",22653 => "11111100",22654 => "01000011",22655 => "10101101",22656 => "01010001",22657 => "00001100",22658 => "10101000",22659 => "01101001",22660 => "00010001",22661 => "00111110",22662 => "01101110",22663 => "01010000",22664 => "11011000",22665 => "10101011",22666 => "01100110",22667 => "00111111",22668 => "10001101",22669 => "00101011",22670 => "01111111",22671 => "01111110",22672 => "10011110",22673 => "01000010",22674 => "11110100",22675 => "01001111",22676 => "11011010",22677 => "10100111",22678 => "10101000",22679 => "10110110",22680 => "10001100",22681 => "10001001",22682 => "00111010",22683 => "10111100",22684 => "11101000",22685 => "11001110",22686 => "01101011",22687 => "10001010",22688 => "10100111",22689 => "10110101",22690 => "00101000",22691 => "11101110",22692 => "11010101",22693 => "00100110",22694 => "10011100",22695 => "11110001",22696 => "00100011",22697 => "01111000",22698 => "10000101",22699 => "00111011",22700 => "01011001",22701 => "01110111",22702 => "10110111",22703 => "00011000",22704 => "01001010",22705 => "11111001",22706 => "11001100",22707 => "00001001",22708 => "11100100",22709 => "10011111",22710 => "01111010",22711 => "01110111",22712 => "10000001",22713 => "11011110",22714 => "10010011",22715 => "01111110",22716 => "11110000",22717 => "00110110",22718 => "10011001",22719 => "00010010",22720 => "11100101",22721 => "00001001",22722 => "01001001",22723 => "00111011",22724 => "00101100",22725 => "00000001",22726 => "01111110",22727 => "01000011",22728 => "11100000",22729 => "11001000",22730 => "01001010",22731 => "10100011",22732 => "10111000",22733 => "11000100",22734 => "10000111",22735 => "10110111",22736 => "00111101",22737 => "00010000",22738 => "10101100",22739 => "10001010",22740 => "01101011",22741 => "10111010",22742 => "10001010",22743 => "01100111",22744 => "11110100",22745 => "11111111",22746 => "11011000",22747 => "01110010",22748 => "01100101",22749 => "00110000",22750 => "00000101",22751 => "11110001",22752 => "01011000",22753 => "00111110",22754 => "10001101",22755 => "10001111",22756 => "01001100",22757 => "11111010",22758 => "10010100",22759 => "01001100",22760 => "00001011",22761 => "10101011",22762 => "11100111",22763 => "01101011",22764 => "10000010",22765 => "00101100",22766 => "10011100",22767 => "11010110",22768 => "00000111",22769 => "10100001",22770 => "01111010",22771 => "11010011",22772 => "00000110",22773 => "01110100",22774 => "00010100",22775 => "01101000",22776 => "10011000",22777 => "10101011",22778 => "11111110",22779 => "01101011",22780 => "11100100",22781 => "01001011",22782 => "01111011",22783 => "11011001",22784 => "11000000",22785 => "11100000",22786 => "11001001",22787 => "10010100",22788 => "10110111",22789 => "10111111",22790 => "01100111",22791 => "00101110",22792 => "00101000",22793 => "01111111",22794 => "10011111",22795 => "11101110",22796 => "01010101",22797 => "00010000",22798 => "11001001",22799 => "00100001",22800 => "10100101",22801 => "10010100",22802 => "01100110",22803 => "11010010",22804 => "00000000",22805 => "11011011",22806 => "11010011",22807 => "11100100",22808 => "01100110",22809 => "10000110",22810 => "00100011",22811 => "10111110",22812 => "11001010",22813 => "11011010",22814 => "10100011",22815 => "00101110",22816 => "10101111",22817 => "10011111",22818 => "11010111",22819 => "11000110",22820 => "01001000",22821 => "00111010",22822 => "10011101",22823 => "00010001",22824 => "00001110",22825 => "10101011",22826 => "10100110",22827 => "10101100",22828 => "00110010",22829 => "00011110",22830 => "10000011",22831 => "00110100",22832 => "01010011",22833 => "11001011",22834 => "10100000",22835 => "11100100",22836 => "10011001",22837 => "11011101",22838 => "10101011",22839 => "11001101",22840 => "00110100",22841 => "10000100",22842 => "10101101",22843 => "01100011",22844 => "10110001",22845 => "11110100",22846 => "11011100",22847 => "10001100",22848 => "00100101",22849 => "00100100",22850 => "00111000",22851 => "11100100",22852 => "01010110",22853 => "00100111",22854 => "01101101",22855 => "01101001",22856 => "01010111",22857 => "10010100",22858 => "10000001",22859 => "11011111",22860 => "00001101",22861 => "11111001",22862 => "11111101",22863 => "10101111",22864 => "00011110",22865 => "10001111",22866 => "10010111",22867 => "01110101",22868 => "00000111",22869 => "11000011",22870 => "10010011",22871 => "11110010",22872 => "01111110",22873 => "10100110",22874 => "01111101",22875 => "00110100",22876 => "11000001",22877 => "01111010",22878 => "11110000",22879 => "00100001",22880 => "00111110",22881 => "10001111",22882 => "10110011",22883 => "01010011",22884 => "11100110",22885 => "10110011",22886 => "11111011",22887 => "11111000",22888 => "11010011",22889 => "00011010",22890 => "10011111",22891 => "00111000",22892 => "00011010",22893 => "01111010",22894 => "10111101",22895 => "11001001",22896 => "01110011",22897 => "11011011",22898 => "11000100",22899 => "11100011",22900 => "11010111",22901 => "01110010",22902 => "00001011",22903 => "01010111",22904 => "00000110",22905 => "11000010",22906 => "11101111",22907 => "11101100",22908 => "10000011",22909 => "10001001",22910 => "01000110",22911 => "11101101",22912 => "11100010",22913 => "00010000",22914 => "10010010",22915 => "11000101",22916 => "11010110",22917 => "10011011",22918 => "01100001",22919 => "10110110",22920 => "10011111",22921 => "11001010",22922 => "10010010",22923 => "00111110",22924 => "10100010",22925 => "01110000",22926 => "10011011",22927 => "11100010",22928 => "00100110",22929 => "01011101",22930 => "10000011",22931 => "00010100",22932 => "01111111",22933 => "10010110",22934 => "11011110",22935 => "00101011",22936 => "11111100",22937 => "01011011",22938 => "01011000",22939 => "00110000",22940 => "10001010",22941 => "01000111",22942 => "10011100",22943 => "10010010",22944 => "11010000",22945 => "00111100",22946 => "01111111",22947 => "00011101",22948 => "10011011",22949 => "00111001",22950 => "01111001",22951 => "00100001",22952 => "00001101",22953 => "00001110",22954 => "01101011",22955 => "01100010",22956 => "00000111",22957 => "00010001",22958 => "10010001",22959 => "01111100",22960 => "01011100",22961 => "11000010",22962 => "10110011",22963 => "01001100",22964 => "01110100",22965 => "11111000",22966 => "01001110",22967 => "10110001",22968 => "11110110",22969 => "10110011",22970 => "11111100",22971 => "10010011",22972 => "01110111",22973 => "11001111",22974 => "11011110",22975 => "01110101",22976 => "10000110",22977 => "11000100",22978 => "00110000",22979 => "11111011",22980 => "11011010",22981 => "11000000",22982 => "10001101",22983 => "10011000",22984 => "00001101",22985 => "11011100",22986 => "10010101",22987 => "00111100",22988 => "11100001",22989 => "01100110",22990 => "00010000",22991 => "00110110",22992 => "01010110",22993 => "11101001",22994 => "11111000",22995 => "10000110",22996 => "11010111",22997 => "11110010",22998 => "10000011",22999 => "01011101",23000 => "10110010",23001 => "01110101",23002 => "10110000",23003 => "11001011",23004 => "00010000",23005 => "00101011",23006 => "01111000",23007 => "10111111",23008 => "11011110",23009 => "11000011",23010 => "11111101",23011 => "11011011",23012 => "01011101",23013 => "11100001",23014 => "10011000",23015 => "00111111",23016 => "01100111",23017 => "01011110",23018 => "01100001",23019 => "01100101",23020 => "01100111",23021 => "00011001",23022 => "11011000",23023 => "10010110",23024 => "01101110",23025 => "00111111",23026 => "10100111",23027 => "01001101",23028 => "00011001",23029 => "00000001",23030 => "11001110",23031 => "11001111",23032 => "01101010",23033 => "01101111",23034 => "11011000",23035 => "11110111",23036 => "00101000",23037 => "01000110",23038 => "01000011",23039 => "01110111",23040 => "10000011",23041 => "00111010",23042 => "11000010",23043 => "01010001",23044 => "00000011",23045 => "11011111",23046 => "00110100",23047 => "11010001",23048 => "10011001",23049 => "10100100",23050 => "11011001",23051 => "01011000",23052 => "00011010",23053 => "01111100",23054 => "11111001",23055 => "00011110",23056 => "01001100",23057 => "00101010",23058 => "10101000",23059 => "10011110",23060 => "01011001",23061 => "00000100",23062 => "11000000",23063 => "11110000",23064 => "00101010",23065 => "11100101",23066 => "00100101",23067 => "00000100",23068 => "01001001",23069 => "11101000",23070 => "10100101",23071 => "11011011",23072 => "11000111",23073 => "00110101",23074 => "00000000",23075 => "01001000",23076 => "11110110",23077 => "01111101",23078 => "00111010",23079 => "00110110",23080 => "10000100",23081 => "10000100",23082 => "11100110",23083 => "01000101",23084 => "11100000",23085 => "11010011",23086 => "10011011",23087 => "00100101",23088 => "01111101",23089 => "10000110",23090 => "01100001",23091 => "00011010",23092 => "10011011",23093 => "10001110",23094 => "00000111",23095 => "11100000",23096 => "00000101",23097 => "10010100",23098 => "00000111",23099 => "11011010",23100 => "11111000",23101 => "11110000",23102 => "01111100",23103 => "00110001",23104 => "11101101",23105 => "11100010",23106 => "10111001",23107 => "01111100",23108 => "01111101",23109 => "10011000",23110 => "11110001",23111 => "01100100",23112 => "11001010",23113 => "01110010",23114 => "01011101",23115 => "00010001",23116 => "11001100",23117 => "11100001",23118 => "01111001",23119 => "01000011",23120 => "11101010",23121 => "11111011",23122 => "00100101",23123 => "01001010",23124 => "00000001",23125 => "11001001",23126 => "11110100",23127 => "00000010",23128 => "00110101",23129 => "10110101",23130 => "00101000",23131 => "11110110",23132 => "00010000",23133 => "00000001",23134 => "11110111",23135 => "11100110",23136 => "11001000",23137 => "10000011",23138 => "11011000",23139 => "10000000",23140 => "10101001",23141 => "11101011",23142 => "00101011",23143 => "11111000",23144 => "01101110",23145 => "10011111",23146 => "00001011",23147 => "10110110",23148 => "11011101",23149 => "10100101",23150 => "01001111",23151 => "01011110",23152 => "11010001",23153 => "11011111",23154 => "10101001",23155 => "11010111",23156 => "01111100",23157 => "01000000",23158 => "01111000",23159 => "00101011",23160 => "00000011",23161 => "11011001",23162 => "01011100",23163 => "10001101",23164 => "10000010",23165 => "01100111",23166 => "01001010",23167 => "10110011",23168 => "10100111",23169 => "01101101",23170 => "11011100",23171 => "00000100",23172 => "01010110",23173 => "00110100",23174 => "10001111",23175 => "01011101",23176 => "11010000",23177 => "11011001",23178 => "11100011",23179 => "10011000",23180 => "01111011",23181 => "11010111",23182 => "11010100",23183 => "01101001",23184 => "01000100",23185 => "10000010",23186 => "11011010",23187 => "00010001",23188 => "01000101",23189 => "11001100",23190 => "01111101",23191 => "01000101",23192 => "00011010",23193 => "10100011",23194 => "00111101",23195 => "00110100",23196 => "11011001",23197 => "10101100",23198 => "10110000",23199 => "01010100",23200 => "00100011",23201 => "01101110",23202 => "11110001",23203 => "00000000",23204 => "00100000",23205 => "01001001",23206 => "11111011",23207 => "11101110",23208 => "10000110",23209 => "10010110",23210 => "01011110",23211 => "01010000",23212 => "01111000",23213 => "11111110",23214 => "00110110",23215 => "10110001",23216 => "00101111",23217 => "11010000",23218 => "11011011",23219 => "01010010",23220 => "11011011",23221 => "10010100",23222 => "01011010",23223 => "11010111",23224 => "10000010",23225 => "11011110",23226 => "01011110",23227 => "11001101",23228 => "00111011",23229 => "11110000",23230 => "00100000",23231 => "10100011",23232 => "00000110",23233 => "10100111",23234 => "10011011",23235 => "11010001",23236 => "01001011",23237 => "10100010",23238 => "00101011",23239 => "11011110",23240 => "11001110",23241 => "00011000",23242 => "11110001",23243 => "11011100",23244 => "01110001",23245 => "11110101",23246 => "11001111",23247 => "11000101",23248 => "01011110",23249 => "10000101",23250 => "11000001",23251 => "00000111",23252 => "10111100",23253 => "10001110",23254 => "11110101",23255 => "10100001",23256 => "11000100",23257 => "01100011",23258 => "01001010",23259 => "11101111",23260 => "00110111",23261 => "01010010",23262 => "01000110",23263 => "00000100",23264 => "00010011",23265 => "11001011",23266 => "10110001",23267 => "00010010",23268 => "01111011",23269 => "00101110",23270 => "01001111",23271 => "10100001",23272 => "11001111",23273 => "10110010",23274 => "11111100",23275 => "11011101",23276 => "10100011",23277 => "00000110",23278 => "01101111",23279 => "01010011",23280 => "00010010",23281 => "00101000",23282 => "10111011",23283 => "00111011",23284 => "00110111",23285 => "10100000",23286 => "11010011",23287 => "10000011",23288 => "10111111",23289 => "01011010",23290 => "10100111",23291 => "00101011",23292 => "00110011",23293 => "10100100",23294 => "10111101",23295 => "10111101",23296 => "01000011",23297 => "00011001",23298 => "00000000",23299 => "11011000",23300 => "01000110",23301 => "10111011",23302 => "00111100",23303 => "01010010",23304 => "00010101",23305 => "10000011",23306 => "10011011",23307 => "00000011",23308 => "01100010",23309 => "01011000",23310 => "01111010",23311 => "11101011",23312 => "10111111",23313 => "01100010",23314 => "01001011",23315 => "01101101",23316 => "01111100",23317 => "00101110",23318 => "10010110",23319 => "10000111",23320 => "11010101",23321 => "11010001",23322 => "11011101",23323 => "10100111",23324 => "10000100",23325 => "11110110",23326 => "10110110",23327 => "00111111",23328 => "00010101",23329 => "00011101",23330 => "00111110",23331 => "01011011",23332 => "00100010",23333 => "00111001",23334 => "10110111",23335 => "01000001",23336 => "01001000",23337 => "10100011",23338 => "11111101",23339 => "01100110",23340 => "11100010",23341 => "00101100",23342 => "10110111",23343 => "01111101",23344 => "11001000",23345 => "11001011",23346 => "00111001",23347 => "00001110",23348 => "11000011",23349 => "01011100",23350 => "00000011",23351 => "01000000",23352 => "10110111",23353 => "11110111",23354 => "00111111",23355 => "00101100",23356 => "01010110",23357 => "00111010",23358 => "10100100",23359 => "01011100",23360 => "01011000",23361 => "01100000",23362 => "00100111",23363 => "01100100",23364 => "00000010",23365 => "10010010",23366 => "00111111",23367 => "01101101",23368 => "10011110",23369 => "11001001",23370 => "10100101",23371 => "11110111",23372 => "00111000",23373 => "00100011",23374 => "00010101",23375 => "11000100",23376 => "10111010",23377 => "01001000",23378 => "00111101",23379 => "00000101",23380 => "11111100",23381 => "11000110",23382 => "00101110",23383 => "01100011",23384 => "10000100",23385 => "11011110",23386 => "00100001",23387 => "10110111",23388 => "10111011",23389 => "00100101",23390 => "11110110",23391 => "01111000",23392 => "10111011",23393 => "11001100",23394 => "00101010",23395 => "00101000",23396 => "10001011",23397 => "01000101",23398 => "10001001",23399 => "01100010",23400 => "00100011",23401 => "11101011",23402 => "10100110",23403 => "00001101",23404 => "11100000",23405 => "11111101",23406 => "00110100",23407 => "01110011",23408 => "00010001",23409 => "11011110",23410 => "11111000",23411 => "00010111",23412 => "10000010",23413 => "10001110",23414 => "10011101",23415 => "10100101",23416 => "10100001",23417 => "00111101",23418 => "01011101",23419 => "10010001",23420 => "01100001",23421 => "10101110",23422 => "01000110",23423 => "11101110",23424 => "00011101",23425 => "01101011",23426 => "00110010",23427 => "10101011",23428 => "11110100",23429 => "10110110",23430 => "10101010",23431 => "00101000",23432 => "11001100",23433 => "01011001",23434 => "01100011",23435 => "10111111",23436 => "01001101",23437 => "11111100",23438 => "00110010",23439 => "11101111",23440 => "11010000",23441 => "00000011",23442 => "01001100",23443 => "11001001",23444 => "10000101",23445 => "01111000",23446 => "00010110",23447 => "10001000",23448 => "11111011",23449 => "10101001",23450 => "01101100",23451 => "00110100",23452 => "00100101",23453 => "10001101",23454 => "00011000",23455 => "00011101",23456 => "10110010",23457 => "11001111",23458 => "11100001",23459 => "01010001",23460 => "10010110",23461 => "00111110",23462 => "00111000",23463 => "11111110",23464 => "00000101",23465 => "01000011",23466 => "11100100",23467 => "01100011",23468 => "10010011",23469 => "11111010",23470 => "11111110",23471 => "11010101",23472 => "11000000",23473 => "11010111",23474 => "10011001",23475 => "11111001",23476 => "01000101",23477 => "00000101",23478 => "01001000",23479 => "10001101",23480 => "11000011",23481 => "11000001",23482 => "10111010",23483 => "10011000",23484 => "11100001",23485 => "11011111",23486 => "11011011",23487 => "01111101",23488 => "00001000",23489 => "11011000",23490 => "01110010",23491 => "01010111",23492 => "10101010",23493 => "10011011",23494 => "01111001",23495 => "11010001",23496 => "00011101",23497 => "01010101",23498 => "11111001",23499 => "01100010",23500 => "10101000",23501 => "01110001",23502 => "11110000",23503 => "10010100",23504 => "00010001",23505 => "11111101",23506 => "01011001",23507 => "01101011",23508 => "00110000",23509 => "01111000",23510 => "11001110",23511 => "11001000",23512 => "11010111",23513 => "11100011",23514 => "11111100",23515 => "01111010",23516 => "01010101",23517 => "01001101",23518 => "00100000",23519 => "10011001",23520 => "01100100",23521 => "11010000",23522 => "11001011",23523 => "01111000",23524 => "11111000",23525 => "01001110",23526 => "10001100",23527 => "11011110",23528 => "01111010",23529 => "01000000",23530 => "00101101",23531 => "10111110",23532 => "01000100",23533 => "00001010",23534 => "00100000",23535 => "00010010",23536 => "00111111",23537 => "10000011",23538 => "10110110",23539 => "11010111",23540 => "00111100",23541 => "10110110",23542 => "10000010",23543 => "00100000",23544 => "01100011",23545 => "00001101",23546 => "10011100",23547 => "10010111",23548 => "10110001",23549 => "01110010",23550 => "10110001",23551 => "01100001",23552 => "10000111",23553 => "11110100",23554 => "11110010",23555 => "10110110",23556 => "00010011",23557 => "00001011",23558 => "10100001",23559 => "00000001",23560 => "10110010",23561 => "01100011",23562 => "11111000",23563 => "01100000",23564 => "11101110",23565 => "00110100",23566 => "10100010",23567 => "11000011",23568 => "01001000",23569 => "11111110",23570 => "00001110",23571 => "10000001",23572 => "10111100",23573 => "01110110",23574 => "01111101",23575 => "10001101",23576 => "01110101",23577 => "01010010",23578 => "00001101",23579 => "10101001",23580 => "10101000",23581 => "00110100",23582 => "00011000",23583 => "01111010",23584 => "01101100",23585 => "11000100",23586 => "10000001",23587 => "11010100",23588 => "11101110",23589 => "11011010",23590 => "01111000",23591 => "01011101",23592 => "00001011",23593 => "00010001",23594 => "01100110",23595 => "01101001",23596 => "00100000",23597 => "01000101",23598 => "10101100",23599 => "10011000",23600 => "11000100",23601 => "11010000",23602 => "00010011",23603 => "01111100",23604 => "11000001",23605 => "01100100",23606 => "11011110",23607 => "10110001",23608 => "00011101",23609 => "01010100",23610 => "10010111",23611 => "10011100",23612 => "10001001",23613 => "01010010",23614 => "01010001",23615 => "11000011",23616 => "01110000",23617 => "11000011",23618 => "10000011",23619 => "00100100",23620 => "11111100",23621 => "01010111",23622 => "01100011",23623 => "01100000",23624 => "11001011",23625 => "10010000",23626 => "10001011",23627 => "11101001",23628 => "10011000",23629 => "00100101",23630 => "11111110",23631 => "00100011",23632 => "00101011",23633 => "10110010",23634 => "01101110",23635 => "01100110",23636 => "01011111",23637 => "11010001",23638 => "01101110",23639 => "11010101",23640 => "10010010",23641 => "01010101",23642 => "10100011",23643 => "01000000",23644 => "11110111",23645 => "11010101",23646 => "11000101",23647 => "01010001",23648 => "01110110",23649 => "10011110",23650 => "11001110",23651 => "01010100",23652 => "01001010",23653 => "00000001",23654 => "11001110",23655 => "00001000",23656 => "01100111",23657 => "00100101",23658 => "00011011",23659 => "11000000",23660 => "10001110",23661 => "10111001",23662 => "10110110",23663 => "11100111",23664 => "01000000",23665 => "00000110",23666 => "01100101",23667 => "10110011",23668 => "00111110",23669 => "11111001",23670 => "10011010",23671 => "00110111",23672 => "11000101",23673 => "10101001",23674 => "11001011",23675 => "11100011",23676 => "10110000",23677 => "11111011",23678 => "11101011",23679 => "01100110",23680 => "01000001",23681 => "11111010",23682 => "11101110",23683 => "11100001",23684 => "11101000",23685 => "10001110",23686 => "01110100",23687 => "01101100",23688 => "01000100",23689 => "10101011",23690 => "11010000",23691 => "00000100",23692 => "11110011",23693 => "10010100",23694 => "01100000",23695 => "01101010",23696 => "11110101",23697 => "10011111",23698 => "10001011",23699 => "01011101",23700 => "01011001",23701 => "10001011",23702 => "11101101",23703 => "00110001",23704 => "00010001",23705 => "00110001",23706 => "01110110",23707 => "01000011",23708 => "00010100",23709 => "00011111",23710 => "11100011",23711 => "01111100",23712 => "01101101",23713 => "00011101",23714 => "00111100",23715 => "10011110",23716 => "11100010",23717 => "10100001",23718 => "11000111",23719 => "10111011",23720 => "11000111",23721 => "11111110",23722 => "01110000",23723 => "10001001",23724 => "10010010",23725 => "10111100",23726 => "00010000",23727 => "10011111",23728 => "01000010",23729 => "00011111",23730 => "10001000",23731 => "11111001",23732 => "01000001",23733 => "11001010",23734 => "00101101",23735 => "11100011",23736 => "00011010",23737 => "11010010",23738 => "00110100",23739 => "10101011",23740 => "00010110",23741 => "11010111",23742 => "00101110",23743 => "11111101",23744 => "00111100",23745 => "01000101",23746 => "00100001",23747 => "00000101",23748 => "00010011",23749 => "11011011",23750 => "00011001",23751 => "10100111",23752 => "00110010",23753 => "11101001",23754 => "10001011",23755 => "01101101",23756 => "01000000",23757 => "00110100",23758 => "00101101",23759 => "10010100",23760 => "11100010",23761 => "01011000",23762 => "11000111",23763 => "01110100",23764 => "11001010",23765 => "10100110",23766 => "11100101",23767 => "01101101",23768 => "01110001",23769 => "01001011",23770 => "01101010",23771 => "11100000",23772 => "01111000",23773 => "11110011",23774 => "00101001",23775 => "01101111",23776 => "01101010",23777 => "10000000",23778 => "01011100",23779 => "10011001",23780 => "01011011",23781 => "00010100",23782 => "01101101",23783 => "11101110",23784 => "10011000",23785 => "00011110",23786 => "00110001",23787 => "00010001",23788 => "11110011",23789 => "11101100",23790 => "10001001",23791 => "00101010",23792 => "01110111",23793 => "01111011",23794 => "10010001",23795 => "10010011",23796 => "10010110",23797 => "01111011",23798 => "01111011",23799 => "01101000",23800 => "00011100",23801 => "11110111",23802 => "11001010",23803 => "01111010",23804 => "00001010",23805 => "00111110",23806 => "10010011",23807 => "01000100",23808 => "01101110",23809 => "00100001",23810 => "01000111",23811 => "10000001",23812 => "11011011",23813 => "11001001",23814 => "10011010",23815 => "00101110",23816 => "11110000",23817 => "10110010",23818 => "11100110",23819 => "01100111",23820 => "10011000",23821 => "11100011",23822 => "00100001",23823 => "11011100",23824 => "10010010",23825 => "11111110",23826 => "11110111",23827 => "10000001",23828 => "01001110",23829 => "10011101",23830 => "00001001",23831 => "01000001",23832 => "11000011",23833 => "00010111",23834 => "10111011",23835 => "00001011",23836 => "00001001",23837 => "10110011",23838 => "00001111",23839 => "10111001",23840 => "10001101",23841 => "00010110",23842 => "01000010",23843 => "01100100",23844 => "01000111",23845 => "01110001",23846 => "10110110",23847 => "11101010",23848 => "10110001",23849 => "10011001",23850 => "10011010",23851 => "10111100",23852 => "10100100",23853 => "11010000",23854 => "11010100",23855 => "00100100",23856 => "10000111",23857 => "10101101",23858 => "10100100",23859 => "00001111",23860 => "10111101",23861 => "00110000",23862 => "10110110",23863 => "10001010",23864 => "00001011",23865 => "10101101",23866 => "10001011",23867 => "11110001",23868 => "00010110",23869 => "00000111",23870 => "00111111",23871 => "11110001",23872 => "10010100",23873 => "01000011",23874 => "01000000",23875 => "10011110",23876 => "01010110",23877 => "00000100",23878 => "01000000",23879 => "10001000",23880 => "01111011",23881 => "01010111",23882 => "10111110",23883 => "01111000",23884 => "10000011",23885 => "01111101",23886 => "00101101",23887 => "00011100",23888 => "00011011",23889 => "10110001",23890 => "11110000",23891 => "01110001",23892 => "10101110",23893 => "10101010",23894 => "10001111",23895 => "11010111",23896 => "11110010",23897 => "10010010",23898 => "01011101",23899 => "10100001",23900 => "00101010",23901 => "00010000",23902 => "01101001",23903 => "11001000",23904 => "10111010",23905 => "01111001",23906 => "01001100",23907 => "00011010",23908 => "10010000",23909 => "00001101",23910 => "01100101",23911 => "00100110",23912 => "10011111",23913 => "10100010",23914 => "10011111",23915 => "01100000",23916 => "10101011",23917 => "01011101",23918 => "00000010",23919 => "10111111",23920 => "00110001",23921 => "11001100",23922 => "01001010",23923 => "00010000",23924 => "00101101",23925 => "01110010",23926 => "01000011",23927 => "11101110",23928 => "00100111",23929 => "00010000",23930 => "01111011",23931 => "10100010",23932 => "11111101",23933 => "11111111",23934 => "10000011",23935 => "10000101",23936 => "11101000",23937 => "01110110",23938 => "10110001",23939 => "10000001",23940 => "10001110",23941 => "10100011",23942 => "01000111",23943 => "00110000",23944 => "00010001",23945 => "00100100",23946 => "10110010",23947 => "01111110",23948 => "01000110",23949 => "10111100",23950 => "00001001",23951 => "01010001",23952 => "11011111",23953 => "01001111",23954 => "00011010",23955 => "11101101",23956 => "01011110",23957 => "00100000",23958 => "10011110",23959 => "00000111",23960 => "00101111",23961 => "10111111",23962 => "00010000",23963 => "00001110",23964 => "11101111",23965 => "10000010",23966 => "11111011",23967 => "00011001",23968 => "11011011",23969 => "00011000",23970 => "01011001",23971 => "00000111",23972 => "10101100",23973 => "00100001",23974 => "11100110",23975 => "01101011",23976 => "10010011",23977 => "01110101",23978 => "00100111",23979 => "01011010",23980 => "10011000",23981 => "00001110",23982 => "10001010",23983 => "01100110",23984 => "00101100",23985 => "10001101",23986 => "00111110",23987 => "11000010",23988 => "00010101",23989 => "00011001",23990 => "10110000",23991 => "10001000",23992 => "00010101",23993 => "11010010",23994 => "01001000",23995 => "00111000",23996 => "10000011",23997 => "11001110",23998 => "10010101",23999 => "11100100",24000 => "00100011",24001 => "01101101",24002 => "11100001",24003 => "01101110",24004 => "01000111",24005 => "01010011",24006 => "11000010",24007 => "01110110",24008 => "10100101",24009 => "01101100",24010 => "01011010",24011 => "11010010",24012 => "01111110",24013 => "10011000",24014 => "11101010",24015 => "10011011",24016 => "11101101",24017 => "01111111",24018 => "01101000",24019 => "10000010",24020 => "00001001",24021 => "00000110",24022 => "11000100",24023 => "11011110",24024 => "01010001",24025 => "11111101",24026 => "10101001",24027 => "00010011",24028 => "10110001",24029 => "10101011",24030 => "10110100",24031 => "11011011",24032 => "11011000",24033 => "01101110",24034 => "01000001",24035 => "00101111",24036 => "01010100",24037 => "10110111",24038 => "10001100",24039 => "10010011",24040 => "01101101",24041 => "01110100",24042 => "00011001",24043 => "11001110",24044 => "10000010",24045 => "00010100",24046 => "01100011",24047 => "01000101",24048 => "00010101",24049 => "11011101",24050 => "00010110",24051 => "11001110",24052 => "01101100",24053 => "00110111",24054 => "01101001",24055 => "11100011",24056 => "11011001",24057 => "10011110",24058 => "10010101",24059 => "00110101",24060 => "00000110",24061 => "00000111",24062 => "01110000",24063 => "01011110",24064 => "00100110",24065 => "01110100",24066 => "10001100",24067 => "01111111",24068 => "11001000",24069 => "00001001",24070 => "11010100",24071 => "01010001",24072 => "11000101",24073 => "11111011",24074 => "00001110",24075 => "11110001",24076 => "10000001",24077 => "11001011",24078 => "00110110",24079 => "00000100",24080 => "11011000",24081 => "10010100",24082 => "00111011",24083 => "01001100",24084 => "00110011",24085 => "01101110",24086 => "10100111",24087 => "01000001",24088 => "11110110",24089 => "10001001",24090 => "10000011",24091 => "00111100",24092 => "11110010",24093 => "10101001",24094 => "00011100",24095 => "01100110",24096 => "11100110",24097 => "01100001",24098 => "10001010",24099 => "11111100",24100 => "00001001",24101 => "00101010",24102 => "11100111",24103 => "11110011",24104 => "10110101",24105 => "11110011",24106 => "00001110",24107 => "01011001",24108 => "00001110",24109 => "10100011",24110 => "00101100",24111 => "10000001",24112 => "11100001",24113 => "11111100",24114 => "10001101",24115 => "10001100",24116 => "00010101",24117 => "11111011",24118 => "01010001",24119 => "00011000",24120 => "11010000",24121 => "11000111",24122 => "01000000",24123 => "00010000",24124 => "00101101",24125 => "11001011",24126 => "01101010",24127 => "00001000",24128 => "11111001",24129 => "10101011",24130 => "00111011",24131 => "10101100",24132 => "00000100",24133 => "00000010",24134 => "11000001",24135 => "11101001",24136 => "01101010",24137 => "10000101",24138 => "01001011",24139 => "11100010",24140 => "11001100",24141 => "11011100",24142 => "01001110",24143 => "10110101",24144 => "01001010",24145 => "11110001",24146 => "01000000",24147 => "00000101",24148 => "01110100",24149 => "00111011",24150 => "10110011",24151 => "10101001",24152 => "00001011",24153 => "00001111",24154 => "11101101",24155 => "00101111",24156 => "01000010",24157 => "11110101",24158 => "01110101",24159 => "01001111",24160 => "01101111",24161 => "11110011",24162 => "11110011",24163 => "11010110",24164 => "11010110",24165 => "00111100",24166 => "01011100",24167 => "01100011",24168 => "01011011",24169 => "01101100",24170 => "00101111",24171 => "11100010",24172 => "00100101",24173 => "01101001",24174 => "11101111",24175 => "11010111",24176 => "11100110",24177 => "00000011",24178 => "11101100",24179 => "11110111",24180 => "10110100",24181 => "10111001",24182 => "11110011",24183 => "01000001",24184 => "11110111",24185 => "00100111",24186 => "01101000",24187 => "10101000",24188 => "10110110",24189 => "11111101",24190 => "01001101",24191 => "11100101",24192 => "11010000",24193 => "01100001",24194 => "00010011",24195 => "00001110",24196 => "00000001",24197 => "00011001",24198 => "01111011",24199 => "10000011",24200 => "10100111",24201 => "10011101",24202 => "10100101",24203 => "00101100",24204 => "00111110",24205 => "10000110",24206 => "00001001",24207 => "10100101",24208 => "11111011",24209 => "11110101",24210 => "00001101",24211 => "01001100",24212 => "10011000",24213 => "01011001",24214 => "01110100",24215 => "10001010",24216 => "00001100",24217 => "10011100",24218 => "00110110",24219 => "00110111",24220 => "11011011",24221 => "00011110",24222 => "11011011",24223 => "01111110",24224 => "11100111",24225 => "11100111",24226 => "11110011",24227 => "11110100",24228 => "10010100",24229 => "01001001",24230 => "11110110",24231 => "01011111",24232 => "11010101",24233 => "00001100",24234 => "00010011",24235 => "01111000",24236 => "00011111",24237 => "00000100",24238 => "10111111",24239 => "11111100",24240 => "00111100",24241 => "01100110",24242 => "11111000",24243 => "10011110",24244 => "10101010",24245 => "10011010",24246 => "11011101",24247 => "01001010",24248 => "00011100",24249 => "10101010",24250 => "10000101",24251 => "11101000",24252 => "10101100",24253 => "10011110",24254 => "01111101",24255 => "01000000",24256 => "01001101",24257 => "10011001",24258 => "01101110",24259 => "10010011",24260 => "00101000",24261 => "00000010",24262 => "01000110",24263 => "10111011",24264 => "01000110",24265 => "10001111",24266 => "00011001",24267 => "00111011",24268 => "01110000",24269 => "10111010",24270 => "00000101",24271 => "00110001",24272 => "11001001",24273 => "10010000",24274 => "00110100",24275 => "00001010",24276 => "00001111",24277 => "10011101",24278 => "11000011",24279 => "11100000",24280 => "11010010",24281 => "00110000",24282 => "10101010",24283 => "10101101",24284 => "00010110",24285 => "00010111",24286 => "00010000",24287 => "00110110",24288 => "10000010",24289 => "10001111",24290 => "10010101",24291 => "01100101",24292 => "11000100",24293 => "01101100",24294 => "10110010",24295 => "00001111",24296 => "11101010",24297 => "01011001",24298 => "10100011",24299 => "00110100",24300 => "11110010",24301 => "11011110",24302 => "00010110",24303 => "00011011",24304 => "10010010",24305 => "01011101",24306 => "01011010",24307 => "10100010",24308 => "10011101",24309 => "10110101",24310 => "11000000",24311 => "01101011",24312 => "00101001",24313 => "10111101",24314 => "10101001",24315 => "10000011",24316 => "10000010",24317 => "01011001",24318 => "11110110",24319 => "10111111",24320 => "01000000",24321 => "01000100",24322 => "11010110",24323 => "01010000",24324 => "00110110",24325 => "10000111",24326 => "10110100",24327 => "10000001",24328 => "01111000",24329 => "10011010",24330 => "11101110",24331 => "00001000",24332 => "11110000",24333 => "11110110",24334 => "00010001",24335 => "11110101",24336 => "11110100",24337 => "01010011",24338 => "11011101",24339 => "00011000",24340 => "00100011",24341 => "00100000",24342 => "10001110",24343 => "01110011",24344 => "11100101",24345 => "10111111",24346 => "11110001",24347 => "01010001",24348 => "01100110",24349 => "11110000",24350 => "10110110",24351 => "11010001",24352 => "11101010",24353 => "10110000",24354 => "01010010",24355 => "10000101",24356 => "00101001",24357 => "00000100",24358 => "11011110",24359 => "01011101",24360 => "01101010",24361 => "00100001",24362 => "01010010",24363 => "01000111",24364 => "10111111",24365 => "00000000",24366 => "10111011",24367 => "10011100",24368 => "11000110",24369 => "00111101",24370 => "01000100",24371 => "01000100",24372 => "00011011",24373 => "01001111",24374 => "01110101",24375 => "11100111",24376 => "10101010",24377 => "10111010",24378 => "00000101",24379 => "00011111",24380 => "10110101",24381 => "10101001",24382 => "00110000",24383 => "01001010",24384 => "11011101",24385 => "00011110",24386 => "01000011",24387 => "10110011",24388 => "00000010",24389 => "10110111",24390 => "10110001",24391 => "01001011",24392 => "11110000",24393 => "11001000",24394 => "01011111",24395 => "01110011",24396 => "10000000",24397 => "11100001",24398 => "00011101",24399 => "11111101",24400 => "11000000",24401 => "01101100",24402 => "11100101",24403 => "01101101",24404 => "00000110",24405 => "10110101",24406 => "00011011",24407 => "11011111",24408 => "01011010",24409 => "10001001",24410 => "11010101",24411 => "01001010",24412 => "01110100",24413 => "00011101",24414 => "11010000",24415 => "10110010",24416 => "00001011",24417 => "00001011",24418 => "10100100",24419 => "00110001",24420 => "11101011",24421 => "01001110",24422 => "11010101",24423 => "01000001",24424 => "11100111",24425 => "01011001",24426 => "10111101",24427 => "11011001",24428 => "10111110",24429 => "01000100",24430 => "11111101",24431 => "10010110",24432 => "11011001",24433 => "01010010",24434 => "11010000",24435 => "11110110",24436 => "01110000",24437 => "01101100",24438 => "00100101",24439 => "11010100",24440 => "11110001",24441 => "10100111",24442 => "11001101",24443 => "00101011",24444 => "01101110",24445 => "10001001",24446 => "00001101",24447 => "00011101",24448 => "11101101",24449 => "11101001",24450 => "00011000",24451 => "00101110",24452 => "10111111",24453 => "11010111",24454 => "11111011",24455 => "00001010",24456 => "10111001",24457 => "11011100",24458 => "01101100",24459 => "00101011",24460 => "00100001",24461 => "11110110",24462 => "10001010",24463 => "11110110",24464 => "01111101",24465 => "11011111",24466 => "00011000",24467 => "10111111",24468 => "10000010",24469 => "10001000",24470 => "10110110",24471 => "10101110",24472 => "10110101",24473 => "11011010",24474 => "00100110",24475 => "00111010",24476 => "10001100",24477 => "01101010",24478 => "10110011",24479 => "01111011",24480 => "01111111",24481 => "01110110",24482 => "01011010",24483 => "10001010",24484 => "10011110",24485 => "11100000",24486 => "00110111",24487 => "11011011",24488 => "11011010",24489 => "11010111",24490 => "01010010",24491 => "10010010",24492 => "11101110",24493 => "01010101",24494 => "00010101",24495 => "00011001",24496 => "00010101",24497 => "10110110",24498 => "01100110",24499 => "10110101",24500 => "00101111",24501 => "00001010",24502 => "11101000",24503 => "00001010",24504 => "10001100",24505 => "10100000",24506 => "00011001",24507 => "11101111",24508 => "10101101",24509 => "01111001",24510 => "10101001",24511 => "10101101",24512 => "01101110",24513 => "10011101",24514 => "11001111",24515 => "01100001",24516 => "11011110",24517 => "11111011",24518 => "10001111",24519 => "00110011",24520 => "00101010",24521 => "00110001",24522 => "10011110",24523 => "11001100",24524 => "00100110",24525 => "10100111",24526 => "01100110",24527 => "11100000",24528 => "00010110",24529 => "00001111",24530 => "00000001",24531 => "01010101",24532 => "10101100",24533 => "01110001",24534 => "00110111",24535 => "10110110",24536 => "10000100",24537 => "00100110",24538 => "10000011",24539 => "10001111",24540 => "00000100",24541 => "00001111",24542 => "00100010",24543 => "11010000",24544 => "11110001",24545 => "10010111",24546 => "10010101",24547 => "11110110",24548 => "01110000",24549 => "00111011",24550 => "11011100",24551 => "11100110",24552 => "01101111",24553 => "11011000",24554 => "00101100",24555 => "10101001",24556 => "01100001",24557 => "00011110",24558 => "01100010",24559 => "00000001",24560 => "11000000",24561 => "00010001",24562 => "11101000",24563 => "11001000",24564 => "00101001",24565 => "11000100",24566 => "11011101",24567 => "10001001",24568 => "11110011",24569 => "00101110",24570 => "01010111",24571 => "01000011",24572 => "10110011",24573 => "10100101",24574 => "01000101",24575 => "10101100",24576 => "01111000",24577 => "11011101",24578 => "11011101",24579 => "10100100",24580 => "01011001",24581 => "10001101",24582 => "00000001",24583 => "00000111",24584 => "01011111",24585 => "00001001",24586 => "01110101",24587 => "11110110",24588 => "00011010",24589 => "10001010",24590 => "11110011",24591 => "01000110",24592 => "11010100",24593 => "11000001",24594 => "10010100",24595 => "01011101",24596 => "10011111",24597 => "01101111",24598 => "01010011",24599 => "10011011",24600 => "00000001",24601 => "11101100",24602 => "00001111",24603 => "11110110",24604 => "00011001",24605 => "10101111",24606 => "10001000",24607 => "01100010",24608 => "01011110",24609 => "01001010",24610 => "11100011",24611 => "10100111",24612 => "01011100",24613 => "11000000",24614 => "00000101",24615 => "11000010",24616 => "01110001",24617 => "01010001",24618 => "01000100",24619 => "00100000",24620 => "01010101",24621 => "01000001",24622 => "11100001",24623 => "11100110",24624 => "00010100",24625 => "10011000",24626 => "11111110",24627 => "00000000",24628 => "11111100",24629 => "00100110",24630 => "00011100",24631 => "10101101",24632 => "01111100",24633 => "10100110",24634 => "10010100",24635 => "00001111",24636 => "10101011",24637 => "00001110",24638 => "10011001",24639 => "10110001",24640 => "00001101",24641 => "11101110",24642 => "01110000",24643 => "11110010",24644 => "11111100",24645 => "00101011",24646 => "00010101",24647 => "10111101",24648 => "10011011",24649 => "00101000",24650 => "10110101",24651 => "11001111",24652 => "01010000",24653 => "00100111",24654 => "00010000",24655 => "01001110",24656 => "11111011",24657 => "01011101",24658 => "00111101",24659 => "00110000",24660 => "00110011",24661 => "11100101",24662 => "00001001",24663 => "00110000",24664 => "01000111",24665 => "10101100",24666 => "10100110",24667 => "00101111",24668 => "01101011",24669 => "01101110",24670 => "00000101",24671 => "11001110",24672 => "00001000",24673 => "11011010",24674 => "00101000",24675 => "10000100",24676 => "11111010",24677 => "00111011",24678 => "00010011",24679 => "00111101",24680 => "00100001",24681 => "11001011",24682 => "11100001",24683 => "00000001",24684 => "00101111",24685 => "11100110",24686 => "11011011",24687 => "00000100",24688 => "11110111",24689 => "00111001",24690 => "11100100",24691 => "01001001",24692 => "00000010",24693 => "01001011",24694 => "00011000",24695 => "00011110",24696 => "00110101",24697 => "10110101",24698 => "01011011",24699 => "00011110",24700 => "11110111",24701 => "11111111",24702 => "00111000",24703 => "10011111",24704 => "00000000",24705 => "11100101",24706 => "01011101",24707 => "00100110",24708 => "11010101",24709 => "10001100",24710 => "01001001",24711 => "10110010",24712 => "11101001",24713 => "01111101",24714 => "11101110",24715 => "10101000",24716 => "01111000",24717 => "10010001",24718 => "01111011",24719 => "01110111",24720 => "01010001",24721 => "10001011",24722 => "10000100",24723 => "11010101",24724 => "10010110",24725 => "01000001",24726 => "10111111",24727 => "11101000",24728 => "01001111",24729 => "11100011",24730 => "10110111",24731 => "11110101",24732 => "00001101",24733 => "11001111",24734 => "11011100",24735 => "01110011",24736 => "10011010",24737 => "00000001",24738 => "01110001",24739 => "10111101",24740 => "01101110",24741 => "11111111",24742 => "01101110",24743 => "10001111",24744 => "01100001",24745 => "01110011",24746 => "01000011",24747 => "00000010",24748 => "11101001",24749 => "00111100",24750 => "11110011",24751 => "01010101",24752 => "01011010",24753 => "01000000",24754 => "10100010",24755 => "00001010",24756 => "10111010",24757 => "00100100",24758 => "01000011",24759 => "11111110",24760 => "01111101",24761 => "11100001",24762 => "01110000",24763 => "10001011",24764 => "11101100",24765 => "11111101",24766 => "11000010",24767 => "00011001",24768 => "01111001",24769 => "00001011",24770 => "10010110",24771 => "00010010",24772 => "00000001",24773 => "01110111",24774 => "01110000",24775 => "10101011",24776 => "10100111",24777 => "11001000",24778 => "00010100",24779 => "01010011",24780 => "11111101",24781 => "01111010",24782 => "01101010",24783 => "10111010",24784 => "01010111",24785 => "00100011",24786 => "10001100",24787 => "01110101",24788 => "10110110",24789 => "11001110",24790 => "00111110",24791 => "10011001",24792 => "10011101",24793 => "00110011",24794 => "10110001",24795 => "10111000",24796 => "10000011",24797 => "10101111",24798 => "11001111",24799 => "00100111",24800 => "10110100",24801 => "01100111",24802 => "11000101",24803 => "00101001",24804 => "01011100",24805 => "10010011",24806 => "00101001",24807 => "01000110",24808 => "00001001",24809 => "00110101",24810 => "00100110",24811 => "00100010",24812 => "01011001",24813 => "11110101",24814 => "00000010",24815 => "10110101",24816 => "10011110",24817 => "01111000",24818 => "01100100",24819 => "01100110",24820 => "01001000",24821 => "11011011",24822 => "11011011",24823 => "11100001",24824 => "01100000",24825 => "00101100",24826 => "10000111",24827 => "11010001",24828 => "11010110",24829 => "11001100",24830 => "01000111",24831 => "01100011",24832 => "01001110",24833 => "10100100",24834 => "00001010",24835 => "00011011",24836 => "10010010",24837 => "11101001",24838 => "11000110",24839 => "00100011",24840 => "11010101",24841 => "00101101",24842 => "00100101",24843 => "00001111",24844 => "10101111",24845 => "00001100",24846 => "00001000",24847 => "00110000",24848 => "01111111",24849 => "01010011",24850 => "11011100",24851 => "00010101",24852 => "11011010",24853 => "01011001",24854 => "01011011",24855 => "00110100",24856 => "01000010",24857 => "00011110",24858 => "00110100",24859 => "01100101",24860 => "11000000",24861 => "10000011",24862 => "10011011",24863 => "01101000",24864 => "10010001",24865 => "11011110",24866 => "00100001",24867 => "01110000",24868 => "00000000",24869 => "00000000",24870 => "01011101",24871 => "01101010",24872 => "01001100",24873 => "10011100",24874 => "01110011",24875 => "11001100",24876 => "01001010",24877 => "00010001",24878 => "11001010",24879 => "10111100",24880 => "01001000",24881 => "00001011",24882 => "10000011",24883 => "11000010",24884 => "01100011",24885 => "01111101",24886 => "10100000",24887 => "10110101",24888 => "00100010",24889 => "11001011",24890 => "10110100",24891 => "11111111",24892 => "00101101",24893 => "01011010",24894 => "00111111",24895 => "10000101",24896 => "10100100",24897 => "11111011",24898 => "00101001",24899 => "00111100",24900 => "01011101",24901 => "00011110",24902 => "01110010",24903 => "01101001",24904 => "11110011",24905 => "01011111",24906 => "11010100",24907 => "11111001",24908 => "01010101",24909 => "11011001",24910 => "01001000",24911 => "11011111",24912 => "01011111",24913 => "10000111",24914 => "11001011",24915 => "00011110",24916 => "10110000",24917 => "10110111",24918 => "00010101",24919 => "11111111",24920 => "10110011",24921 => "10001001",24922 => "11110001",24923 => "01110001",24924 => "11001110",24925 => "11111111",24926 => "11011100",24927 => "00010101",24928 => "00110111",24929 => "10001000",24930 => "10111101",24931 => "10100100",24932 => "10100111",24933 => "11010010",24934 => "10001101",24935 => "01110000",24936 => "10010101",24937 => "00101111",24938 => "00110010",24939 => "01110110",24940 => "01000100",24941 => "00111100",24942 => "00011001",24943 => "00101100",24944 => "00001010",24945 => "01111011",24946 => "11011100",24947 => "01100101",24948 => "11111010",24949 => "10000011",24950 => "01101011",24951 => "01110100",24952 => "00010100",24953 => "11101001",24954 => "00011001",24955 => "11000111",24956 => "10111000",24957 => "10001110",24958 => "11001010",24959 => "01100110",24960 => "00000010",24961 => "00101001",24962 => "11110111",24963 => "10011010",24964 => "01101101",24965 => "01110001",24966 => "11000011",24967 => "11100111",24968 => "11010010",24969 => "00110010",24970 => "01111011",24971 => "10010101",24972 => "10110010",24973 => "11100100",24974 => "10110111",24975 => "10100001",24976 => "01000000",24977 => "10101111",24978 => "01110001",24979 => "10011111",24980 => "01011011",24981 => "10001110",24982 => "01000011",24983 => "00101011",24984 => "00100001",24985 => "10111001",24986 => "10010010",24987 => "10001010",24988 => "10001110",24989 => "00100110",24990 => "11001001",24991 => "00110001",24992 => "01111000",24993 => "10100001",24994 => "00001111",24995 => "00101001",24996 => "10101001",24997 => "01100111",24998 => "11010010",24999 => "10111010",25000 => "00100000",25001 => "10100110",25002 => "00011001",25003 => "01000011",25004 => "00000011",25005 => "00000000",25006 => "11001000",25007 => "00101001",25008 => "11110110",25009 => "00110111",25010 => "10101100",25011 => "01100100",25012 => "11101110",25013 => "01110001",25014 => "01001000",25015 => "01101010",25016 => "01011010",25017 => "00111000",25018 => "11001001",25019 => "01011011",25020 => "01101101",25021 => "10101100",25022 => "01011100",25023 => "10101010",25024 => "00110100",25025 => "11111100",25026 => "10100111",25027 => "11000111",25028 => "00010101",25029 => "10011111",25030 => "11110010",25031 => "00101001",25032 => "11110001",25033 => "11111100",25034 => "00111101",25035 => "11101001",25036 => "01100111",25037 => "11111110",25038 => "01101001",25039 => "11111111",25040 => "11100101",25041 => "01010100",25042 => "11010011",25043 => "11010100",25044 => "10000011",25045 => "00010111",25046 => "10011110",25047 => "01011111",25048 => "11100100",25049 => "11110001",25050 => "00010010",25051 => "00010111",25052 => "11010100",25053 => "01101101",25054 => "11011110",25055 => "11000110",25056 => "10010111",25057 => "00110101",25058 => "10000011",25059 => "00000001",25060 => "01110010",25061 => "00111110",25062 => "01001000",25063 => "11010110",25064 => "11010100",25065 => "01001010",25066 => "01101101",25067 => "10110100",25068 => "11110011",25069 => "11011111",25070 => "10110001",25071 => "01000010",25072 => "10001011",25073 => "01111100",25074 => "00110111",25075 => "10111000",25076 => "01101100",25077 => "11111011",25078 => "10110010",25079 => "11000110",25080 => "10110011",25081 => "10101001",25082 => "10000001",25083 => "01101011",25084 => "11101000",25085 => "00001000",25086 => "01101100",25087 => "11110110",25088 => "11100100",25089 => "10100000",25090 => "10111111",25091 => "01100101",25092 => "00111001",25093 => "00101010",25094 => "10001010",25095 => "11011010",25096 => "00001100",25097 => "11100110",25098 => "11011111",25099 => "11100010",25100 => "01001011",25101 => "11100000",25102 => "11010000",25103 => "11001011",25104 => "11010100",25105 => "10110011",25106 => "10111011",25107 => "10111011",25108 => "00110011",25109 => "00000100",25110 => "00110011",25111 => "10011111",25112 => "00110010",25113 => "00000010",25114 => "01010000",25115 => "01001011",25116 => "11110111",25117 => "10111010",25118 => "01100000",25119 => "00101001",25120 => "10010001",25121 => "11101110",25122 => "11110001",25123 => "10011010",25124 => "00110000",25125 => "11010011",25126 => "01100010",25127 => "10011011",25128 => "01111000",25129 => "10011010",25130 => "11011111",25131 => "00101100",25132 => "01111000",25133 => "11001011",25134 => "01001101",25135 => "11010010",25136 => "11010001",25137 => "10000111",25138 => "11011100",25139 => "11010001",25140 => "01111010",25141 => "01000010",25142 => "00110000",25143 => "10101111",25144 => "11010100",25145 => "00001110",25146 => "10100110",25147 => "00010001",25148 => "10110010",25149 => "11101000",25150 => "01000110",25151 => "01010010",25152 => "11100000",25153 => "00011110",25154 => "01110011",25155 => "01011111",25156 => "11101110",25157 => "10011100",25158 => "11000010",25159 => "00110011",25160 => "01011000",25161 => "01111110",25162 => "00110010",25163 => "00011101",25164 => "11111110",25165 => "00010001",25166 => "11100110",25167 => "11010111",25168 => "11010000",25169 => "10010100",25170 => "11000011",25171 => "11111111",25172 => "11000101",25173 => "00100101",25174 => "01110010",25175 => "11101001",25176 => "01011111",25177 => "00001101",25178 => "10011001",25179 => "10110001",25180 => "10111111",25181 => "00010010",25182 => "11010100",25183 => "10011110",25184 => "11100001",25185 => "01001000",25186 => "00001110",25187 => "01100101",25188 => "01110000",25189 => "10110111",25190 => "10101000",25191 => "10100110",25192 => "10000011",25193 => "10101111",25194 => "10111001",25195 => "10010001",25196 => "11001011",25197 => "01111010",25198 => "11111010",25199 => "00011101",25200 => "10111100",25201 => "10110000",25202 => "01011000",25203 => "10000001",25204 => "10110011",25205 => "01010010",25206 => "00010011",25207 => "10010111",25208 => "01100011",25209 => "11101111",25210 => "01010011",25211 => "10111110",25212 => "00110101",25213 => "11101101",25214 => "10111100",25215 => "01100110",25216 => "10111010",25217 => "01101010",25218 => "01000101",25219 => "00010101",25220 => "00000001",25221 => "00100000",25222 => "10110111",25223 => "01011010",25224 => "10001000",25225 => "00011111",25226 => "10010110",25227 => "01100001",25228 => "11010110",25229 => "11001010",25230 => "00101001",25231 => "11010001",25232 => "11011000",25233 => "00011011",25234 => "10111000",25235 => "11011000",25236 => "01101101",25237 => "10100110",25238 => "01000010",25239 => "01011011",25240 => "01000100",25241 => "00100011",25242 => "10001001",25243 => "01101101",25244 => "10010000",25245 => "11000101",25246 => "01110001",25247 => "11111010",25248 => "10101100",25249 => "10001111",25250 => "10001010",25251 => "00010110",25252 => "10001001",25253 => "11110011",25254 => "01101001",25255 => "10001000",25256 => "11001100",25257 => "11011101",25258 => "10101110",25259 => "10000100",25260 => "01101100",25261 => "01111011",25262 => "10111101",25263 => "01101100",25264 => "10110011",25265 => "11011011",25266 => "11100001",25267 => "00100101",25268 => "11001000",25269 => "10010000",25270 => "11000010",25271 => "10111110",25272 => "10000101",25273 => "01100110",25274 => "01100110",25275 => "10010101",25276 => "11010111",25277 => "01001010",25278 => "01101001",25279 => "01100100",25280 => "10100100",25281 => "01100010",25282 => "11110011",25283 => "11001010",25284 => "01000011",25285 => "11000000",25286 => "10110111",25287 => "11011100",25288 => "00100011",25289 => "00110000",25290 => "01100001",25291 => "10111011",25292 => "01101101",25293 => "10010100",25294 => "01010100",25295 => "00010100",25296 => "00100100",25297 => "11101110",25298 => "10000100",25299 => "00100101",25300 => "01111001",25301 => "00000100",25302 => "01111110",25303 => "01110111",25304 => "00001100",25305 => "01100101",25306 => "00010101",25307 => "01100001",25308 => "01110010",25309 => "01110001",25310 => "11100111",25311 => "01010000",25312 => "10101001",25313 => "00000100",25314 => "01000000",25315 => "00100001",25316 => "10101010",25317 => "01111101",25318 => "10111001",25319 => "10001111",25320 => "10001000",25321 => "11000111",25322 => "11111011",25323 => "11110010",25324 => "01001011",25325 => "10100011",25326 => "00010110",25327 => "11001111",25328 => "01110010",25329 => "10001110",25330 => "00010100",25331 => "11100110",25332 => "10010101",25333 => "11111000",25334 => "00110011",25335 => "10110100",25336 => "00010010",25337 => "11111111",25338 => "00111010",25339 => "10001111",25340 => "01001010",25341 => "10000111",25342 => "00001001",25343 => "00000100",25344 => "10000011",25345 => "01110000",25346 => "00000011",25347 => "10111110",25348 => "11110110",25349 => "01001111",25350 => "01111010",25351 => "11100101",25352 => "01100101",25353 => "01011111",25354 => "00100000",25355 => "00111000",25356 => "01111110",25357 => "10101101",25358 => "00010110",25359 => "11110100",25360 => "00010001",25361 => "11111010",25362 => "00001101",25363 => "01010111",25364 => "01110011",25365 => "01110011",25366 => "00110011",25367 => "00110110",25368 => "10000100",25369 => "10110111",25370 => "11111101",25371 => "11101011",25372 => "00000101",25373 => "10010010",25374 => "01111010",25375 => "01011111",25376 => "11110000",25377 => "01010001",25378 => "00110110",25379 => "00001011",25380 => "01111000",25381 => "01110001",25382 => "01001010",25383 => "00100011",25384 => "10110011",25385 => "01101001",25386 => "01001000",25387 => "11010101",25388 => "01101101",25389 => "10111110",25390 => "00010111",25391 => "10101100",25392 => "01010001",25393 => "01110100",25394 => "10000010",25395 => "11001001",25396 => "01001101",25397 => "11000000",25398 => "11100110",25399 => "11100000",25400 => "01101100",25401 => "01000111",25402 => "10111000",25403 => "11100010",25404 => "01111100",25405 => "01000011",25406 => "01001011",25407 => "10011100",25408 => "00000101",25409 => "01101011",25410 => "00111100",25411 => "01011110",25412 => "10111100",25413 => "11101100",25414 => "10100111",25415 => "10111011",25416 => "10001100",25417 => "10001010",25418 => "11101101",25419 => "00111110",25420 => "11100010",25421 => "00011110",25422 => "00001000",25423 => "10001010",25424 => "11001111",25425 => "10011000",25426 => "00000101",25427 => "01011100",25428 => "00000110",25429 => "01100001",25430 => "00011101",25431 => "11001101",25432 => "11000010",25433 => "11010100",25434 => "00011001",25435 => "01000011",25436 => "01000101",25437 => "10011110",25438 => "11011001",25439 => "01101101",25440 => "10100011",25441 => "11100100",25442 => "00011111",25443 => "00111000",25444 => "01111110",25445 => "01010110",25446 => "11011101",25447 => "11000001",25448 => "01111011",25449 => "11110011",25450 => "00100011",25451 => "11100001",25452 => "11001110",25453 => "00011100",25454 => "01100010",25455 => "01000110",25456 => "01000001",25457 => "11101101",25458 => "00011011",25459 => "01000101",25460 => "01101111",25461 => "11111101",25462 => "01010111",25463 => "10110110",25464 => "10001010",25465 => "01010001",25466 => "01011010",25467 => "00101000",25468 => "00111011",25469 => "11001010",25470 => "00111110",25471 => "01010111",25472 => "10111100",25473 => "11010010",25474 => "10100111",25475 => "00011111",25476 => "00100101",25477 => "01101010",25478 => "01110001",25479 => "01101111",25480 => "00000110",25481 => "10011101",25482 => "10100111",25483 => "00011010",25484 => "10000010",25485 => "11010101",25486 => "00011011",25487 => "10011110",25488 => "01000100",25489 => "10100110",25490 => "10111111",25491 => "11000110",25492 => "01101011",25493 => "00000000",25494 => "00101100",25495 => "10000000",25496 => "00111110",25497 => "01001101",25498 => "10110000",25499 => "11111000",25500 => "00101101",25501 => "10111000",25502 => "10100010",25503 => "11010101",25504 => "11000110",25505 => "11100000",25506 => "01011001",25507 => "10001100",25508 => "10010111",25509 => "00010101",25510 => "00111100",25511 => "01011110",25512 => "11011101",25513 => "00001010",25514 => "10010100",25515 => "00100001",25516 => "11001100",25517 => "10100111",25518 => "00011001",25519 => "11101001",25520 => "00011100",25521 => "01111010",25522 => "10011111",25523 => "01000111",25524 => "11001010",25525 => "01101110",25526 => "10000111",25527 => "11111100",25528 => "01001100",25529 => "11001101",25530 => "11100001",25531 => "00110010",25532 => "10101010",25533 => "00110111",25534 => "00010101",25535 => "11100111",25536 => "00100001",25537 => "11101101",25538 => "11001101",25539 => "00110101",25540 => "10101100",25541 => "00100110",25542 => "11001000",25543 => "00100011",25544 => "10001001",25545 => "00000110",25546 => "00000011",25547 => "11011110",25548 => "10010100",25549 => "00001110",25550 => "00111110",25551 => "10011111",25552 => "01001110",25553 => "00001011",25554 => "11110010",25555 => "10001110",25556 => "01000101",25557 => "00110011",25558 => "01000001",25559 => "10111110",25560 => "00001100",25561 => "01000001",25562 => "00100101",25563 => "11011011",25564 => "00111011",25565 => "11011111",25566 => "01100000",25567 => "10100000",25568 => "00101101",25569 => "01101101",25570 => "01001101",25571 => "01100000",25572 => "00000100",25573 => "10110010",25574 => "00100001",25575 => "11010110",25576 => "10101101",25577 => "00101010",25578 => "00011100",25579 => "10111000",25580 => "01101010",25581 => "01101111",25582 => "01101100",25583 => "10001000",25584 => "10001110",25585 => "10011001",25586 => "10100011",25587 => "11110001",25588 => "10111100",25589 => "00000110",25590 => "01110000",25591 => "01011101",25592 => "10100010",25593 => "10010001",25594 => "00010101",25595 => "00101000",25596 => "11011000",25597 => "00011111",25598 => "10100000",25599 => "00100011",25600 => "11101001",25601 => "11100000",25602 => "00111000",25603 => "11010001",25604 => "10001001",25605 => "01011111",25606 => "11010100",25607 => "11011111",25608 => "01111001",25609 => "01010010",25610 => "01110111",25611 => "11001111",25612 => "00010101",25613 => "10111110",25614 => "10101110",25615 => "00100001",25616 => "00011110",25617 => "00111101",25618 => "00110100",25619 => "10010001",25620 => "01000100",25621 => "00100111",25622 => "10001001",25623 => "01011011",25624 => "10011101",25625 => "00011001",25626 => "01011010",25627 => "00001010",25628 => "11101110",25629 => "01001101",25630 => "01111101",25631 => "10111011",25632 => "01001101",25633 => "01101001",25634 => "01001101",25635 => "00000100",25636 => "00001001",25637 => "00101001",25638 => "10011010",25639 => "01111001",25640 => "01101100",25641 => "01111100",25642 => "00000011",25643 => "11010100",25644 => "10100000",25645 => "00101001",25646 => "11010111",25647 => "01111001",25648 => "00000011",25649 => "11000011",25650 => "11010100",25651 => "10111100",25652 => "11010001",25653 => "10100001",25654 => "11011100",25655 => "00110101",25656 => "11000111",25657 => "00001101",25658 => "01011000",25659 => "10100100",25660 => "11010000",25661 => "01001110",25662 => "11110100",25663 => "01101111",25664 => "10100110",25665 => "11000010",25666 => "11110000",25667 => "10101101",25668 => "11011110",25669 => "00110010",25670 => "01001101",25671 => "00001110",25672 => "00110100",25673 => "01111010",25674 => "00000000",25675 => "10010001",25676 => "10110000",25677 => "11000110",25678 => "10000110",25679 => "01100011",25680 => "01001101",25681 => "00001110",25682 => "01100001",25683 => "00011001",25684 => "00010011",25685 => "00001110",25686 => "00000001",25687 => "01100100",25688 => "11111110",25689 => "11000111",25690 => "11110001",25691 => "10001110",25692 => "10001000",25693 => "00110100",25694 => "11011101",25695 => "11110010",25696 => "01001100",25697 => "11101001",25698 => "11001011",25699 => "11010011",25700 => "11010001",25701 => "11010100",25702 => "11110011",25703 => "00001000",25704 => "11011110",25705 => "10001111",25706 => "00110011",25707 => "01101010",25708 => "00110010",25709 => "00011010",25710 => "11011110",25711 => "11010011",25712 => "11111100",25713 => "01110101",25714 => "01100111",25715 => "00111100",25716 => "11110110",25717 => "01000001",25718 => "10000111",25719 => "00011011",25720 => "01100010",25721 => "10001010",25722 => "01101100",25723 => "01011000",25724 => "01110111",25725 => "11110001",25726 => "00001100",25727 => "00101101",25728 => "00010111",25729 => "10001011",25730 => "11100101",25731 => "01111001",25732 => "10111101",25733 => "00110110",25734 => "01100010",25735 => "00001101",25736 => "00100110",25737 => "00101101",25738 => "00001110",25739 => "11010100",25740 => "11101010",25741 => "11101010",25742 => "01100111",25743 => "10011100",25744 => "01100011",25745 => "00111110",25746 => "11101011",25747 => "11000010",25748 => "01010000",25749 => "11000101",25750 => "00000100",25751 => "10101101",25752 => "00000100",25753 => "00000011",25754 => "00000110",25755 => "11010011",25756 => "01000110",25757 => "10011000",25758 => "10001011",25759 => "01110011",25760 => "11010101",25761 => "01110000",25762 => "00100100",25763 => "01100010",25764 => "10101010",25765 => "01001101",25766 => "00100101",25767 => "01010000",25768 => "00011101",25769 => "00100111",25770 => "11101101",25771 => "11110010",25772 => "11111001",25773 => "11101000",25774 => "00010000",25775 => "00100000",25776 => "00001011",25777 => "00001000",25778 => "01111101",25779 => "10111101",25780 => "01010101",25781 => "10001100",25782 => "01010001",25783 => "01010000",25784 => "10100101",25785 => "11010100",25786 => "10011100",25787 => "01111101",25788 => "01011101",25789 => "00101100",25790 => "10001110",25791 => "01011110",25792 => "10100001",25793 => "11110110",25794 => "00100001",25795 => "00101010",25796 => "00101011",25797 => "00001001",25798 => "11001101",25799 => "11010110",25800 => "01101111",25801 => "10000011",25802 => "10110111",25803 => "00011100",25804 => "10100000",25805 => "01100001",25806 => "00110000",25807 => "11101010",25808 => "00001010",25809 => "00100000",25810 => "10110111",25811 => "01100110",25812 => "10000010",25813 => "01100000",25814 => "01110011",25815 => "10001101",25816 => "00101101",25817 => "00000111",25818 => "10111111",25819 => "01101011",25820 => "01111110",25821 => "10011000",25822 => "01010101",25823 => "10101000",25824 => "01010010",25825 => "01001111",25826 => "11010000",25827 => "10101110",25828 => "10000111",25829 => "11001001",25830 => "11001100",25831 => "00101100",25832 => "10100101",25833 => "10000111",25834 => "10011010",25835 => "00111100",25836 => "10101011",25837 => "11111101",25838 => "00111111",25839 => "10110100",25840 => "11101101",25841 => "10010011",25842 => "11111101",25843 => "00010011",25844 => "01111011",25845 => "01111001",25846 => "00110011",25847 => "11001110",25848 => "11100111",25849 => "10000111",25850 => "11100101",25851 => "01001001",25852 => "01011111",25853 => "11101000",25854 => "00111011",25855 => "01111110",25856 => "10011000",25857 => "00001010",25858 => "11100111",25859 => "01011100",25860 => "01001011",25861 => "00101011",25862 => "00011010",25863 => "00010101",25864 => "01001010",25865 => "10110010",25866 => "11001011",25867 => "11111010",25868 => "00010001",25869 => "00101001",25870 => "01010101",25871 => "01000100",25872 => "01100110",25873 => "01000011",25874 => "10110110",25875 => "01111111",25876 => "11001110",25877 => "01111101",25878 => "01011011",25879 => "00011100",25880 => "11001100",25881 => "01010010",25882 => "11110111",25883 => "00110001",25884 => "10110000",25885 => "11100011",25886 => "10000000",25887 => "00011001",25888 => "01001000",25889 => "10001010",25890 => "00100110",25891 => "10111110",25892 => "00111001",25893 => "01101000",25894 => "11001110",25895 => "00011110",25896 => "11101011",25897 => "00001011",25898 => "00101010",25899 => "00100011",25900 => "00100000",25901 => "10000011",25902 => "00010100",25903 => "10101001",25904 => "10010101",25905 => "01011110",25906 => "10101100",25907 => "10001111",25908 => "11100100",25909 => "10100000",25910 => "10011010",25911 => "00110011",25912 => "01111100",25913 => "11011000",25914 => "10010001",25915 => "01001011",25916 => "01100100",25917 => "00100110",25918 => "00011101",25919 => "10100111",25920 => "11100000",25921 => "01001000",25922 => "01010000",25923 => "00011100",25924 => "01011100",25925 => "00101101",25926 => "00010100",25927 => "11111111",25928 => "01100010",25929 => "11110010",25930 => "11011111",25931 => "00000101",25932 => "11100001",25933 => "00111110",25934 => "00100011",25935 => "00010100",25936 => "01010100",25937 => "11000111",25938 => "11011010",25939 => "00101000",25940 => "10010111",25941 => "01011001",25942 => "10000001",25943 => "00101110",25944 => "00111001",25945 => "01101111",25946 => "10110101",25947 => "10011110",25948 => "11110010",25949 => "01100110",25950 => "11101010",25951 => "11110111",25952 => "10000111",25953 => "01000001",25954 => "10100010",25955 => "00000111",25956 => "10100111",25957 => "01010000",25958 => "11110101",25959 => "01011000",25960 => "10100001",25961 => "11101110",25962 => "01101001",25963 => "01101010",25964 => "00110101",25965 => "11011011",25966 => "00100010",25967 => "00111011",25968 => "00001010",25969 => "00110001",25970 => "11001101",25971 => "00001111",25972 => "00100101",25973 => "11011100",25974 => "10100000",25975 => "01010101",25976 => "01110000",25977 => "11010101",25978 => "00110001",25979 => "11111010",25980 => "01001000",25981 => "11010000",25982 => "10100000",25983 => "01000100",25984 => "01101010",25985 => "01010000",25986 => "00010110",25987 => "10011000",25988 => "11111010",25989 => "11010111",25990 => "10100111",25991 => "00111100",25992 => "11000111",25993 => "10111111",25994 => "11010101",25995 => "10100011",25996 => "01001100",25997 => "01010100",25998 => "10100111",25999 => "10110101",26000 => "11110101",26001 => "10010011",26002 => "11111011",26003 => "00011111",26004 => "11001001",26005 => "10100100",26006 => "00101100",26007 => "11111010",26008 => "00101100",26009 => "01100011",26010 => "10000001",26011 => "00110100",26012 => "10010010",26013 => "10010001",26014 => "11101001",26015 => "01000101",26016 => "01001000",26017 => "00011000",26018 => "11110011",26019 => "01001100",26020 => "11011010",26021 => "11001100",26022 => "11001010",26023 => "10101110",26024 => "00011000",26025 => "10000110",26026 => "11111000",26027 => "10010111",26028 => "11000111",26029 => "00100010",26030 => "11000010",26031 => "10000010",26032 => "11110010",26033 => "11001010",26034 => "10000011",26035 => "11001110",26036 => "00110110",26037 => "00101111",26038 => "00000010",26039 => "01100111",26040 => "11011110",26041 => "00101001",26042 => "10011001",26043 => "10101101",26044 => "01010010",26045 => "01110010",26046 => "00001001",26047 => "00100011",26048 => "10110110",26049 => "00000010",26050 => "11100011",26051 => "11001011",26052 => "01110101",26053 => "01010000",26054 => "01011010",26055 => "10011011",26056 => "00100111",26057 => "11001100",26058 => "10100101",26059 => "00110100",26060 => "01100001",26061 => "10100011",26062 => "10011011",26063 => "01101111",26064 => "10111101",26065 => "11101000",26066 => "11110111",26067 => "10001000",26068 => "11001011",26069 => "00001001",26070 => "00011010",26071 => "11101110",26072 => "00001100",26073 => "01101001",26074 => "00010001",26075 => "11000011",26076 => "00001111",26077 => "00000100",26078 => "01010100",26079 => "00011110",26080 => "11110100",26081 => "00010001",26082 => "11111111",26083 => "00010111",26084 => "11111000",26085 => "11010001",26086 => "00001001",26087 => "11100001",26088 => "00111101",26089 => "10011001",26090 => "11111110",26091 => "01100011",26092 => "11110001",26093 => "10111101",26094 => "10011111",26095 => "10110010",26096 => "10101010",26097 => "00010011",26098 => "11110000",26099 => "00101000",26100 => "11011000",26101 => "10001110",26102 => "10010001",26103 => "00111001",26104 => "11000101",26105 => "01000010",26106 => "11000011",26107 => "11000101",26108 => "11111010",26109 => "10011011",26110 => "01111100",26111 => "00101001",26112 => "10011011",26113 => "11101101",26114 => "01000001",26115 => "10001001",26116 => "00001001",26117 => "01100111",26118 => "00110101",26119 => "00101101",26120 => "11011111",26121 => "10101111",26122 => "00100001",26123 => "11101010",26124 => "10110010",26125 => "10010011",26126 => "10101111",26127 => "01001111",26128 => "00110110",26129 => "10010100",26130 => "00001001",26131 => "11110101",26132 => "10100111",26133 => "11001000",26134 => "01110100",26135 => "11011111",26136 => "11001110",26137 => "01110011",26138 => "10111010",26139 => "11001011",26140 => "11000000",26141 => "00110101",26142 => "11011100",26143 => "10110111",26144 => "11111001",26145 => "01010100",26146 => "00110100",26147 => "10000010",26148 => "00110110",26149 => "10010101",26150 => "10100001",26151 => "00111000",26152 => "01110110",26153 => "01110011",26154 => "00110110",26155 => "10000001",26156 => "10101100",26157 => "00001110",26158 => "01111110",26159 => "10100101",26160 => "10111100",26161 => "01000001",26162 => "01100110",26163 => "10101110",26164 => "01010000",26165 => "01000011",26166 => "10101010",26167 => "00010110",26168 => "01101011",26169 => "10101101",26170 => "01100101",26171 => "00001110",26172 => "01010101",26173 => "01010101",26174 => "11001010",26175 => "11100110",26176 => "11101010",26177 => "10100110",26178 => "01101100",26179 => "11111101",26180 => "11110001",26181 => "00100001",26182 => "10011111",26183 => "11011101",26184 => "11001110",26185 => "10110001",26186 => "11011010",26187 => "01001101",26188 => "01001111",26189 => "11010100",26190 => "01000010",26191 => "10111010",26192 => "00100010",26193 => "00000111",26194 => "00001100",26195 => "10111111",26196 => "10010100",26197 => "01010000",26198 => "00110101",26199 => "11110111",26200 => "11010110",26201 => "11111101",26202 => "01101011",26203 => "00011000",26204 => "10110101",26205 => "10110111",26206 => "10001111",26207 => "01100010",26208 => "01011101",26209 => "10110111",26210 => "01001100",26211 => "00011010",26212 => "10011001",26213 => "00011000",26214 => "10001110",26215 => "00001101",26216 => "00000000",26217 => "11100011",26218 => "00011001",26219 => "10000100",26220 => "11111011",26221 => "00001110",26222 => "11011100",26223 => "10011001",26224 => "11101100",26225 => "00001100",26226 => "10110011",26227 => "01111110",26228 => "00111110",26229 => "00001000",26230 => "01000100",26231 => "11111100",26232 => "01001110",26233 => "01011010",26234 => "10010011",26235 => "01101100",26236 => "11001000",26237 => "11110101",26238 => "00000001",26239 => "11100000",26240 => "10000010",26241 => "00101010",26242 => "10111000",26243 => "01111011",26244 => "00000111",26245 => "01100111",26246 => "01110100",26247 => "10010000",26248 => "11100001",26249 => "01111111",26250 => "10001011",26251 => "00111001",26252 => "11111011",26253 => "01101110",26254 => "10011101",26255 => "00101111",26256 => "01001011",26257 => "01011101",26258 => "00001110",26259 => "11001101",26260 => "11001111",26261 => "10011101",26262 => "10000011",26263 => "00101000",26264 => "10010100",26265 => "10011010",26266 => "11010010",26267 => "01011000",26268 => "10000100",26269 => "10000110",26270 => "11001101",26271 => "10011000",26272 => "00100000",26273 => "11100001",26274 => "10111100",26275 => "11101101",26276 => "10100100",26277 => "01011001",26278 => "00000011",26279 => "00100001",26280 => "10110100",26281 => "00101111",26282 => "11111111",26283 => "01111000",26284 => "11000001",26285 => "11111000",26286 => "10110001",26287 => "10110101",26288 => "10011010",26289 => "00100001",26290 => "00111111",26291 => "10010100",26292 => "00011110",26293 => "11101111",26294 => "01010110",26295 => "11010000",26296 => "01100000",26297 => "01101101",26298 => "01111100",26299 => "10101001",26300 => "11000010",26301 => "01101111",26302 => "00101110",26303 => "01000011",26304 => "11000000",26305 => "11100111",26306 => "10101001",26307 => "10100011",26308 => "11101000",26309 => "10010100",26310 => "10001010",26311 => "01101111",26312 => "11001111",26313 => "11010010",26314 => "01010010",26315 => "00000111",26316 => "00100001",26317 => "11011010",26318 => "00111001",26319 => "00001000",26320 => "01001101",26321 => "10010111",26322 => "01100110",26323 => "11010100",26324 => "10011100",26325 => "10000101",26326 => "00000101",26327 => "00001001",26328 => "11111001",26329 => "01011100",26330 => "10101101",26331 => "11111111",26332 => "11111111",26333 => "00110001",26334 => "00100000",26335 => "01111100",26336 => "01111000",26337 => "10101111",26338 => "00111001",26339 => "00000110",26340 => "11100001",26341 => "01011011",26342 => "11111100",26343 => "01010010",26344 => "11110100",26345 => "00110100",26346 => "10110011",26347 => "00100111",26348 => "00111111",26349 => "01100011",26350 => "10111001",26351 => "01011101",26352 => "01111100",26353 => "01100100",26354 => "01100001",26355 => "10001010",26356 => "00111001",26357 => "00000001",26358 => "00100101",26359 => "11000100",26360 => "11111100",26361 => "11010110",26362 => "10110010",26363 => "00000100",26364 => "00110101",26365 => "10101000",26366 => "00111100",26367 => "11001010",26368 => "00100110",26369 => "10110011",26370 => "00011101",26371 => "10001101",26372 => "11001011",26373 => "00011001",26374 => "00011101",26375 => "00000001",26376 => "10001011",26377 => "11110111",26378 => "01110111",26379 => "01010010",26380 => "10111001",26381 => "00101010",26382 => "00101111",26383 => "10001001",26384 => "11111100",26385 => "11111011",26386 => "00001100",26387 => "10111111",26388 => "00111100",26389 => "01111100",26390 => "00010100",26391 => "00000010",26392 => "11010000",26393 => "11111100",26394 => "01000011",26395 => "00011001",26396 => "01100001",26397 => "01011110",26398 => "01110011",26399 => "01101111",26400 => "11100101",26401 => "00000001",26402 => "01101011",26403 => "01101110",26404 => "11101100",26405 => "11010011",26406 => "10111110",26407 => "00101010",26408 => "01101000",26409 => "00110111",26410 => "11010100",26411 => "11000000",26412 => "00100001",26413 => "01111110",26414 => "00101100",26415 => "10010001",26416 => "11011011",26417 => "10110111",26418 => "01100101",26419 => "00110101",26420 => "10000100",26421 => "01001010",26422 => "11001100",26423 => "10011010",26424 => "01101000",26425 => "00010110",26426 => "10001110",26427 => "01001110",26428 => "11010100",26429 => "11100111",26430 => "01001001",26431 => "00010001",26432 => "11110010",26433 => "11100001",26434 => "10111010",26435 => "11010111",26436 => "00100001",26437 => "01010111",26438 => "10011010",26439 => "01111100",26440 => "11111100",26441 => "01011110",26442 => "00011011",26443 => "01010001",26444 => "01111011",26445 => "11010011",26446 => "11110111",26447 => "11101001",26448 => "00100000",26449 => "00001100",26450 => "11011101",26451 => "01111011",26452 => "00110010",26453 => "01000000",26454 => "00110011",26455 => "00101101",26456 => "11110010",26457 => "01011101",26458 => "01000011",26459 => "00011111",26460 => "10001010",26461 => "11011100",26462 => "11000000",26463 => "11100010",26464 => "10111011",26465 => "00011000",26466 => "10101101",26467 => "00011111",26468 => "11111001",26469 => "10000110",26470 => "00000001",26471 => "01111010",26472 => "10110001",26473 => "01001000",26474 => "00000110",26475 => "01111011",26476 => "11100111",26477 => "11000001",26478 => "11111110",26479 => "00111111",26480 => "01000110",26481 => "10100110",26482 => "11101101",26483 => "00011100",26484 => "11111111",26485 => "11000101",26486 => "11010010",26487 => "00001110",26488 => "00000110",26489 => "00100001",26490 => "01001001",26491 => "10000011",26492 => "01101001",26493 => "11001000",26494 => "01000010",26495 => "00101000",26496 => "10010101",26497 => "01100011",26498 => "10000101",26499 => "10101001",26500 => "00011001",26501 => "11111011",26502 => "00000010",26503 => "11011111",26504 => "01000010",26505 => "10110011",26506 => "11011100",26507 => "11010100",26508 => "01110001",26509 => "11010010",26510 => "10110100",26511 => "10101100",26512 => "11111001",26513 => "00001110",26514 => "10000000",26515 => "11000000",26516 => "11110000",26517 => "11110100",26518 => "00011001",26519 => "11010000",26520 => "11110000",26521 => "11101111",26522 => "00000111",26523 => "00000100",26524 => "01110000",26525 => "01110101",26526 => "00010010",26527 => "11011010",26528 => "00111111",26529 => "10110100",26530 => "11001101",26531 => "11111110",26532 => "00101001",26533 => "00001100",26534 => "00010111",26535 => "11111000",26536 => "00100010",26537 => "10010010",26538 => "11001010",26539 => "10011110",26540 => "11010010",26541 => "01110110",26542 => "00100111",26543 => "10101001",26544 => "11100000",26545 => "01000110",26546 => "00100010",26547 => "00100101",26548 => "10000110",26549 => "00011101",26550 => "00111101",26551 => "01100010",26552 => "01111000",26553 => "00011110",26554 => "00110101",26555 => "00010100",26556 => "00111001",26557 => "00010111",26558 => "00101101",26559 => "11010010",26560 => "10111000",26561 => "00010010",26562 => "11111000",26563 => "11001101",26564 => "11110111",26565 => "10110101",26566 => "00001110",26567 => "10100011",26568 => "00111000",26569 => "11100100",26570 => "00011110",26571 => "11110100",26572 => "00111011",26573 => "00000000",26574 => "10010110",26575 => "00001011",26576 => "10111111",26577 => "10001110",26578 => "01100110",26579 => "11000001",26580 => "01111011",26581 => "01100110",26582 => "00011110",26583 => "00001010",26584 => "00010010",26585 => "00011011",26586 => "01001001",26587 => "11010001",26588 => "10010011",26589 => "11000001",26590 => "01011110",26591 => "11001110",26592 => "11111010",26593 => "10011101",26594 => "00110001",26595 => "01001001",26596 => "11000010",26597 => "11101100",26598 => "10110111",26599 => "01011000",26600 => "01111001",26601 => "11011010",26602 => "10100101",26603 => "01101111",26604 => "11000110",26605 => "10100011",26606 => "10000011",26607 => "11111100",26608 => "11110011",26609 => "11011110",26610 => "10001011",26611 => "00001011",26612 => "11100100",26613 => "01101000",26614 => "11111110",26615 => "01001110",26616 => "01000000",26617 => "01111110",26618 => "11000000",26619 => "11101011",26620 => "10110111",26621 => "11011101",26622 => "11111110",26623 => "01000111",26624 => "01001101",26625 => "00010000",26626 => "00110100",26627 => "01011111",26628 => "10100011",26629 => "01000100",26630 => "10111010",26631 => "01010111",26632 => "11100100",26633 => "01111001",26634 => "00001011",26635 => "11100000",26636 => "11011110",26637 => "11111110",26638 => "11101101",26639 => "11011100",26640 => "00111100",26641 => "00011011",26642 => "01111101",26643 => "01000011",26644 => "00101010",26645 => "01101111",26646 => "10011010",26647 => "00010101",26648 => "10100000",26649 => "11100000",26650 => "11101000",26651 => "11000100",26652 => "00111001",26653 => "10100110",26654 => "11000010",26655 => "00001111",26656 => "11100010",26657 => "01100100",26658 => "10100101",26659 => "01100100",26660 => "00110100",26661 => "00100011",26662 => "00100101",26663 => "00001101",26664 => "00110000",26665 => "11100001",26666 => "01110001",26667 => "11101100",26668 => "01110011",26669 => "00001110",26670 => "00100010",26671 => "11000100",26672 => "01111001",26673 => "01100011",26674 => "01010110",26675 => "00100000",26676 => "01100101",26677 => "01011111",26678 => "00010011",26679 => "11010011",26680 => "00101101",26681 => "01000000",26682 => "01100110",26683 => "00001101",26684 => "11001101",26685 => "11011010",26686 => "01100100",26687 => "11010011",26688 => "11100000",26689 => "01000010",26690 => "10111110",26691 => "11011111",26692 => "10001010",26693 => "01101110",26694 => "10001101",26695 => "10110000",26696 => "00100001",26697 => "01101100",26698 => "10110100",26699 => "10001000",26700 => "01100011",26701 => "01100110",26702 => "11001010",26703 => "00111011",26704 => "00111101",26705 => "11001111",26706 => "10011010",26707 => "11010111",26708 => "11101110",26709 => "11111001",26710 => "01001100",26711 => "10101000",26712 => "11010111",26713 => "01000000",26714 => "11100111",26715 => "01010010",26716 => "00100111",26717 => "01000011",26718 => "10010111",26719 => "11110000",26720 => "01110110",26721 => "11100010",26722 => "10001011",26723 => "01111000",26724 => "01010100",26725 => "00101100",26726 => "01011000",26727 => "00001000",26728 => "01000001",26729 => "01111100",26730 => "10011001",26731 => "01111111",26732 => "01110011",26733 => "10011000",26734 => "01011011",26735 => "00110100",26736 => "00011000",26737 => "11101001",26738 => "10110011",26739 => "11110100",26740 => "11111100",26741 => "01101101",26742 => "00101110",26743 => "00001000",26744 => "10111111",26745 => "00010011",26746 => "01110000",26747 => "11101100",26748 => "00101000",26749 => "00001010",26750 => "01110000",26751 => "10001010",26752 => "10011101",26753 => "10100001",26754 => "01110100",26755 => "00010110",26756 => "11111001",26757 => "01000110",26758 => "01001000",26759 => "11111000",26760 => "10000000",26761 => "10000111",26762 => "01000101",26763 => "01010100",26764 => "11011101",26765 => "01110100",26766 => "01011001",26767 => "11010111",26768 => "10101110",26769 => "10101000",26770 => "10011001",26771 => "01000011",26772 => "00111010",26773 => "11000011",26774 => "01001000",26775 => "00000110",26776 => "01110000",26777 => "11000000",26778 => "01011110",26779 => "00111110",26780 => "00100011",26781 => "10100101",26782 => "11100001",26783 => "10001110",26784 => "01100000",26785 => "01010010",26786 => "00011011",26787 => "11111000",26788 => "01010110",26789 => "01111101",26790 => "11010100",26791 => "11010110",26792 => "10101110",26793 => "10101010",26794 => "11000100",26795 => "00001101",26796 => "00110010",26797 => "01001110",26798 => "11001001",26799 => "10110100",26800 => "10100001",26801 => "11010011",26802 => "01010010",26803 => "10010000",26804 => "11100000",26805 => "01110011",26806 => "11101010",26807 => "10111111",26808 => "11100000",26809 => "00000000",26810 => "01100100",26811 => "10001010",26812 => "01101100",26813 => "00100111",26814 => "10011011",26815 => "00100011",26816 => "00101011",26817 => "10001101",26818 => "11001101",26819 => "01010011",26820 => "00011011",26821 => "01101100",26822 => "01001101",26823 => "01000010",26824 => "11011111",26825 => "10101011",26826 => "01100010",26827 => "01001111",26828 => "01010100",26829 => "01010110",26830 => "00011010",26831 => "01111110",26832 => "11001000",26833 => "10011100",26834 => "11100011",26835 => "00110000",26836 => "01001011",26837 => "00011100",26838 => "10001011",26839 => "11101000",26840 => "11100001",26841 => "11001000",26842 => "00000111",26843 => "11011010",26844 => "00011101",26845 => "00111000",26846 => "10001001",26847 => "01010101",26848 => "11101101",26849 => "00011001",26850 => "01111101",26851 => "00000111",26852 => "11110011",26853 => "10110010",26854 => "00010000",26855 => "00100000",26856 => "11101111",26857 => "00001001",26858 => "11010000",26859 => "01011101",26860 => "10101011",26861 => "11000011",26862 => "10010100",26863 => "00110110",26864 => "11101111",26865 => "01010101",26866 => "00011001",26867 => "01100000",26868 => "01001111",26869 => "11100110",26870 => "10011111",26871 => "11000000",26872 => "11010110",26873 => "00000001",26874 => "10101111",26875 => "00001101",26876 => "11000000",26877 => "11010010",26878 => "10010001",26879 => "00101000",26880 => "00001010",26881 => "10010000",26882 => "10111111",26883 => "11100001",26884 => "00100001",26885 => "11101000",26886 => "10011100",26887 => "11100000",26888 => "10001111",26889 => "01001001",26890 => "11100010",26891 => "11110100",26892 => "10011110",26893 => "11110111",26894 => "00110010",26895 => "00010010",26896 => "00101100",26897 => "11111010",26898 => "00010101",26899 => "11110001",26900 => "00001001",26901 => "11110010",26902 => "10101010",26903 => "01101001",26904 => "01000100",26905 => "01111101",26906 => "11110001",26907 => "00100001",26908 => "10101010",26909 => "10000100",26910 => "11111100",26911 => "10010000",26912 => "01010111",26913 => "10001010",26914 => "01001111",26915 => "10101101",26916 => "01101101",26917 => "01100011",26918 => "01111100",26919 => "10101101",26920 => "10011111",26921 => "11001101",26922 => "10010101",26923 => "01101101",26924 => "10010001",26925 => "00100001",26926 => "11011100",26927 => "01001100",26928 => "00110011",26929 => "11110111",26930 => "10000100",26931 => "11101011",26932 => "11110011",26933 => "11110110",26934 => "01110010",26935 => "10010000",26936 => "01100110",26937 => "01111001",26938 => "11111110",26939 => "00100011",26940 => "10100001",26941 => "10000111",26942 => "01100100",26943 => "10001001",26944 => "00010001",26945 => "10000100",26946 => "10000001",26947 => "01111011",26948 => "11001011",26949 => "10101111",26950 => "10111001",26951 => "00001100",26952 => "00010111",26953 => "01011010",26954 => "11000000",26955 => "11011110",26956 => "11011100",26957 => "00110111",26958 => "00101100",26959 => "10110100",26960 => "10010100",26961 => "00100001",26962 => "11111111",26963 => "01111011",26964 => "11001000",26965 => "11001110",26966 => "01100101",26967 => "00110001",26968 => "10011010",26969 => "10011001",26970 => "11100111",26971 => "11011101",26972 => "00110010",26973 => "00011101",26974 => "01010011",26975 => "11001001",26976 => "11111110",26977 => "10011111",26978 => "11111000",26979 => "00100000",26980 => "01001000",26981 => "11100000",26982 => "01111110",26983 => "01100000",26984 => "00001111",26985 => "10010001",26986 => "11011001",26987 => "01101001",26988 => "11100111",26989 => "00000001",26990 => "10101110",26991 => "10010101",26992 => "00000110",26993 => "01010110",26994 => "01001101",26995 => "10001110",26996 => "00100101",26997 => "01111110",26998 => "01111010",26999 => "11001111",27000 => "00011111",27001 => "11011111",27002 => "11010111",27003 => "01011111",27004 => "10110000",27005 => "11001000",27006 => "00000110",27007 => "01011000",27008 => "10010010",27009 => "10000101",27010 => "01101000",27011 => "01000011",27012 => "10110011",27013 => "11010111",27014 => "10000111",27015 => "11011010",27016 => "10101001",27017 => "10110001",27018 => "01100100",27019 => "11101101",27020 => "01101111",27021 => "01011001",27022 => "11001001",27023 => "11101010",27024 => "00111110",27025 => "10110111",27026 => "10011000",27027 => "10100110",27028 => "11100010",27029 => "01101000",27030 => "11110111",27031 => "11110110",27032 => "11100001",27033 => "10110111",27034 => "10100011",27035 => "01100101",27036 => "01100111",27037 => "01001010",27038 => "00101001",27039 => "01101000",27040 => "10100110",27041 => "01100010",27042 => "01101011",27043 => "11011110",27044 => "00001100",27045 => "11000101",27046 => "01100011",27047 => "01001100",27048 => "01101100",27049 => "11100000",27050 => "10001010",27051 => "00001000",27052 => "10100111",27053 => "01110111",27054 => "01110101",27055 => "11100101",27056 => "00011000",27057 => "00111000",27058 => "01011011",27059 => "01110011",27060 => "01101011",27061 => "11111100",27062 => "01000110",27063 => "00110001",27064 => "00001100",27065 => "00010110",27066 => "10011000",27067 => "00000110",27068 => "00001001",27069 => "10110100",27070 => "11010000",27071 => "10011110",27072 => "01000100",27073 => "01000011",27074 => "10110011",27075 => "10001000",27076 => "10101111",27077 => "11100111",27078 => "00110100",27079 => "11111110",27080 => "10000011",27081 => "00111100",27082 => "00000101",27083 => "01100001",27084 => "00110101",27085 => "11001111",27086 => "00000011",27087 => "00000001",27088 => "11110100",27089 => "00001011",27090 => "01010000",27091 => "10110110",27092 => "01101011",27093 => "00001111",27094 => "00001011",27095 => "01010000",27096 => "11110110",27097 => "00111110",27098 => "00001010",27099 => "00111000",27100 => "11111111",27101 => "01011101",27102 => "00111100",27103 => "00100100",27104 => "11010010",27105 => "11010001",27106 => "10100110",27107 => "10000000",27108 => "11010100",27109 => "01000010",27110 => "10000101",27111 => "10001010",27112 => "11111010",27113 => "00111011",27114 => "10011001",27115 => "00011001",27116 => "10010110",27117 => "10101000",27118 => "00111000",27119 => "10010111",27120 => "00011010",27121 => "11001101",27122 => "10001010",27123 => "00011110",27124 => "01111111",27125 => "11101000",27126 => "01110110",27127 => "00111111",27128 => "01000111",27129 => "11011111",27130 => "11100001",27131 => "11010011",27132 => "01010000",27133 => "11010000",27134 => "00110010",27135 => "10100000",27136 => "01000111",27137 => "10010101",27138 => "11001100",27139 => "01100110",27140 => "10001111",27141 => "10011010",27142 => "10110100",27143 => "11011011",27144 => "00011111",27145 => "11101001",27146 => "11110000",27147 => "01011001",27148 => "11101001",27149 => "01110101",27150 => "10011010",27151 => "10100100",27152 => "10101100",27153 => "01111110",27154 => "10011000",27155 => "10100010",27156 => "00100001",27157 => "10101111",27158 => "01100011",27159 => "01011010",27160 => "10000100",27161 => "11000111",27162 => "11010101",27163 => "10110100",27164 => "11110110",27165 => "10111100",27166 => "01001100",27167 => "10010000",27168 => "00111000",27169 => "00101111",27170 => "00000110",27171 => "01000000",27172 => "00111100",27173 => "00110011",27174 => "11111000",27175 => "10011000",27176 => "11001011",27177 => "00011101",27178 => "11001100",27179 => "11101001",27180 => "00100110",27181 => "01010100",27182 => "00100011",27183 => "10101110",27184 => "01111111",27185 => "00101101",27186 => "01011010",27187 => "01100000",27188 => "10110101",27189 => "11011011",27190 => "01000011",27191 => "10011110",27192 => "01001010",27193 => "10111011",27194 => "11111001",27195 => "10001110",27196 => "10011111",27197 => "00000110",27198 => "10001010",27199 => "11101111",27200 => "11001001",27201 => "11111000",27202 => "10100110",27203 => "00110110",27204 => "10010011",27205 => "10110101",27206 => "11011000",27207 => "10111000",27208 => "00011000",27209 => "10101100",27210 => "00011110",27211 => "10001111",27212 => "01111100",27213 => "10100110",27214 => "01001100",27215 => "00011101",27216 => "01001000",27217 => "11011000",27218 => "00001000",27219 => "10010010",27220 => "10011010",27221 => "00001001",27222 => "10000100",27223 => "01000100",27224 => "01001110",27225 => "10010010",27226 => "00111101",27227 => "00111101",27228 => "00011111",27229 => "10100110",27230 => "10011011",27231 => "01111100",27232 => "00100101",27233 => "01111000",27234 => "00110000",27235 => "00000011",27236 => "10010011",27237 => "00110100",27238 => "01001010",27239 => "11110001",27240 => "01010010",27241 => "00011100",27242 => "00111011",27243 => "10110000",27244 => "00000010",27245 => "11111010",27246 => "00101101",27247 => "10100101",27248 => "01110111",27249 => "10100110",27250 => "10001000",27251 => "01110110",27252 => "01010100",27253 => "10001111",27254 => "10000001",27255 => "01001010",27256 => "10101001",27257 => "00010010",27258 => "10001111",27259 => "01100010",27260 => "01000101",27261 => "10001010",27262 => "01010101",27263 => "00011001",27264 => "11111000",27265 => "00011110",27266 => "00110100",27267 => "01001011",27268 => "11101110",27269 => "10001011",27270 => "00111100",27271 => "01111000",27272 => "00100100",27273 => "10101111",27274 => "11101001",27275 => "11011011",27276 => "10010011",27277 => "10101110",27278 => "10001100",27279 => "00001010",27280 => "11011110",27281 => "10011101",27282 => "00101011",27283 => "00100000",27284 => "11101101",27285 => "11000000",27286 => "01110101",27287 => "01001011",27288 => "10001001",27289 => "00100010",27290 => "11110010",27291 => "11110000",27292 => "00111010",27293 => "10011101",27294 => "11001010",27295 => "11010110",27296 => "11100001",27297 => "10000100",27298 => "11010101",27299 => "11001011",27300 => "00101010",27301 => "10110011",27302 => "01100001",27303 => "11110001",27304 => "11011111",27305 => "00000001",27306 => "01101100",27307 => "11010001",27308 => "11110010",27309 => "10100101",27310 => "00010111",27311 => "00111010",27312 => "01110101",27313 => "10011110",27314 => "01100111",27315 => "00111000",27316 => "10011101",27317 => "11001110",27318 => "10001101",27319 => "11100011",27320 => "00010000",27321 => "00100011",27322 => "01110001",27323 => "01111100",27324 => "01001101",27325 => "10110100",27326 => "10011110",27327 => "10010000",27328 => "01010011",27329 => "01110001",27330 => "10001011",27331 => "11111001",27332 => "01000110",27333 => "00011001",27334 => "11110111",27335 => "01111111",27336 => "10111001",27337 => "00000110",27338 => "10001011",27339 => "00010111",27340 => "11011101",27341 => "11101110",27342 => "01011101",27343 => "10001001",27344 => "00011110",27345 => "01111110",27346 => "10000001",27347 => "01101111",27348 => "11100010",27349 => "11010100",27350 => "10110000",27351 => "01011111",27352 => "11000111",27353 => "10101011",27354 => "10000100",27355 => "01101011",27356 => "00111001",27357 => "11011011",27358 => "01011000",27359 => "10111100",27360 => "01010111",27361 => "00000011",27362 => "10010110",27363 => "01111001",27364 => "01110001",27365 => "01000011",27366 => "01111000",27367 => "01100101",27368 => "10101111",27369 => "00110011",27370 => "01111100",27371 => "00110110",27372 => "01101101",27373 => "10010011",27374 => "00000110",27375 => "10011111",27376 => "01100101",27377 => "10000010",27378 => "00001110",27379 => "10101101",27380 => "00111001",27381 => "11111010",27382 => "01000010",27383 => "00010001",27384 => "01111000",27385 => "00100011",27386 => "11111010",27387 => "11101101",27388 => "10011001",27389 => "01101110",27390 => "10101101",27391 => "10011000",27392 => "10000001",27393 => "01101000",27394 => "11110110",27395 => "10100110",27396 => "10010110",27397 => "01101011",27398 => "11110000",27399 => "10111110",27400 => "10000001",27401 => "10010100",27402 => "01001011",27403 => "10001100",27404 => "10100001",27405 => "01101010",27406 => "01110100",27407 => "10000001",27408 => "10001111",27409 => "00100110",27410 => "00110010",27411 => "01110000",27412 => "01001100",27413 => "01101110",27414 => "11101010",27415 => "00001000",27416 => "11111101",27417 => "01010100",27418 => "11100000",27419 => "10001110",27420 => "11110000",27421 => "01011010",27422 => "01101111",27423 => "01100011",27424 => "10111011",27425 => "11101111",27426 => "11111000",27427 => "10011110",27428 => "00101111",27429 => "00011100",27430 => "00110010",27431 => "11000110",27432 => "11011111",27433 => "11111010",27434 => "01101011",27435 => "01001110",27436 => "11110011",27437 => "11100011",27438 => "10011101",27439 => "01001010",27440 => "00000000",27441 => "00100111",27442 => "11000000",27443 => "01111000",27444 => "10110101",27445 => "01110001",27446 => "01010100",27447 => "00111001",27448 => "10100100",27449 => "10101010",27450 => "10001010",27451 => "00011001",27452 => "11100100",27453 => "00110111",27454 => "01110010",27455 => "10001111",27456 => "01111110",27457 => "00000110",27458 => "11101101",27459 => "00111000",27460 => "11110100",27461 => "01110001",27462 => "10010011",27463 => "00111100",27464 => "00100101",27465 => "00000100",27466 => "10100010",27467 => "10110110",27468 => "00101111",27469 => "11110011",27470 => "01000100",27471 => "01101100",27472 => "10001000",27473 => "11001000",27474 => "01000010",27475 => "00110101",27476 => "11011010",27477 => "10001001",27478 => "00100101",27479 => "10001011",27480 => "11101101",27481 => "11101111",27482 => "11101100",27483 => "11101001",27484 => "00111001",27485 => "01000100",27486 => "01000010",27487 => "00110111",27488 => "00111000",27489 => "11100010",27490 => "01010000",27491 => "00011010",27492 => "01001000",27493 => "00111101",27494 => "01110100",27495 => "11111001",27496 => "11110001",27497 => "11101011",27498 => "11110110",27499 => "01010101",27500 => "00011000",27501 => "01010001",27502 => "11001010",27503 => "01100000",27504 => "00110000",27505 => "10100011",27506 => "11001011",27507 => "11001100",27508 => "00001001",27509 => "10111101",27510 => "00000011",27511 => "10100010",27512 => "10011000",27513 => "00000111",27514 => "10101010",27515 => "01011101",27516 => "11001011",27517 => "01101001",27518 => "11110000",27519 => "01001011",27520 => "00010001",27521 => "01000001",27522 => "01010001",27523 => "00010001",27524 => "00110101",27525 => "01000100",27526 => "00011001",27527 => "00110111",27528 => "11101100",27529 => "00000011",27530 => "00110001",27531 => "00111010",27532 => "01000010",27533 => "01001011",27534 => "10001110",27535 => "01001110",27536 => "10001010",27537 => "10110110",27538 => "00011100",27539 => "10001100",27540 => "01011101",27541 => "10011000",27542 => "00100101",27543 => "00111001",27544 => "00011100",27545 => "10001100",27546 => "10010111",27547 => "01010100",27548 => "11110000",27549 => "11111011",27550 => "01101101",27551 => "00010100",27552 => "10111110",27553 => "10100110",27554 => "10011001",27555 => "11011001",27556 => "10100000",27557 => "00111100",27558 => "00000110",27559 => "10011010",27560 => "11110010",27561 => "11001011",27562 => "00111111",27563 => "00111011",27564 => "00010010",27565 => "10111100",27566 => "00010010",27567 => "11100011",27568 => "00001100",27569 => "10010000",27570 => "00001010",27571 => "11111101",27572 => "11010100",27573 => "00001101",27574 => "11011010",27575 => "11011011",27576 => "10110011",27577 => "10001001",27578 => "10101001",27579 => "10010111",27580 => "00100101",27581 => "01001111",27582 => "11000110",27583 => "11110001",27584 => "11001001",27585 => "10100011",27586 => "01100100",27587 => "00100011",27588 => "00100001",27589 => "11010000",27590 => "01111101",27591 => "00001100",27592 => "11110011",27593 => "11101101",27594 => "10100011",27595 => "10100001",27596 => "10111001",27597 => "10111011",27598 => "11111100",27599 => "11101100",27600 => "11011000",27601 => "01110101",27602 => "00000111",27603 => "00010110",27604 => "00100111",27605 => "01011110",27606 => "00100001",27607 => "10011100",27608 => "10001100",27609 => "01011100",27610 => "01010100",27611 => "11000000",27612 => "01100111",27613 => "10010101",27614 => "10100101",27615 => "00010011",27616 => "00000101",27617 => "01110111",27618 => "01111100",27619 => "11100100",27620 => "10110010",27621 => "11100101",27622 => "01011001",27623 => "10100010",27624 => "01100010",27625 => "11110000",27626 => "11101001",27627 => "00010010",27628 => "10111000",27629 => "00101101",27630 => "00101110",27631 => "00110000",27632 => "00010101",27633 => "11111010",27634 => "11001010",27635 => "10011000",27636 => "01011011",27637 => "01001010",27638 => "11010010",27639 => "11100101",27640 => "01000101",27641 => "10001111",27642 => "01001010",27643 => "11000011",27644 => "10111000",27645 => "11111001",27646 => "01010000",27647 => "01111111",27648 => "00001001",27649 => "11100110",27650 => "11111111",27651 => "11101111",27652 => "01100100",27653 => "11111011",27654 => "10011111",27655 => "00110011",27656 => "00100111",27657 => "00110011",27658 => "11010101",27659 => "11101010",27660 => "10100011",27661 => "10111011",27662 => "01100110",27663 => "10010001",27664 => "00011011",27665 => "11011110",27666 => "00010001",27667 => "01011111",27668 => "11101101",27669 => "00110111",27670 => "00001110",27671 => "01011001",27672 => "10011110",27673 => "11110100",27674 => "01001111",27675 => "00101001",27676 => "11111001",27677 => "10101011",27678 => "10000010",27679 => "00101100",27680 => "01100010",27681 => "11010110",27682 => "00111011",27683 => "10011110",27684 => "01011010",27685 => "00100011",27686 => "10111101",27687 => "00111101",27688 => "11011100",27689 => "11011010",27690 => "00001100",27691 => "11110100",27692 => "10001000",27693 => "11110000",27694 => "01001101",27695 => "10011100",27696 => "10100010",27697 => "00100011",27698 => "01011000",27699 => "01010010",27700 => "01100000",27701 => "01000010",27702 => "10110111",27703 => "10000011",27704 => "10011111",27705 => "11001111",27706 => "11111011",27707 => "00010100",27708 => "00110011",27709 => "00000101",27710 => "11001000",27711 => "11011100",27712 => "01100110",27713 => "11101110",27714 => "10101100",27715 => "00111011",27716 => "10001110",27717 => "11110101",27718 => "00110000",27719 => "11011101",27720 => "10101110",27721 => "10110111",27722 => "11010001",27723 => "11001110",27724 => "00110010",27725 => "11111011",27726 => "10010000",27727 => "01000011",27728 => "01110010",27729 => "00011000",27730 => "01010111",27731 => "00001011",27732 => "11110011",27733 => "00110000",27734 => "01110001",27735 => "01010100",27736 => "10001100",27737 => "11001001",27738 => "00001100",27739 => "00010100",27740 => "01000110",27741 => "00101000",27742 => "10100110",27743 => "10100100",27744 => "11110111",27745 => "01000100",27746 => "11001101",27747 => "10000111",27748 => "00011111",27749 => "00101010",27750 => "10000101",27751 => "00111111",27752 => "01000001",27753 => "10101011",27754 => "10011110",27755 => "01101011",27756 => "01110110",27757 => "10011010",27758 => "01100100",27759 => "00011000",27760 => "00110100",27761 => "00110001",27762 => "00111101",27763 => "00111100",27764 => "00100010",27765 => "01001001",27766 => "11101100",27767 => "01001001",27768 => "10011100",27769 => "00010100",27770 => "01110011",27771 => "01100000",27772 => "01110100",27773 => "00110101",27774 => "00011010",27775 => "01100011",27776 => "11010000",27777 => "10111101",27778 => "11111011",27779 => "01011111",27780 => "01101000",27781 => "11000100",27782 => "01000001",27783 => "11100010",27784 => "10111010",27785 => "00100101",27786 => "11100000",27787 => "11011001",27788 => "00101110",27789 => "11111010",27790 => "00101110",27791 => "11001110",27792 => "00000100",27793 => "11000010",27794 => "00111101",27795 => "10101010",27796 => "01101000",27797 => "00001111",27798 => "11001111",27799 => "11101111",27800 => "11001110",27801 => "10111101",27802 => "11101110",27803 => "10000011",27804 => "11000101",27805 => "01100110",27806 => "01100001",27807 => "11010001",27808 => "01101100",27809 => "00100001",27810 => "11111011",27811 => "00011011",27812 => "01010011",27813 => "00101100",27814 => "11001110",27815 => "10111010",27816 => "11001111",27817 => "11000011",27818 => "11000111",27819 => "01100001",27820 => "11111111",27821 => "01010011",27822 => "00111101",27823 => "10110100",27824 => "01010111",27825 => "00101111",27826 => "10001010",27827 => "10000100",27828 => "01110111",27829 => "10101111",27830 => "00011111",27831 => "00111011",27832 => "01001010",27833 => "10101000",27834 => "10011010",27835 => "11101110",27836 => "11010100",27837 => "00100100",27838 => "10001100",27839 => "00010010",27840 => "11001001",27841 => "00110011",27842 => "01101000",27843 => "11010001",27844 => "11100110",27845 => "01100010",27846 => "10001001",27847 => "11100110",27848 => "10001011",27849 => "11010110",27850 => "01110011",27851 => "11111000",27852 => "11000010",27853 => "11100010",27854 => "00100001",27855 => "01010010",27856 => "01111101",27857 => "01100111",27858 => "11010010",27859 => "11100100",27860 => "01101100",27861 => "00010001",27862 => "00101111",27863 => "00001101",27864 => "01100110",27865 => "00101010",27866 => "10010001",27867 => "10001011",27868 => "00011000",27869 => "11111100",27870 => "11100101",27871 => "11110110",27872 => "10101110",27873 => "00000011",27874 => "00011000",27875 => "00110110",27876 => "11000010",27877 => "01100010",27878 => "11111010",27879 => "01110110",27880 => "11100100",27881 => "11111100",27882 => "01101000",27883 => "00110100",27884 => "01110000",27885 => "10010111",27886 => "11110111",27887 => "10100001",27888 => "10010010",27889 => "10001111",27890 => "01111101",27891 => "00111011",27892 => "11010010",27893 => "01110000",27894 => "01000110",27895 => "11101001",27896 => "10100101",27897 => "01101000",27898 => "00110001",27899 => "00001011",27900 => "11101010",27901 => "11111010",27902 => "10101100",27903 => "11111011",27904 => "11001111",27905 => "10001101",27906 => "10001011",27907 => "00000100",27908 => "00110001",27909 => "11110010",27910 => "10010000",27911 => "11010110",27912 => "10010110",27913 => "10001100",27914 => "00001100",27915 => "10101100",27916 => "01001011",27917 => "10111110",27918 => "01110111",27919 => "10000000",27920 => "01001010",27921 => "00011110",27922 => "00110001",27923 => "11001010",27924 => "00101011",27925 => "00110101",27926 => "01100111",27927 => "01011001",27928 => "10100111",27929 => "00100000",27930 => "10001010",27931 => "01111110",27932 => "10001101",27933 => "00110000",27934 => "01010000",27935 => "11000110",27936 => "00101001",27937 => "10001110",27938 => "00101011",27939 => "00110010",27940 => "11000101",27941 => "10110100",27942 => "00011110",27943 => "10001110",27944 => "10110000",27945 => "01000000",27946 => "00010010",27947 => "00100100",27948 => "11111000",27949 => "11100000",27950 => "10110100",27951 => "11110111",27952 => "01100010",27953 => "00111001",27954 => "10100011",27955 => "00000010",27956 => "11011001",27957 => "10010011",27958 => "01011011",27959 => "01010110",27960 => "01011010",27961 => "11001000",27962 => "01000011",27963 => "10101111",27964 => "10110111",27965 => "11110001",27966 => "11110111",27967 => "11111001",27968 => "01011011",27969 => "11010110",27970 => "11000101",27971 => "00011011",27972 => "01011101",27973 => "11110000",27974 => "10001011",27975 => "00000001",27976 => "00101001",27977 => "01111011",27978 => "10011110",27979 => "00001110",27980 => "00011101",27981 => "00001000",27982 => "11000001",27983 => "11110110",27984 => "01101111",27985 => "11001111",27986 => "11001010",27987 => "11001101",27988 => "01010010",27989 => "10100100",27990 => "00000010",27991 => "01011100",27992 => "10111001",27993 => "10110011",27994 => "00110111",27995 => "01000010",27996 => "11101010",27997 => "00001000",27998 => "10010000",27999 => "11101000",28000 => "11100011",28001 => "10111001",28002 => "11101110",28003 => "01010100",28004 => "10001111",28005 => "10010011",28006 => "01000001",28007 => "00011101",28008 => "10000100",28009 => "00001100",28010 => "10010001",28011 => "01111011",28012 => "01010000",28013 => "11110110",28014 => "00010111",28015 => "01100001",28016 => "11000100",28017 => "01000101",28018 => "00010011",28019 => "10101100",28020 => "00010111",28021 => "00101011",28022 => "01010001",28023 => "10011001",28024 => "00110011",28025 => "11110101",28026 => "10100000",28027 => "10110100",28028 => "00101111",28029 => "01100000",28030 => "01011000",28031 => "10100010",28032 => "10001010",28033 => "10100100",28034 => "11111000",28035 => "01110010",28036 => "00101111",28037 => "00001101",28038 => "11001010",28039 => "11111100",28040 => "00000110",28041 => "10111000",28042 => "10010010",28043 => "00010011",28044 => "10101011",28045 => "01010110",28046 => "00100101",28047 => "00101010",28048 => "11111011",28049 => "01100000",28050 => "01010010",28051 => "00001101",28052 => "01110000",28053 => "10110000",28054 => "00010111",28055 => "11100010",28056 => "10100000",28057 => "10100011",28058 => "11111000",28059 => "00000100",28060 => "11001100",28061 => "01011011",28062 => "10010101",28063 => "11100111",28064 => "00010000",28065 => "11101001",28066 => "11011110",28067 => "00001100",28068 => "10101100",28069 => "00010010",28070 => "10011111",28071 => "11001010",28072 => "01110001",28073 => "11100100",28074 => "00010111",28075 => "01010110",28076 => "01101110",28077 => "01100001",28078 => "10001000",28079 => "11001001",28080 => "10010001",28081 => "01010101",28082 => "10011101",28083 => "01101011",28084 => "10110010",28085 => "00110101",28086 => "10110001",28087 => "01011000",28088 => "00010010",28089 => "01010010",28090 => "00100010",28091 => "11100110",28092 => "01001000",28093 => "11011001",28094 => "10101101",28095 => "00001011",28096 => "00000100",28097 => "10000111",28098 => "10001111",28099 => "01011001",28100 => "01111101",28101 => "00010001",28102 => "01001011",28103 => "00100001",28104 => "01111111",28105 => "01001110",28106 => "01100100",28107 => "11111001",28108 => "00000110",28109 => "10110001",28110 => "01011111",28111 => "00011110",28112 => "01010101",28113 => "10110100",28114 => "00110011",28115 => "11000010",28116 => "01111101",28117 => "11101011",28118 => "01000100",28119 => "01110111",28120 => "00101001",28121 => "01100110",28122 => "00100110",28123 => "11000110",28124 => "11010001",28125 => "10010011",28126 => "10011100",28127 => "01001100",28128 => "11100001",28129 => "01101011",28130 => "11100001",28131 => "00010001",28132 => "00110011",28133 => "11011110",28134 => "10101010",28135 => "00111011",28136 => "10111000",28137 => "00101010",28138 => "10110100",28139 => "11011111",28140 => "00011100",28141 => "11101100",28142 => "01100110",28143 => "11001101",28144 => "01001111",28145 => "10110101",28146 => "01011001",28147 => "00010101",28148 => "10000001",28149 => "00011000",28150 => "00101001",28151 => "11010010",28152 => "01011011",28153 => "11110101",28154 => "11100000",28155 => "00010111",28156 => "11000101",28157 => "11011111",28158 => "10010011",28159 => "00100000",28160 => "00110001",28161 => "11111001",28162 => "10001000",28163 => "11111110",28164 => "00101001",28165 => "10101100",28166 => "11101100",28167 => "10101100",28168 => "01110000",28169 => "11011011",28170 => "10111111",28171 => "10011110",28172 => "10101110",28173 => "10100110",28174 => "01101010",28175 => "11101000",28176 => "10110011",28177 => "01101111",28178 => "10100000",28179 => "11100001",28180 => "00111000",28181 => "10011110",28182 => "00111000",28183 => "10011111",28184 => "00100100",28185 => "00110110",28186 => "10011100",28187 => "00110010",28188 => "00011111",28189 => "10001110",28190 => "10111100",28191 => "00100111",28192 => "01111101",28193 => "11101111",28194 => "10101001",28195 => "10011111",28196 => "00110000",28197 => "10000001",28198 => "11010110",28199 => "01001000",28200 => "10100111",28201 => "01001001",28202 => "01011011",28203 => "11011111",28204 => "00010111",28205 => "10111101",28206 => "00111011",28207 => "11010111",28208 => "01001000",28209 => "11100001",28210 => "10101101",28211 => "10110010",28212 => "01010001",28213 => "00001001",28214 => "00111001",28215 => "10001110",28216 => "01110001",28217 => "10011100",28218 => "11110011",28219 => "01001011",28220 => "10111100",28221 => "10001001",28222 => "01010000",28223 => "10101100",28224 => "00101000",28225 => "10001100",28226 => "00111011",28227 => "11101001",28228 => "01101110",28229 => "11110111",28230 => "00000000",28231 => "01011101",28232 => "10011111",28233 => "11001010",28234 => "01011001",28235 => "00101110",28236 => "00001001",28237 => "10001111",28238 => "11111011",28239 => "10010100",28240 => "11010101",28241 => "00110101",28242 => "00001111",28243 => "11100101",28244 => "00001111",28245 => "01110010",28246 => "01000110",28247 => "10111100",28248 => "11111010",28249 => "00000101",28250 => "11101011",28251 => "01110110",28252 => "00110001",28253 => "11100100",28254 => "01111111",28255 => "11010000",28256 => "00110001",28257 => "11000100",28258 => "11111000",28259 => "11011101",28260 => "01001010",28261 => "10110000",28262 => "00110011",28263 => "01110000",28264 => "00100000",28265 => "10110111",28266 => "00010111",28267 => "00000101",28268 => "10011001",28269 => "10110011",28270 => "10100011",28271 => "11100001",28272 => "10111001",28273 => "00111010",28274 => "10101111",28275 => "11010110",28276 => "10110000",28277 => "11000010",28278 => "01011110",28279 => "00101111",28280 => "00111000",28281 => "10010011",28282 => "00000100",28283 => "11001101",28284 => "01001111",28285 => "11111110",28286 => "11110111",28287 => "01110001",28288 => "10100001",28289 => "00100100",28290 => "11100100",28291 => "11110100",28292 => "10000001",28293 => "00010001",28294 => "11010100",28295 => "10111010",28296 => "11010011",28297 => "11011000",28298 => "10001110",28299 => "11011111",28300 => "00001001",28301 => "11110001",28302 => "00011111",28303 => "01011010",28304 => "01111100",28305 => "01010011",28306 => "01100010",28307 => "10011110",28308 => "10010010",28309 => "10111101",28310 => "00100101",28311 => "00110011",28312 => "10011000",28313 => "00111001",28314 => "00100100",28315 => "11001000",28316 => "11101011",28317 => "11011101",28318 => "00011110",28319 => "01101011",28320 => "10011001",28321 => "00001111",28322 => "11110101",28323 => "00110110",28324 => "11001100",28325 => "01011011",28326 => "00101111",28327 => "01110001",28328 => "00100110",28329 => "00111010",28330 => "11111111",28331 => "11101111",28332 => "00011011",28333 => "00100001",28334 => "10110101",28335 => "01011101",28336 => "01011010",28337 => "10100011",28338 => "00110011",28339 => "01011000",28340 => "10110010",28341 => "10111010",28342 => "01010110",28343 => "10111101",28344 => "01011111",28345 => "00100001",28346 => "10000010",28347 => "01001000",28348 => "01111110",28349 => "11111010",28350 => "00101100",28351 => "01110111",28352 => "11010110",28353 => "01011011",28354 => "01110001",28355 => "10100000",28356 => "11111101",28357 => "00001111",28358 => "10010001",28359 => "01011001",28360 => "00001110",28361 => "10000111",28362 => "00101010",28363 => "00110000",28364 => "11010000",28365 => "01100010",28366 => "11010000",28367 => "10001001",28368 => "11100110",28369 => "11111001",28370 => "11111101",28371 => "00010001",28372 => "11011101",28373 => "11110101",28374 => "11101111",28375 => "01000001",28376 => "11101111",28377 => "10101101",28378 => "11001111",28379 => "00110011",28380 => "11111110",28381 => "10111111",28382 => "11100100",28383 => "00111010",28384 => "01100000",28385 => "01101100",28386 => "11101110",28387 => "01100010",28388 => "11001000",28389 => "11110000",28390 => "10000010",28391 => "00100011",28392 => "00010011",28393 => "01000111",28394 => "10011101",28395 => "11011100",28396 => "00001010",28397 => "01111011",28398 => "11001101",28399 => "01100011",28400 => "11000001",28401 => "00011111",28402 => "11011001",28403 => "00010001",28404 => "01010110",28405 => "10011101",28406 => "11110011",28407 => "01110000",28408 => "01110000",28409 => "00101111",28410 => "00100010",28411 => "10010110",28412 => "00101000",28413 => "10111101",28414 => "01001100",28415 => "01111110",28416 => "00110011",28417 => "10011111",28418 => "01101010",28419 => "10001001",28420 => "01111111",28421 => "00000000",28422 => "10001111",28423 => "10000100",28424 => "10001001",28425 => "10000100",28426 => "10011011",28427 => "11001010",28428 => "01010110",28429 => "10000101",28430 => "10101101",28431 => "01000011",28432 => "10011111",28433 => "11101000",28434 => "11110101",28435 => "00110011",28436 => "01110001",28437 => "10000110",28438 => "10010111",28439 => "10011111",28440 => "11000001",28441 => "01001011",28442 => "11100000",28443 => "01010101",28444 => "11010000",28445 => "11001100",28446 => "01111100",28447 => "01111001",28448 => "10110100",28449 => "10000110",28450 => "00011111",28451 => "01111110",28452 => "11101001",28453 => "10000100",28454 => "11101111",28455 => "11000101",28456 => "11010010",28457 => "00111100",28458 => "00011110",28459 => "00101110",28460 => "01111111",28461 => "01100001",28462 => "10101101",28463 => "01011001",28464 => "00010101",28465 => "11001101",28466 => "01001111",28467 => "10011110",28468 => "00000111",28469 => "01011100",28470 => "00100001",28471 => "11100011",28472 => "00010101",28473 => "01000100",28474 => "00101100",28475 => "00111000",28476 => "00001011",28477 => "10100010",28478 => "11101101",28479 => "01100111",28480 => "10000110",28481 => "10100001",28482 => "11111110",28483 => "00101100",28484 => "00011011",28485 => "10110010",28486 => "11111101",28487 => "00110110",28488 => "00100100",28489 => "10011101",28490 => "01001100",28491 => "00010110",28492 => "10001110",28493 => "00001001",28494 => "00101111",28495 => "01101100",28496 => "11010011",28497 => "00011011",28498 => "00010000",28499 => "01100111",28500 => "00111101",28501 => "01111100",28502 => "10100100",28503 => "01101001",28504 => "11001100",28505 => "11111111",28506 => "00000101",28507 => "10000001",28508 => "00010110",28509 => "00110000",28510 => "00111011",28511 => "10111010",28512 => "00100001",28513 => "11100111",28514 => "11000111",28515 => "01111011",28516 => "01000001",28517 => "00111011",28518 => "01111011",28519 => "10110110",28520 => "10000110",28521 => "11100100",28522 => "00110101",28523 => "01001100",28524 => "00011001",28525 => "11111111",28526 => "00100000",28527 => "00000101",28528 => "01011110",28529 => "01100100",28530 => "00100111",28531 => "01010100",28532 => "01000101",28533 => "00111101",28534 => "11111100",28535 => "11001110",28536 => "11010001",28537 => "10101001",28538 => "00111001",28539 => "11111011",28540 => "01110111",28541 => "00000101",28542 => "00100101",28543 => "01000110",28544 => "01101001",28545 => "00100111",28546 => "10111000",28547 => "10010001",28548 => "01000101",28549 => "11111011",28550 => "11100101",28551 => "01010110",28552 => "01111100",28553 => "11011101",28554 => "11111100",28555 => "11111110",28556 => "10011000",28557 => "01101100",28558 => "11001001",28559 => "01000100",28560 => "01001101",28561 => "00100000",28562 => "10000111",28563 => "11011011",28564 => "01001100",28565 => "10001100",28566 => "10111011",28567 => "10010100",28568 => "01101011",28569 => "11110101",28570 => "00101100",28571 => "10101111",28572 => "10100101",28573 => "11101110",28574 => "00011110",28575 => "10000100",28576 => "00100010",28577 => "00001101",28578 => "00010101",28579 => "01001111",28580 => "00001101",28581 => "10011100",28582 => "10011000",28583 => "11100010",28584 => "01011101",28585 => "01110000",28586 => "11000000",28587 => "00110101",28588 => "10010010",28589 => "10011100",28590 => "11101010",28591 => "01111100",28592 => "11000100",28593 => "10100011",28594 => "11001000",28595 => "10111101",28596 => "01111111",28597 => "11111100",28598 => "10111001",28599 => "10111101",28600 => "10100001",28601 => "11001101",28602 => "11101001",28603 => "11110001",28604 => "01110101",28605 => "11011000",28606 => "11010001",28607 => "11001011",28608 => "00100000",28609 => "00111010",28610 => "00011110",28611 => "01111011",28612 => "00000101",28613 => "11000000",28614 => "11000111",28615 => "00101110",28616 => "00111001",28617 => "01100011",28618 => "11000011",28619 => "10111110",28620 => "11100010",28621 => "01100011",28622 => "11010000",28623 => "01100000",28624 => "11101000",28625 => "10100101",28626 => "10111111",28627 => "10010000",28628 => "11100000",28629 => "11101000",28630 => "01100010",28631 => "00100011",28632 => "11000101",28633 => "11010010",28634 => "01010101",28635 => "11100010",28636 => "01001010",28637 => "11010011",28638 => "00111111",28639 => "01111110",28640 => "00101010",28641 => "01000111",28642 => "11111101",28643 => "00111111",28644 => "00011000",28645 => "10010111",28646 => "10001001",28647 => "00011000",28648 => "01101110",28649 => "01001000",28650 => "01010100",28651 => "00010101",28652 => "01000010",28653 => "10000000",28654 => "10000110",28655 => "01110010",28656 => "10110001",28657 => "01100001",28658 => "00000101",28659 => "11010100",28660 => "10110100",28661 => "11100100",28662 => "10101110",28663 => "01111010",28664 => "00000001",28665 => "11001101",28666 => "00011000",28667 => "00001100",28668 => "11011000",28669 => "01110101",28670 => "11000111",28671 => "11111010",28672 => "10110100",28673 => "00000000",28674 => "00011100",28675 => "01000000",28676 => "00001110",28677 => "10100000",28678 => "01111011",28679 => "10110001",28680 => "11010010",28681 => "00001000",28682 => "11011101",28683 => "01001101",28684 => "11101001",28685 => "01011011",28686 => "10111000",28687 => "10011001",28688 => "00010010",28689 => "01110100",28690 => "01110010",28691 => "01011010",28692 => "00111101",28693 => "10010110",28694 => "10101011",28695 => "11011110",28696 => "01011011",28697 => "01000100",28698 => "01010010",28699 => "00011010",28700 => "11001110",28701 => "01000110",28702 => "11110000",28703 => "11110001",28704 => "01101111",28705 => "01100110",28706 => "00010010",28707 => "10001011",28708 => "10001111",28709 => "00011011",28710 => "11011101",28711 => "10000111",28712 => "01100111",28713 => "01010000",28714 => "01001001",28715 => "00101011",28716 => "01011010",28717 => "10010010",28718 => "00001000",28719 => "00000011",28720 => "11010000",28721 => "11001001",28722 => "01111101",28723 => "00010011",28724 => "01100000",28725 => "00101111",28726 => "10110100",28727 => "11100101",28728 => "10011111",28729 => "11011011",28730 => "11001101",28731 => "01000000",28732 => "00100101",28733 => "01001011",28734 => "00000110",28735 => "10000110",28736 => "10001001",28737 => "11010010",28738 => "01001011",28739 => "11011100",28740 => "11001101",28741 => "11111110",28742 => "00110111",28743 => "10010111",28744 => "01011111",28745 => "11010111",28746 => "10011111",28747 => "10111000",28748 => "00001001",28749 => "01100011",28750 => "00111100",28751 => "10011111",28752 => "01000001",28753 => "01000001",28754 => "10011001",28755 => "10000100",28756 => "11110110",28757 => "00110111",28758 => "01010100",28759 => "11101011",28760 => "01110111",28761 => "11111000",28762 => "11101010",28763 => "00101101",28764 => "11110001",28765 => "01011000",28766 => "10100011",28767 => "10110100",28768 => "00000110",28769 => "01001001",28770 => "11001110",28771 => "00101011",28772 => "10010110",28773 => "00111101",28774 => "11100010",28775 => "01110100",28776 => "00111011",28777 => "01010001",28778 => "01001100",28779 => "00010000",28780 => "00011101",28781 => "01000110",28782 => "01101110",28783 => "00001111",28784 => "10001010",28785 => "10010001",28786 => "11010000",28787 => "10011111",28788 => "01101110",28789 => "10101110",28790 => "10001000",28791 => "11011010",28792 => "00110011",28793 => "01000101",28794 => "01101001",28795 => "10001000",28796 => "00111011",28797 => "11110010",28798 => "10001010",28799 => "00010100",28800 => "01011010",28801 => "01001010",28802 => "11101110",28803 => "00101010",28804 => "11100100",28805 => "01101000",28806 => "01011101",28807 => "10111101",28808 => "00100110",28809 => "01100010",28810 => "10100000",28811 => "11001100",28812 => "11111110",28813 => "01000100",28814 => "10010011",28815 => "01010100",28816 => "01011010",28817 => "10110010",28818 => "11001101",28819 => "01010101",28820 => "11000111",28821 => "10100101",28822 => "01001111",28823 => "01101001",28824 => "10101100",28825 => "00001001",28826 => "10111010",28827 => "10101100",28828 => "10011100",28829 => "11110100",28830 => "10001100",28831 => "10111000",28832 => "11111100",28833 => "00000110",28834 => "10001111",28835 => "01110101",28836 => "10001001",28837 => "10100111",28838 => "01100111",28839 => "11001001",28840 => "00000001",28841 => "11110110",28842 => "00000010",28843 => "10100001",28844 => "01111010",28845 => "01011010",28846 => "00111111",28847 => "11001011",28848 => "01011011",28849 => "00110010",28850 => "10010011",28851 => "00100101",28852 => "11111010",28853 => "11101000",28854 => "01111110",28855 => "11110011",28856 => "00010001",28857 => "01101101",28858 => "01111101",28859 => "11001101",28860 => "00000010",28861 => "01110011",28862 => "10010100",28863 => "11011000",28864 => "11101111",28865 => "00010100",28866 => "11010001",28867 => "01010101",28868 => "10001011",28869 => "11111110",28870 => "11101010",28871 => "10001001",28872 => "00011110",28873 => "00110110",28874 => "11110111",28875 => "10111111",28876 => "11011111",28877 => "10100001",28878 => "00001100",28879 => "11110001",28880 => "10001111",28881 => "11101011",28882 => "10100110",28883 => "11010100",28884 => "11001000",28885 => "11101111",28886 => "10101000",28887 => "01101010",28888 => "10101110",28889 => "11011011",28890 => "00101010",28891 => "00000000",28892 => "10110001",28893 => "10101011",28894 => "00110101",28895 => "11010110",28896 => "01101111",28897 => "10011000",28898 => "00000111",28899 => "00011111",28900 => "01001011",28901 => "10111101",28902 => "01101111",28903 => "11011000",28904 => "01011011",28905 => "11101011",28906 => "00001000",28907 => "10101110",28908 => "11110100",28909 => "01111110",28910 => "00011010",28911 => "11110100",28912 => "01110110",28913 => "11000001",28914 => "00000011",28915 => "11100010",28916 => "00001010",28917 => "00001110",28918 => "01001010",28919 => "00011011",28920 => "01001001",28921 => "01100110",28922 => "00110110",28923 => "00000000",28924 => "11111100",28925 => "00100010",28926 => "01001100",28927 => "10101101",28928 => "11011011",28929 => "00010110",28930 => "00010111",28931 => "00011100",28932 => "11001010",28933 => "00100011",28934 => "00001110",28935 => "11001011",28936 => "01000111",28937 => "11101111",28938 => "00001101",28939 => "11001011",28940 => "11111110",28941 => "01000111",28942 => "10010011",28943 => "11100000",28944 => "10100010",28945 => "10001111",28946 => "00111101",28947 => "00000110",28948 => "00011011",28949 => "11000000",28950 => "00100110",28951 => "01111001",28952 => "00111001",28953 => "01000111",28954 => "00111111",28955 => "10110010",28956 => "10101100",28957 => "01001011",28958 => "10000000",28959 => "10011111",28960 => "00010101",28961 => "10110011",28962 => "11110000",28963 => "11111010",28964 => "10011101",28965 => "11101101",28966 => "01100001",28967 => "10111000",28968 => "00101101",28969 => "00000100",28970 => "00011101",28971 => "00110010",28972 => "00111000",28973 => "11110010",28974 => "10101011",28975 => "00101110",28976 => "00011010",28977 => "11011110",28978 => "01011011",28979 => "01100101",28980 => "01011101",28981 => "00100111",28982 => "01100001",28983 => "01001101",28984 => "10110100",28985 => "00001101",28986 => "00100000",28987 => "11111010",28988 => "11011000",28989 => "01100111",28990 => "11000001",28991 => "00001110",28992 => "01011010",28993 => "10011101",28994 => "00000011",28995 => "10111110",28996 => "10010101",28997 => "11110011",28998 => "10010110",28999 => "00101000",29000 => "01111001",29001 => "10100000",29002 => "11110010",29003 => "01111000",29004 => "11010111",29005 => "00000010",29006 => "10100001",29007 => "11000010",29008 => "11101111",29009 => "10001110",29010 => "00111001",29011 => "10000100",29012 => "00101000",29013 => "10000110",29014 => "00001101",29015 => "11100110",29016 => "10011011",29017 => "01000000",29018 => "00110000",29019 => "10111011",29020 => "01111011",29021 => "01001111",29022 => "11100110",29023 => "00000001",29024 => "11010010",29025 => "10010011",29026 => "11110101",29027 => "11101111",29028 => "00011011",29029 => "11101100",29030 => "01010001",29031 => "11011011",29032 => "11101010",29033 => "10010110",29034 => "11111100",29035 => "11100101",29036 => "01100111",29037 => "11110010",29038 => "11100000",29039 => "11101000",29040 => "11100100",29041 => "01001000",29042 => "00111110",29043 => "00100000",29044 => "01000100",29045 => "00010101",29046 => "00011011",29047 => "01111101",29048 => "00100100",29049 => "01111011",29050 => "10010101",29051 => "10111010",29052 => "10000001",29053 => "01010110",29054 => "00110000",29055 => "10011101",29056 => "10100010",29057 => "00010110",29058 => "01111100",29059 => "10010010",29060 => "01011010",29061 => "10001101",29062 => "01000011",29063 => "10011100",29064 => "01100001",29065 => "01001110",29066 => "01011100",29067 => "10101110",29068 => "11101000",29069 => "11100011",29070 => "11001000",29071 => "01110001",29072 => "01100100",29073 => "10101000",29074 => "01100101",29075 => "10110101",29076 => "11110011",29077 => "01010000",29078 => "10000001",29079 => "11011000",29080 => "01110001",29081 => "11000100",29082 => "00010011",29083 => "11100110",29084 => "10011000",29085 => "00011100",29086 => "00100001",29087 => "10111111",29088 => "11010011",29089 => "10000001",29090 => "00011011",29091 => "10100010",29092 => "11001111",29093 => "00011010",29094 => "01011010",29095 => "10101011",29096 => "00100001",29097 => "10010111",29098 => "11110100",29099 => "10100100",29100 => "11011101",29101 => "01001101",29102 => "10100111",29103 => "00100110",29104 => "10001111",29105 => "11111011",29106 => "01111111",29107 => "01110011",29108 => "10000101",29109 => "00111000",29110 => "00001110",29111 => "10001000",29112 => "11000101",29113 => "10011110",29114 => "10001111",29115 => "01111010",29116 => "00111001",29117 => "00011011",29118 => "11001000",29119 => "11000001",29120 => "10011000",29121 => "01111110",29122 => "00000111",29123 => "01101111",29124 => "10010111",29125 => "01001110",29126 => "11110001",29127 => "00110110",29128 => "01001100",29129 => "11111011",29130 => "00001001",29131 => "00111010",29132 => "01010010",29133 => "00110001",29134 => "11000111",29135 => "10110011",29136 => "11000011",29137 => "00001001",29138 => "10111111",29139 => "01000001",29140 => "11100001",29141 => "01011110",29142 => "01010000",29143 => "10001110",29144 => "00001001",29145 => "01011101",29146 => "11110110",29147 => "11100111",29148 => "00110010",29149 => "11101000",29150 => "01000111",29151 => "11110101",29152 => "11101001",29153 => "10100010",29154 => "01111011",29155 => "10001110",29156 => "01101011",29157 => "10110001",29158 => "00111000",29159 => "11100011",29160 => "00111000",29161 => "01110100",29162 => "10100111",29163 => "10010011",29164 => "11111001",29165 => "01101000",29166 => "00000100",29167 => "01100000",29168 => "10000111",29169 => "01110011",29170 => "01011000",29171 => "10000111",29172 => "10011100",29173 => "00000100",29174 => "00010101",29175 => "00101111",29176 => "00010111",29177 => "00001010",29178 => "11101000",29179 => "00011111",29180 => "00100101",29181 => "00111110",29182 => "01101110",29183 => "01000010",29184 => "11011001",29185 => "01111100",29186 => "01101101",29187 => "00101111",29188 => "11111111",29189 => "00011111",29190 => "11010101",29191 => "11011001",29192 => "11001011",29193 => "00100010",29194 => "11100111",29195 => "01000101",29196 => "00011000",29197 => "00110110",29198 => "01110011",29199 => "00110000",29200 => "11110101",29201 => "10111011",29202 => "01011100",29203 => "01100101",29204 => "00110001",29205 => "00100000",29206 => "00000111",29207 => "10011100",29208 => "10001011",29209 => "00010100",29210 => "11001101",29211 => "11110011",29212 => "01010010",29213 => "10101101",29214 => "10110001",29215 => "10110110",29216 => "01110101",29217 => "10100010",29218 => "01100000",29219 => "00101100",29220 => "00011000",29221 => "11001011",29222 => "01101101",29223 => "00000110",29224 => "10110000",29225 => "00000010",29226 => "00111101",29227 => "00001111",29228 => "10010101",29229 => "11010101",29230 => "11100110",29231 => "10100011",29232 => "11100111",29233 => "11101100",29234 => "00101101",29235 => "10010001",29236 => "01110101",29237 => "11000110",29238 => "10011111",29239 => "10101001",29240 => "11011000",29241 => "11100101",29242 => "11010010",29243 => "10001001",29244 => "10001110",29245 => "00111001",29246 => "10000111",29247 => "10110011",29248 => "10011000",29249 => "10011111",29250 => "01111011",29251 => "10000110",29252 => "10010001",29253 => "11011001",29254 => "00111111",29255 => "11011011",29256 => "00101000",29257 => "11000001",29258 => "00010001",29259 => "00011011",29260 => "00010101",29261 => "11010100",29262 => "01011011",29263 => "01010110",29264 => "11010010",29265 => "10111100",29266 => "10000111",29267 => "11100000",29268 => "00110000",29269 => "11010010",29270 => "11100100",29271 => "00011001",29272 => "00111111",29273 => "01000010",29274 => "10000000",29275 => "01011001",29276 => "00010000",29277 => "11001101",29278 => "10101001",29279 => "11011100",29280 => "00101101",29281 => "01011111",29282 => "00010111",29283 => "01100110",29284 => "10110110",29285 => "00001000",29286 => "10011111",29287 => "01010000",29288 => "01010000",29289 => "00001010",29290 => "10111111",29291 => "00111000",29292 => "01101100",29293 => "10111110",29294 => "10011111",29295 => "11111010",29296 => "00100001",29297 => "01110100",29298 => "01010001",29299 => "11101101",29300 => "10001100",29301 => "00010101",29302 => "10100100",29303 => "10110010",29304 => "11011000",29305 => "01100100",29306 => "00111110",29307 => "01111100",29308 => "10110100",29309 => "10001111",29310 => "00001000",29311 => "10010000",29312 => "10100111",29313 => "11101010",29314 => "11110110",29315 => "01000001",29316 => "11010000",29317 => "00000011",29318 => "10010001",29319 => "11001001",29320 => "01111100",29321 => "01001010",29322 => "01111110",29323 => "10101101",29324 => "11111111",29325 => "10101010",29326 => "11011101",29327 => "10100011",29328 => "11111110",29329 => "01100110",29330 => "00110111",29331 => "11101101",29332 => "10110100",29333 => "01101100",29334 => "10011110",29335 => "00110011",29336 => "00100110",29337 => "00010100",29338 => "11101100",29339 => "01100001",29340 => "11000100",29341 => "00001001",29342 => "00001110",29343 => "01010011",29344 => "11000010",29345 => "11101000",29346 => "10111101",29347 => "11100001",29348 => "11110001",29349 => "10000010",29350 => "01100101",29351 => "00001000",29352 => "11000100",29353 => "00011110",29354 => "00010100",29355 => "10101101",29356 => "01111010",29357 => "11000100",29358 => "10110001",29359 => "10010001",29360 => "00100011",29361 => "00010111",29362 => "11110001",29363 => "10110100",29364 => "01001110",29365 => "10100011",29366 => "00011111",29367 => "11011110",29368 => "11101010",29369 => "10011011",29370 => "01101000",29371 => "10110001",29372 => "00001001",29373 => "01100000",29374 => "11101110",29375 => "11110101",29376 => "01111101",29377 => "11101001",29378 => "11101011",29379 => "01111010",29380 => "10101000",29381 => "01010100",29382 => "00100010",29383 => "01000110",29384 => "11100101",29385 => "00010010",29386 => "10011001",29387 => "01000111",29388 => "01101000",29389 => "10011001",29390 => "00101101",29391 => "11001000",29392 => "01000101",29393 => "10111010",29394 => "10111100",29395 => "00001010",29396 => "11000011",29397 => "01110110",29398 => "11101101",29399 => "01100100",29400 => "10110100",29401 => "01101111",29402 => "11011100",29403 => "10111000",29404 => "01101111",29405 => "11111101",29406 => "10101001",29407 => "10011010",29408 => "01110100",29409 => "01111001",29410 => "10100110",29411 => "01001110",29412 => "11011010",29413 => "01101111",29414 => "11000111",29415 => "10001001",29416 => "00100010",29417 => "10110011",29418 => "00010000",29419 => "00111001",29420 => "00000011",29421 => "10010101",29422 => "11100111",29423 => "11100000",29424 => "10011100",29425 => "01011100",29426 => "00010100",29427 => "00010111",29428 => "10001001",29429 => "00111110",29430 => "01001000",29431 => "10110000",29432 => "00110001",29433 => "11100011",29434 => "00000011",29435 => "00110100",29436 => "01011011",29437 => "01111111",29438 => "01100110",29439 => "00001010",29440 => "11101001",29441 => "00111011",29442 => "11011100",29443 => "01100111",29444 => "11011110",29445 => "01100111",29446 => "00110110",29447 => "01001011",29448 => "10001101",29449 => "10000011",29450 => "11100000",29451 => "00001001",29452 => "10010010",29453 => "01001011",29454 => "01010111",29455 => "10001111",29456 => "10111011",29457 => "00101101",29458 => "10011010",29459 => "10001011",29460 => "00011011",29461 => "00011010",29462 => "00011101",29463 => "00110100",29464 => "01101010",29465 => "11110001",29466 => "00110111",29467 => "11101011",29468 => "00001100",29469 => "00111100",29470 => "01101000",29471 => "01000001",29472 => "01011010",29473 => "00101110",29474 => "10111001",29475 => "00011010",29476 => "00010101",29477 => "11011100",29478 => "01011101",29479 => "00110010",29480 => "01101011",29481 => "11110111",29482 => "01001000",29483 => "01100000",29484 => "00111011",29485 => "00011110",29486 => "00101110",29487 => "00001000",29488 => "11101101",29489 => "10011110",29490 => "10100110",29491 => "10110011",29492 => "11110010",29493 => "01000010",29494 => "11101001",29495 => "10110110",29496 => "10110011",29497 => "01101111",29498 => "01110001",29499 => "11011111",29500 => "00110011",29501 => "01011111",29502 => "00011011",29503 => "10101001",29504 => "01000010",29505 => "01110101",29506 => "11101100",29507 => "01010111",29508 => "01110000",29509 => "11110110",29510 => "10111011",29511 => "11011110",29512 => "11000011",29513 => "10110000",29514 => "01011110",29515 => "00110100",29516 => "11011001",29517 => "00000011",29518 => "10001000",29519 => "11101100",29520 => "11001100",29521 => "01001111",29522 => "00000100",29523 => "10101101",29524 => "10100110",29525 => "10110011",29526 => "11111001",29527 => "10001100",29528 => "00000011",29529 => "00101101",29530 => "00111010",29531 => "11100101",29532 => "00110100",29533 => "11100001",29534 => "10110011",29535 => "10111010",29536 => "10010101",29537 => "00111110",29538 => "00110001",29539 => "10101010",29540 => "10001101",29541 => "10110110",29542 => "01000111",29543 => "01110111",29544 => "10110010",29545 => "00000000",29546 => "11010111",29547 => "10010001",29548 => "10001101",29549 => "10010011",29550 => "00111011",29551 => "01001110",29552 => "00011110",29553 => "01011100",29554 => "10000000",29555 => "11100001",29556 => "01010001",29557 => "01111001",29558 => "11110000",29559 => "11010000",29560 => "11000010",29561 => "00110000",29562 => "01110000",29563 => "00100011",29564 => "00001011",29565 => "10101010",29566 => "00010100",29567 => "11000101",29568 => "00100000",29569 => "00111101",29570 => "00111001",29571 => "11001111",29572 => "00100010",29573 => "10101100",29574 => "01010010",29575 => "00100110",29576 => "11000011",29577 => "10001100",29578 => "10111010",29579 => "01111011",29580 => "11101110",29581 => "01001110",29582 => "01011010",29583 => "01010110",29584 => "00001111",29585 => "01110000",29586 => "10101000",29587 => "01000001",29588 => "10010001",29589 => "00001010",29590 => "01101001",29591 => "01101010",29592 => "11001100",29593 => "00001100",29594 => "10101010",29595 => "11100000",29596 => "10110101",29597 => "00111111",29598 => "11011110",29599 => "01100100",29600 => "10101110",29601 => "11000011",29602 => "10010001",29603 => "00011010",29604 => "00101010",29605 => "11100100",29606 => "00111110",29607 => "11101000",29608 => "00100011",29609 => "01011101",29610 => "01000110",29611 => "00000111",29612 => "10010001",29613 => "11111101",29614 => "01000100",29615 => "10110010",29616 => "10001101",29617 => "10110000",29618 => "11101101",29619 => "10011001",29620 => "11100010",29621 => "11011111",29622 => "11001110",29623 => "00111111",29624 => "11100101",29625 => "10010000",29626 => "10000011",29627 => "11110111",29628 => "01110001",29629 => "10111100",29630 => "10010001",29631 => "10111010",29632 => "10010010",29633 => "00001001",29634 => "11010001",29635 => "11001111",29636 => "00000110",29637 => "01101110",29638 => "00000001",29639 => "01111011",29640 => "10111000",29641 => "11000110",29642 => "00010000",29643 => "10010000",29644 => "11010000",29645 => "11100001",29646 => "11011000",29647 => "00010011",29648 => "10001101",29649 => "11001001",29650 => "10111111",29651 => "01000001",29652 => "11010000",29653 => "00001001",29654 => "11111101",29655 => "11110101",29656 => "11000000",29657 => "01001011",29658 => "11111010",29659 => "11111101",29660 => "11100001",29661 => "11010101",29662 => "11001010",29663 => "10100000",29664 => "01011100",29665 => "10010111",29666 => "11011101",29667 => "00000111",29668 => "01010010",29669 => "10111101",29670 => "00001111",29671 => "01010100",29672 => "11011000",29673 => "00010100",29674 => "01100011",29675 => "01100011",29676 => "00001000",29677 => "10011010",29678 => "00111101",29679 => "11101010",29680 => "10111100",29681 => "01110000",29682 => "10001011",29683 => "00011100",29684 => "10001000",29685 => "10100001",29686 => "01100011",29687 => "11111000",29688 => "00110101",29689 => "11110101",29690 => "10110111",29691 => "10110011",29692 => "00011111",29693 => "11010000",29694 => "10110011",29695 => "10011111",29696 => "11101001",29697 => "00110001",29698 => "00111110",29699 => "01110110",29700 => "01111101",29701 => "01100001",29702 => "01001100",29703 => "11000011",29704 => "00010100",29705 => "01011010",29706 => "11010101",29707 => "11110110",29708 => "11110111",29709 => "01110110",29710 => "00111001",29711 => "10010111",29712 => "01010000",29713 => "10110111",29714 => "10110011",29715 => "11011101",29716 => "00011110",29717 => "11111111",29718 => "10010011",29719 => "10111101",29720 => "00011110",29721 => "01111011",29722 => "10010011",29723 => "00001100",29724 => "01100111",29725 => "11011010",29726 => "10000111",29727 => "11010100",29728 => "00101101",29729 => "10111000",29730 => "10010110",29731 => "00110111",29732 => "01010000",29733 => "01111101",29734 => "10010110",29735 => "01000011",29736 => "01111000",29737 => "10101010",29738 => "10011110",29739 => "01101011",29740 => "01111111",29741 => "00110011",29742 => "11110101",29743 => "01100111",29744 => "00101100",29745 => "01111100",29746 => "11000010",29747 => "01001010",29748 => "11010010",29749 => "11011011",29750 => "10110111",29751 => "00010101",29752 => "11100001",29753 => "10111111",29754 => "10011010",29755 => "10101011",29756 => "01010101",29757 => "10000001",29758 => "00101000",29759 => "01011001",29760 => "00111111",29761 => "01011100",29762 => "00010001",29763 => "01000101",29764 => "11110101",29765 => "11100111",29766 => "00001100",29767 => "11011110",29768 => "01011111",29769 => "00110110",29770 => "11110001",29771 => "01010100",29772 => "10001011",29773 => "10100111",29774 => "10101011",29775 => "00011001",29776 => "00001111",29777 => "01011000",29778 => "11000101",29779 => "01010100",29780 => "10100010",29781 => "01100111",29782 => "11111101",29783 => "11000001",29784 => "10001001",29785 => "00001001",29786 => "10100110",29787 => "00000110",29788 => "11011010",29789 => "00101011",29790 => "11100001",29791 => "11011000",29792 => "10111111",29793 => "00000111",29794 => "11011011",29795 => "10001010",29796 => "01101010",29797 => "11010011",29798 => "10011100",29799 => "00110111",29800 => "11000111",29801 => "00100111",29802 => "11010011",29803 => "11011010",29804 => "01010100",29805 => "11100011",29806 => "01001010",29807 => "00101110",29808 => "00111001",29809 => "01011111",29810 => "10110101",29811 => "00011001",29812 => "10000000",29813 => "11000101",29814 => "00111001",29815 => "00101001",29816 => "01000001",29817 => "00100101",29818 => "00011011",29819 => "11011001",29820 => "01010101",29821 => "11010000",29822 => "10111000",29823 => "10011001",29824 => "10100101",29825 => "00101011",29826 => "10000100",29827 => "11000010",29828 => "00111101",29829 => "11010011",29830 => "00001011",29831 => "10000111",29832 => "11110110",29833 => "10110111",29834 => "00111110",29835 => "11110110",29836 => "10001110",29837 => "01101110",29838 => "01101011",29839 => "11010001",29840 => "10011011",29841 => "00010110",29842 => "11100101",29843 => "00100111",29844 => "00110010",29845 => "11000000",29846 => "10000010",29847 => "10101111",29848 => "10011000",29849 => "11001000",29850 => "00000011",29851 => "00010110",29852 => "10111000",29853 => "11000001",29854 => "11000111",29855 => "01000100",29856 => "11011001",29857 => "01001001",29858 => "10100111",29859 => "10010011",29860 => "11100000",29861 => "00011001",29862 => "11111001",29863 => "10000001",29864 => "00110001",29865 => "01101010",29866 => "00000010",29867 => "10100010",29868 => "01100111",29869 => "01101011",29870 => "10111111",29871 => "01010001",29872 => "00110000",29873 => "01110111",29874 => "11110110",29875 => "01010111",29876 => "00011111",29877 => "00111010",29878 => "10111100",29879 => "01000000",29880 => "01111100",29881 => "11101010",29882 => "00101001",29883 => "10100110",29884 => "00010101",29885 => "01101000",29886 => "01000011",29887 => "00010111",29888 => "01011011",29889 => "01101010",29890 => "01100111",29891 => "01100100",29892 => "00011110",29893 => "00011110",29894 => "10011010",29895 => "01111011",29896 => "00100010",29897 => "10110011",29898 => "00101010",29899 => "11011011",29900 => "01000010",29901 => "10100100",29902 => "00101110",29903 => "10100100",29904 => "00110010",29905 => "01110000",29906 => "00110100",29907 => "01101010",29908 => "10001110",29909 => "01100101",29910 => "10010110",29911 => "10010100",29912 => "10110100",29913 => "00001001",29914 => "01010100",29915 => "11100010",29916 => "00010011",29917 => "11011000",29918 => "00110110",29919 => "11000101",29920 => "11010101",29921 => "01100010",29922 => "00001000",29923 => "00000000",29924 => "00010010",29925 => "00110000",29926 => "00101001",29927 => "10101000",29928 => "01110000",29929 => "10010010",29930 => "01010011",29931 => "11111100",29932 => "10011110",29933 => "01000100",29934 => "01100111",29935 => "01010111",29936 => "00110110",29937 => "10110011",29938 => "10001110",29939 => "10111000",29940 => "11010010",29941 => "00111011",29942 => "01001011",29943 => "00000100",29944 => "01111100",29945 => "01010111",29946 => "00100100",29947 => "10101000",29948 => "10100000",29949 => "10010000",29950 => "11000100",29951 => "11110100",29952 => "01011000",29953 => "10000110",29954 => "10101000",29955 => "10000001",29956 => "11100100",29957 => "00001110",29958 => "00111000",29959 => "00001010",29960 => "00100100",29961 => "11110010",29962 => "10100110",29963 => "10001111",29964 => "10101110",29965 => "01110110",29966 => "11111100",29967 => "00010100",29968 => "10110010",29969 => "11101110",29970 => "00000101",29971 => "00100010",29972 => "11101001",29973 => "10000111",29974 => "00101010",29975 => "00000010",29976 => "01100000",29977 => "10101011",29978 => "11000100",29979 => "00110000",29980 => "01100010",29981 => "00100101",29982 => "10110001",29983 => "00100000",29984 => "10100010",29985 => "11110001",29986 => "01000110",29987 => "00010001",29988 => "11100110",29989 => "11110101",29990 => "00000010",29991 => "01010000",29992 => "00010101",29993 => "11001000",29994 => "00101110",29995 => "11010101",29996 => "11001111",29997 => "10111010",29998 => "10000101",29999 => "01111000",30000 => "11100011",30001 => "00010000",30002 => "11110111",30003 => "00111100",30004 => "00000001",30005 => "11111101",30006 => "00010110",30007 => "11001001",30008 => "00000100",30009 => "00111111",30010 => "10100100",30011 => "11010000",30012 => "10110100",30013 => "10101110",30014 => "11100100",30015 => "01011110",30016 => "11110110",30017 => "00011100",30018 => "01000000",30019 => "11111001",30020 => "10101000",30021 => "00001100",30022 => "01111100",30023 => "10101001",30024 => "00001101",30025 => "01110111",30026 => "01100001",30027 => "00001010",30028 => "01000100",30029 => "00100101",30030 => "00011111",30031 => "00101011",30032 => "00011001",30033 => "11011010",30034 => "01111000",30035 => "01010000",30036 => "11111010",30037 => "00100111",30038 => "10110101",30039 => "10010100",30040 => "00001100",30041 => "01011011",30042 => "10000010",30043 => "11111101",30044 => "11011110",30045 => "11111000",30046 => "10010111",30047 => "00000011",30048 => "11010011",30049 => "01000010",30050 => "01000001",30051 => "10100010",30052 => "11000100",30053 => "10110111",30054 => "11110010",30055 => "01111001",30056 => "11010100",30057 => "01011011",30058 => "11100010",30059 => "11101000",30060 => "01110000",30061 => "11010001",30062 => "00001010",30063 => "01001000",30064 => "11010110",30065 => "11011100",30066 => "11101010",30067 => "01000011",30068 => "00101100",30069 => "01001010",30070 => "01011111",30071 => "00101110",30072 => "00011011",30073 => "10000001",30074 => "00001011",30075 => "11100101",30076 => "10101100",30077 => "10110001",30078 => "00001001",30079 => "11101001",30080 => "11000111",30081 => "11011101",30082 => "10101111",30083 => "00110111",30084 => "11110110",30085 => "00110010",30086 => "11110000",30087 => "11111111",30088 => "10010110",30089 => "00110111",30090 => "00000110",30091 => "01111101",30092 => "01111011",30093 => "00010000",30094 => "11001111",30095 => "00000010",30096 => "11111000",30097 => "01010001",30098 => "10101110",30099 => "00101100",30100 => "10100011",30101 => "01101110",30102 => "00000110",30103 => "00110000",30104 => "10100000",30105 => "01011011",30106 => "00000111",30107 => "10000101",30108 => "11101111",30109 => "01010000",30110 => "11000100",30111 => "10111110",30112 => "01101011",30113 => "11010100",30114 => "10101101",30115 => "10110111",30116 => "00010011",30117 => "10100110",30118 => "10100110",30119 => "00011111",30120 => "11000001",30121 => "01000011",30122 => "11100100",30123 => "10010110",30124 => "00010011",30125 => "00110010",30126 => "11110010",30127 => "01000011",30128 => "10000111",30129 => "00000111",30130 => "11101101",30131 => "11100000",30132 => "00010010",30133 => "10110101",30134 => "10101111",30135 => "10001011",30136 => "00011100",30137 => "10011101",30138 => "00010100",30139 => "00101110",30140 => "01010111",30141 => "11000000",30142 => "10110011",30143 => "00110011",30144 => "10110011",30145 => "11100110",30146 => "11110001",30147 => "10010100",30148 => "10001101",30149 => "11100000",30150 => "11110101",30151 => "01111100",30152 => "11001111",30153 => "11001101",30154 => "01010001",30155 => "11110100",30156 => "10001011",30157 => "11111001",30158 => "11011110",30159 => "11111000",30160 => "10111011",30161 => "11010000",30162 => "01001101",30163 => "00111111",30164 => "10000111",30165 => "11101110",30166 => "11110100",30167 => "11000010",30168 => "00111111",30169 => "01001101",30170 => "00101000",30171 => "11110110",30172 => "01000011",30173 => "10110100",30174 => "00101100",30175 => "11001000",30176 => "10000011",30177 => "01100010",30178 => "10010100",30179 => "01101110",30180 => "00001101",30181 => "11110110",30182 => "00101001",30183 => "01000110",30184 => "10111101",30185 => "10101100",30186 => "00011010",30187 => "11110101",30188 => "01000100",30189 => "01000000",30190 => "10000111",30191 => "01011000",30192 => "01011100",30193 => "10010101",30194 => "10100000",30195 => "01101000",30196 => "00000101",30197 => "11100100",30198 => "11100011",30199 => "10010001",30200 => "11110011",30201 => "01010000",30202 => "00111110",30203 => "10110101",30204 => "11111100",30205 => "10010100",30206 => "11101011",30207 => "00010001",30208 => "00111001",30209 => "11011001",30210 => "11011111",30211 => "11010110",30212 => "00011011",30213 => "10111010",30214 => "00100100",30215 => "01010111",30216 => "10010100",30217 => "00011011",30218 => "01111001",30219 => "01001001",30220 => "00111011",30221 => "10001111",30222 => "10001000",30223 => "00011101",30224 => "00001100",30225 => "01101011",30226 => "01011000",30227 => "01101001",30228 => "11011111",30229 => "10001010",30230 => "11101101",30231 => "01101111",30232 => "01101011",30233 => "01101000",30234 => "10011011",30235 => "00011101",30236 => "00011001",30237 => "00110000",30238 => "11100100",30239 => "10010000",30240 => "11001100",30241 => "11000111",30242 => "01111101",30243 => "00000100",30244 => "10000010",30245 => "10000001",30246 => "01101000",30247 => "01110101",30248 => "01001011",30249 => "10001001",30250 => "11101000",30251 => "01110000",30252 => "00110110",30253 => "11000101",30254 => "10010000",30255 => "10001100",30256 => "10101000",30257 => "01011001",30258 => "10001111",30259 => "10001001",30260 => "00000110",30261 => "11011101",30262 => "10100101",30263 => "11011000",30264 => "10011010",30265 => "11011100",30266 => "11100111",30267 => "00100110",30268 => "10010110",30269 => "00101001",30270 => "01010011",30271 => "11100010",30272 => "11110010",30273 => "10010111",30274 => "01010110",30275 => "00000001",30276 => "10000111",30277 => "00010101",30278 => "01011111",30279 => "10001111",30280 => "10011101",30281 => "11101000",30282 => "01100010",30283 => "11100011",30284 => "01111100",30285 => "00101010",30286 => "00110011",30287 => "00101000",30288 => "01010111",30289 => "11011000",30290 => "01001000",30291 => "01110001",30292 => "10010111",30293 => "00111001",30294 => "01000010",30295 => "01000001",30296 => "01001000",30297 => "11010100",30298 => "00111111",30299 => "10101110",30300 => "10111000",30301 => "01111100",30302 => "11010011",30303 => "00011010",30304 => "01110101",30305 => "11011001",30306 => "01000100",30307 => "01111101",30308 => "00110001",30309 => "11011010",30310 => "01101111",30311 => "10101000",30312 => "00111011",30313 => "00100011",30314 => "10010110",30315 => "00111011",30316 => "01111001",30317 => "11010000",30318 => "10000111",30319 => "01111111",30320 => "10001011",30321 => "01011111",30322 => "11010110",30323 => "11010011",30324 => "00000100",30325 => "01011111",30326 => "00000111",30327 => "01100011",30328 => "11000011",30329 => "01111000",30330 => "10110011",30331 => "10010000",30332 => "00000011",30333 => "01101100",30334 => "11001000",30335 => "10101101",30336 => "10000011",30337 => "11111111",30338 => "10101000",30339 => "01010001",30340 => "00000111",30341 => "01011001",30342 => "10001001",30343 => "01100000",30344 => "00000110",30345 => "01100000",30346 => "00100100",30347 => "11001101",30348 => "10111000",30349 => "01100010",30350 => "10010000",30351 => "00101110",30352 => "10100010",30353 => "11001001",30354 => "01000111",30355 => "00100001",30356 => "10101111",30357 => "11001010",30358 => "11111110",30359 => "11100010",30360 => "10111001",30361 => "10011101",30362 => "11111000",30363 => "10111000",30364 => "11010111",30365 => "01001110",30366 => "11001011",30367 => "10001001",30368 => "10010111",30369 => "10000100",30370 => "01100101",30371 => "00011010",30372 => "01011011",30373 => "01111010",30374 => "10111101",30375 => "01111110",30376 => "01001001",30377 => "11011011",30378 => "11111101",30379 => "11100010",30380 => "10100111",30381 => "01100000",30382 => "01110011",30383 => "00010100",30384 => "01000010",30385 => "00111000",30386 => "10101100",30387 => "10100001",30388 => "10011110",30389 => "11110010",30390 => "11100001",30391 => "01100011",30392 => "10001010",30393 => "00001100",30394 => "01001010",30395 => "00011111",30396 => "00011111",30397 => "10000110",30398 => "01100101",30399 => "01101111",30400 => "01001010",30401 => "10011101",30402 => "01011010",30403 => "00100011",30404 => "11111001",30405 => "00101111",30406 => "10000000",30407 => "11111010",30408 => "00001111",30409 => "01101000",30410 => "00010010",30411 => "10001111",30412 => "10010011",30413 => "00111100",30414 => "11000001",30415 => "10101011",30416 => "01100000",30417 => "10111001",30418 => "11110001",30419 => "00100101",30420 => "11011011",30421 => "00101100",30422 => "01010101",30423 => "01011000",30424 => "11101110",30425 => "01101011",30426 => "00011001",30427 => "10010000",30428 => "00100011",30429 => "11000011",30430 => "10100100",30431 => "10100010",30432 => "11111000",30433 => "10100110",30434 => "01001000",30435 => "11010010",30436 => "10110100",30437 => "01111101",30438 => "10011111",30439 => "00111100",30440 => "00101100",30441 => "11011001",30442 => "01011000",30443 => "01101111",30444 => "00100000",30445 => "11011110",30446 => "00111001",30447 => "00110001",30448 => "11011010",30449 => "10110100",30450 => "10001011",30451 => "10100001",30452 => "10001000",30453 => "00001110",30454 => "00010011",30455 => "01110111",30456 => "00111000",30457 => "00110011",30458 => "01110010",30459 => "01101011",30460 => "00000100",30461 => "11010010",30462 => "01100001",30463 => "01000101",30464 => "01011101",30465 => "00011111",30466 => "10111001",30467 => "11000110",30468 => "00011100",30469 => "10000010",30470 => "00010010",30471 => "00011111",30472 => "11100001",30473 => "01001001",30474 => "11011001",30475 => "01011111",30476 => "00100000",30477 => "01010110",30478 => "01111101",30479 => "10110111",30480 => "01010111",30481 => "00111101",30482 => "00010000",30483 => "10111101",30484 => "01000111",30485 => "01110100",30486 => "11001111",30487 => "11011011",30488 => "01011000",30489 => "00111000",30490 => "00000111",30491 => "11011111",30492 => "10010101",30493 => "00000011",30494 => "11010011",30495 => "00001011",30496 => "01101010",30497 => "00101010",30498 => "10010001",30499 => "11111000",30500 => "01001011",30501 => "10001011",30502 => "00111110",30503 => "11100111",30504 => "00001110",30505 => "10001101",30506 => "10000110",30507 => "01001010",30508 => "00101111",30509 => "00101110",30510 => "10100101",30511 => "11001101",30512 => "11000110",30513 => "00100110",30514 => "11111001",30515 => "00100101",30516 => "00011110",30517 => "11110100",30518 => "11101010",30519 => "10011000",30520 => "11111010",30521 => "10011100",30522 => "01010000",30523 => "00010101",30524 => "00110000",30525 => "10100100",30526 => "00000010",30527 => "00110000",30528 => "10111110",30529 => "10000110",30530 => "01110110",30531 => "00101000",30532 => "01011001",30533 => "10011100",30534 => "11111011",30535 => "01000011",30536 => "01101110",30537 => "10101111",30538 => "00111001",30539 => "01000110",30540 => "10110001",30541 => "01011011",30542 => "10101011",30543 => "10010110",30544 => "01100101",30545 => "11100111",30546 => "10001101",30547 => "10110110",30548 => "11111010",30549 => "01000000",30550 => "01111001",30551 => "10110111",30552 => "01010010",30553 => "10010001",30554 => "00010111",30555 => "00110010",30556 => "01011100",30557 => "11110100",30558 => "11110011",30559 => "11111100",30560 => "10111101",30561 => "01110001",30562 => "10100011",30563 => "01010100",30564 => "00101101",30565 => "11000100",30566 => "01011001",30567 => "00000000",30568 => "01001011",30569 => "11110111",30570 => "11111100",30571 => "11110001",30572 => "01011101",30573 => "01100110",30574 => "10101101",30575 => "01000010",30576 => "01111011",30577 => "11011001",30578 => "10110001",30579 => "00011001",30580 => "00000110",30581 => "00000001",30582 => "11111011",30583 => "01111011",30584 => "10101101",30585 => "01010001",30586 => "01100101",30587 => "11111001",30588 => "11100101",30589 => "11010011",30590 => "10111101",30591 => "10011100",30592 => "10010000",30593 => "00110011",30594 => "11101111",30595 => "10110000",30596 => "00001100",30597 => "11010000",30598 => "11111100",30599 => "01101011",30600 => "11011110",30601 => "10010101",30602 => "01011010",30603 => "00000001",30604 => "10100100",30605 => "01101001",30606 => "00101111",30607 => "10011110",30608 => "01110101",30609 => "01101000",30610 => "01110000",30611 => "11110000",30612 => "11101110",30613 => "00000000",30614 => "11010100",30615 => "11010001",30616 => "00010010",30617 => "11111111",30618 => "01001001",30619 => "01100000",30620 => "10011011",30621 => "01000000",30622 => "01010100",30623 => "00010011",30624 => "00100010",30625 => "10111111",30626 => "10101011",30627 => "11100100",30628 => "00000011",30629 => "11001010",30630 => "00011000",30631 => "00110110",30632 => "10110010",30633 => "10110011",30634 => "11100110",30635 => "00110100",30636 => "11001101",30637 => "00100101",30638 => "10110110",30639 => "11001100",30640 => "00111001",30641 => "01111101",30642 => "01111011",30643 => "00110010",30644 => "01010001",30645 => "01101110",30646 => "01011111",30647 => "00001001",30648 => "00100010",30649 => "00101111",30650 => "11101011",30651 => "11001101",30652 => "00110000",30653 => "10000000",30654 => "10011011",30655 => "11011110",30656 => "00101010",30657 => "10111010",30658 => "01001110",30659 => "10111000",30660 => "10001100",30661 => "00001100",30662 => "01100000",30663 => "00001010",30664 => "10110111",30665 => "11011001",30666 => "00100100",30667 => "01010101",30668 => "11100000",30669 => "10010111",30670 => "01111000",30671 => "11011001",30672 => "01011000",30673 => "11010111",30674 => "10100001",30675 => "10100000",30676 => "10010101",30677 => "01001111",30678 => "10101010",30679 => "00101101",30680 => "11111111",30681 => "10101000",30682 => "00100011",30683 => "01010001",30684 => "00010100",30685 => "01000000",30686 => "00101111",30687 => "00110101",30688 => "10011001",30689 => "10011111",30690 => "10100000",30691 => "01100011",30692 => "10000011",30693 => "11111111",30694 => "11001010",30695 => "00101010",30696 => "10101010",30697 => "00001111",30698 => "10111101",30699 => "10111100",30700 => "00111111",30701 => "10110011",30702 => "11101001",30703 => "00011101",30704 => "00000000",30705 => "01110001",30706 => "11101111",30707 => "00111111",30708 => "00000111",30709 => "11110001",30710 => "11100010",30711 => "10011101",30712 => "00101100",30713 => "00000101",30714 => "11011111",30715 => "00100000",30716 => "01111101",30717 => "11001111",30718 => "00100101",30719 => "10011111",30720 => "11100011",30721 => "10101110",30722 => "01011001",30723 => "00111110",30724 => "11100001",30725 => "00101001",30726 => "10110100",30727 => "11111010",30728 => "01111100",30729 => "01010001",30730 => "00011010",30731 => "11100110",30732 => "10111101",30733 => "01110101",30734 => "10111110",30735 => "01011110",30736 => "10100011",30737 => "10110100",30738 => "11100111",30739 => "00111011",30740 => "10110011",30741 => "00000001",30742 => "00010010",30743 => "00000000",30744 => "10011111",30745 => "01111000",30746 => "11100001",30747 => "10000000",30748 => "01100101",30749 => "01001011",30750 => "10111010",30751 => "11110010",30752 => "01111000",30753 => "10000101",30754 => "00111101",30755 => "11111001",30756 => "10001101",30757 => "11000000",30758 => "11001011",30759 => "10101101",30760 => "01111010",30761 => "01010110",30762 => "10111101",30763 => "11000111",30764 => "01110111",30765 => "01100000",30766 => "01011111",30767 => "11100100",30768 => "11111011",30769 => "10010011",30770 => "01111110",30771 => "10101011",30772 => "11010011",30773 => "11010101",30774 => "00000001",30775 => "11110011",30776 => "10001110",30777 => "01111101",30778 => "10100111",30779 => "11101110",30780 => "10010010",30781 => "00111110",30782 => "00011000",30783 => "01000111",30784 => "10111000",30785 => "11101110",30786 => "11001010",30787 => "11010100",30788 => "11110111",30789 => "00100110",30790 => "11110001",30791 => "11111000",30792 => "10110010",30793 => "00011110",30794 => "10011111",30795 => "00000010",30796 => "01000001",30797 => "00111101",30798 => "10100100",30799 => "01000101",30800 => "00001010",30801 => "00110100",30802 => "11001010",30803 => "00111110",30804 => "10100111",30805 => "11111000",30806 => "00001101",30807 => "11100110",30808 => "01010011",30809 => "10010101",30810 => "11100010",30811 => "01111001",30812 => "11001100",30813 => "01100010",30814 => "00011000",30815 => "01101100",30816 => "00110001",30817 => "11101100",30818 => "11000010",30819 => "11110000",30820 => "11111010",30821 => "11001111",30822 => "01110000",30823 => "10101001",30824 => "01000010",30825 => "01010001",30826 => "10111100",30827 => "01100000",30828 => "10000010",30829 => "11001100",30830 => "00101111",30831 => "01111000",30832 => "01011111",30833 => "00011110",30834 => "10101101",30835 => "10010101",30836 => "11001101",30837 => "01110111",30838 => "00001101",30839 => "00010001",30840 => "10001110",30841 => "11101111",30842 => "00001110",30843 => "11011100",30844 => "00100011",30845 => "11101011",30846 => "00011001",30847 => "10111100",30848 => "00011000",30849 => "10100010",30850 => "11000101",30851 => "00011100",30852 => "10100010",30853 => "00111001",30854 => "00110011",30855 => "01011000",30856 => "11100000",30857 => "10000110",30858 => "11111101",30859 => "00100001",30860 => "00011001",30861 => "11111011",30862 => "11110011",30863 => "10101111",30864 => "10111000",30865 => "00101100",30866 => "11011001",30867 => "01001011",30868 => "11100011",30869 => "10100101",30870 => "10000010",30871 => "11001000",30872 => "10111010",30873 => "00100111",30874 => "10110000",30875 => "00011110",30876 => "01100001",30877 => "11101000",30878 => "10001011",30879 => "01001001",30880 => "11010000",30881 => "11010010",30882 => "01110100",30883 => "11001101",30884 => "01110010",30885 => "01001010",30886 => "10011111",30887 => "11110100",30888 => "01001000",30889 => "11111001",30890 => "00000010",30891 => "11110000",30892 => "10110011",30893 => "10001011",30894 => "00111001",30895 => "11010010",30896 => "11010011",30897 => "10010011",30898 => "11111000",30899 => "11100100",30900 => "00011001",30901 => "10010100",30902 => "00101000",30903 => "11111000",30904 => "10110001",30905 => "01001101",30906 => "11100010",30907 => "10100010",30908 => "00001101",30909 => "00001001",30910 => "00010010",30911 => "01001110",30912 => "11000010",30913 => "00111111",30914 => "11011100",30915 => "11110001",30916 => "10100011",30917 => "10011000",30918 => "01101010",30919 => "01111110",30920 => "00010100",30921 => "01101101",30922 => "11111000",30923 => "01100100",30924 => "01111111",30925 => "01101001",30926 => "11010101",30927 => "10110100",30928 => "11000001",30929 => "01010000",30930 => "10000111",30931 => "00111100",30932 => "00010011",30933 => "00100010",30934 => "00111110",30935 => "11010110",30936 => "01100011",30937 => "01110111",30938 => "10011111",30939 => "11110001",30940 => "00000101",30941 => "11110000",30942 => "11101100",30943 => "00110100",30944 => "10111010",30945 => "11111010",30946 => "10011101",30947 => "01011111",30948 => "00001101",30949 => "11000110",30950 => "01100101",30951 => "01100000",30952 => "11101111",30953 => "10110010",30954 => "11111001",30955 => "10001011",30956 => "01000111",30957 => "11110001",30958 => "11101101",30959 => "10110000",30960 => "01010100",30961 => "00111101",30962 => "00100100",30963 => "11000100",30964 => "11110011",30965 => "00000111",30966 => "10000011",30967 => "10011011",30968 => "11101111",30969 => "01001001",30970 => "00100111",30971 => "10011010",30972 => "10110001",30973 => "11111110",30974 => "10111000",30975 => "10011101",30976 => "10101110",30977 => "10110011",30978 => "01100011",30979 => "00111110",30980 => "00010001",30981 => "01010111",30982 => "11000111",30983 => "00111100",30984 => "10001001",30985 => "10010100",30986 => "01111000",30987 => "01000000",30988 => "11011110",30989 => "00110111",30990 => "01111100",30991 => "10001100",30992 => "11011010",30993 => "11010111",30994 => "11111010",30995 => "01110110",30996 => "00001101",30997 => "10101001",30998 => "00100011",30999 => "11000101",31000 => "10101000",31001 => "01110000",31002 => "01101001",31003 => "11011011",31004 => "00111011",31005 => "00110011",31006 => "11001100",31007 => "11111101",31008 => "01111111",31009 => "10000100",31010 => "00000000",31011 => "11001001",31012 => "00110000",31013 => "10010101",31014 => "11110100",31015 => "01000001",31016 => "10001101",31017 => "00110110",31018 => "10010010",31019 => "10010110",31020 => "00101010",31021 => "00001101",31022 => "11010101",31023 => "10100011",31024 => "01000011",31025 => "10000000",31026 => "10001001",31027 => "10111101",31028 => "01011011",31029 => "11110100",31030 => "00101100",31031 => "10001011",31032 => "00100001",31033 => "01111010",31034 => "11011000",31035 => "10101100",31036 => "10101011",31037 => "11111101",31038 => "00011101",31039 => "01011001",31040 => "11111010",31041 => "11111100",31042 => "00001000",31043 => "11100001",31044 => "01011001",31045 => "00101100",31046 => "01101100",31047 => "11110110",31048 => "10101110",31049 => "00011010",31050 => "11111100",31051 => "10110000",31052 => "10101101",31053 => "10100100",31054 => "10010011",31055 => "01110011",31056 => "10110100",31057 => "00011100",31058 => "00101100",31059 => "11001101",31060 => "11110001",31061 => "11111110",31062 => "01001000",31063 => "10001000",31064 => "10001100",31065 => "10001010",31066 => "10111101",31067 => "11110101",31068 => "01101100",31069 => "00011001",31070 => "10110111",31071 => "01011000",31072 => "11111010",31073 => "00001011",31074 => "00101001",31075 => "10000101",31076 => "01100100",31077 => "11110001",31078 => "00111100",31079 => "10011010",31080 => "00010100",31081 => "10000011",31082 => "10100111",31083 => "10000100",31084 => "00110101",31085 => "01001110",31086 => "10111000",31087 => "10101111",31088 => "00000000",31089 => "11110111",31090 => "10000001",31091 => "00000001",31092 => "11101000",31093 => "11110110",31094 => "11010010",31095 => "10000011",31096 => "10000000",31097 => "00001111",31098 => "01100111",31099 => "00101100",31100 => "01110010",31101 => "10001000",31102 => "11111000",31103 => "01010011",31104 => "01111000",31105 => "11011100",31106 => "11011010",31107 => "10101110",31108 => "01110101",31109 => "00010101",31110 => "00000100",31111 => "11100100",31112 => "11101100",31113 => "00110110",31114 => "11100011",31115 => "11111001",31116 => "10010110",31117 => "01110000",31118 => "11111010",31119 => "00000001",31120 => "01011110",31121 => "11000000",31122 => "00001111",31123 => "11011110",31124 => "00001110",31125 => "11110110",31126 => "10010001",31127 => "10100001",31128 => "11110001",31129 => "00100001",31130 => "11000011",31131 => "10001111",31132 => "00010011",31133 => "00111100",31134 => "00100110",31135 => "01011111",31136 => "00110000",31137 => "11100011",31138 => "10111100",31139 => "00011100",31140 => "01101100",31141 => "11010010",31142 => "01111011",31143 => "01110010",31144 => "11111101",31145 => "00101000",31146 => "10111111",31147 => "10000100",31148 => "00011110",31149 => "11100100",31150 => "01111000",31151 => "01010011",31152 => "10010100",31153 => "11111100",31154 => "11101011",31155 => "01101101",31156 => "10011111",31157 => "01010101",31158 => "01100011",31159 => "00000001",31160 => "01110100",31161 => "00011101",31162 => "11011101",31163 => "10111111",31164 => "10110111",31165 => "01111011",31166 => "00010001",31167 => "00001110",31168 => "00110000",31169 => "10100000",31170 => "00100110",31171 => "10011100",31172 => "11111110",31173 => "10100011",31174 => "10000111",31175 => "00010010",31176 => "00100010",31177 => "10110010",31178 => "11100101",31179 => "10101000",31180 => "00110101",31181 => "11111000",31182 => "10000000",31183 => "10010111",31184 => "10101000",31185 => "01010000",31186 => "00001110",31187 => "00110100",31188 => "01001101",31189 => "10001100",31190 => "00000001",31191 => "11010111",31192 => "00011000",31193 => "10001011",31194 => "11000010",31195 => "11101111",31196 => "00101110",31197 => "00111000",31198 => "11000010",31199 => "00001100",31200 => "01110101",31201 => "11111000",31202 => "01111011",31203 => "11111001",31204 => "10111111",31205 => "11110111",31206 => "01100110",31207 => "10101000",31208 => "10110000",31209 => "10001101",31210 => "00110101",31211 => "11011101",31212 => "01100100",31213 => "11111010",31214 => "00110111",31215 => "10100011",31216 => "01011100",31217 => "00101011",31218 => "01101010",31219 => "00011111",31220 => "11101000",31221 => "00000001",31222 => "00101010",31223 => "01111111",31224 => "10000011",31225 => "10001100",31226 => "00011111",31227 => "01110010",31228 => "00100111",31229 => "10010111",31230 => "00011000",31231 => "01011000",31232 => "00010011",31233 => "01101100",31234 => "00000010",31235 => "11001110",31236 => "00000101",31237 => "11001101",31238 => "01101010",31239 => "00100011",31240 => "01110111",31241 => "10110111",31242 => "10110101",31243 => "00101101",31244 => "00111111",31245 => "00111000",31246 => "11100100",31247 => "10000011",31248 => "01001010",31249 => "00011000",31250 => "01010000",31251 => "10100111",31252 => "00001001",31253 => "00010110",31254 => "00001001",31255 => "11001001",31256 => "00100100",31257 => "01101110",31258 => "11100001",31259 => "01111111",31260 => "01011011",31261 => "01110001",31262 => "10010110",31263 => "11001010",31264 => "00001011",31265 => "01111000",31266 => "10010000",31267 => "10010011",31268 => "01110111",31269 => "00100101",31270 => "01111110",31271 => "01111010",31272 => "01101111",31273 => "01001110",31274 => "10110101",31275 => "00011011",31276 => "01010100",31277 => "01010101",31278 => "10001101",31279 => "11101001",31280 => "01111001",31281 => "10111100",31282 => "00010110",31283 => "11100011",31284 => "01101111",31285 => "11110111",31286 => "11011001",31287 => "01010111",31288 => "10000110",31289 => "11101101",31290 => "01100011",31291 => "11000101",31292 => "10001100",31293 => "11011011",31294 => "01001110",31295 => "00101000",31296 => "00101101",31297 => "00011010",31298 => "00010010",31299 => "00011100",31300 => "10100100",31301 => "10101000",31302 => "00010101",31303 => "01100111",31304 => "11110100",31305 => "00100001",31306 => "01111010",31307 => "11110001",31308 => "01100000",31309 => "01001110",31310 => "01000001",31311 => "10101101",31312 => "01000110",31313 => "00000101",31314 => "10111010",31315 => "00001000",31316 => "00101101",31317 => "10101110",31318 => "11111011",31319 => "11100110",31320 => "00110000",31321 => "10101101",31322 => "10111010",31323 => "10111101",31324 => "00101110",31325 => "11010101",31326 => "10010001",31327 => "11111010",31328 => "10011100",31329 => "01100100",31330 => "01110100",31331 => "00011010",31332 => "10100001",31333 => "00100011",31334 => "00100101",31335 => "01001010",31336 => "10001111",31337 => "11001101",31338 => "00111011",31339 => "00001110",31340 => "00010010",31341 => "00111100",31342 => "01000001",31343 => "00001100",31344 => "00001011",31345 => "01001100",31346 => "01101000",31347 => "10011000",31348 => "11111111",31349 => "11001101",31350 => "11001101",31351 => "11011110",31352 => "01001100",31353 => "00101001",31354 => "10110011",31355 => "11101100",31356 => "00001101",31357 => "11001111",31358 => "00010111",31359 => "11110111",31360 => "11101011",31361 => "00010000",31362 => "10011001",31363 => "10001010",31364 => "11000000",31365 => "10001101",31366 => "00101110",31367 => "00100111",31368 => "00000100",31369 => "11110001",31370 => "01101101",31371 => "01001000",31372 => "10111100",31373 => "10010010",31374 => "01011000",31375 => "01010101",31376 => "01110010",31377 => "00000110",31378 => "01111101",31379 => "10001111",31380 => "01011110",31381 => "11101100",31382 => "00101011",31383 => "01010000",31384 => "11010001",31385 => "10001000",31386 => "10111111",31387 => "10011111",31388 => "00110111",31389 => "10010100",31390 => "01100010",31391 => "00110010",31392 => "11001011",31393 => "01000111",31394 => "11101001",31395 => "01010001",31396 => "01000000",31397 => "11001001",31398 => "00111010",31399 => "11111100",31400 => "00101100",31401 => "00101110",31402 => "11100011",31403 => "00001111",31404 => "01000110",31405 => "11100100",31406 => "10100001",31407 => "11101001",31408 => "00111110",31409 => "00010111",31410 => "10011011",31411 => "00111001",31412 => "11110111",31413 => "10110001",31414 => "00110110",31415 => "10100011",31416 => "11111101",31417 => "00011101",31418 => "11111101",31419 => "01110011",31420 => "11100110",31421 => "00000001",31422 => "00101101",31423 => "11110000",31424 => "00110111",31425 => "00100111",31426 => "00111100",31427 => "00010011",31428 => "00100101",31429 => "11010011",31430 => "10110100",31431 => "10000011",31432 => "01000101",31433 => "10011100",31434 => "10011100",31435 => "10001001",31436 => "10111010",31437 => "10001111",31438 => "10000101",31439 => "11010100",31440 => "00000000",31441 => "01111000",31442 => "00101100",31443 => "01111011",31444 => "10000100",31445 => "10000101",31446 => "11110001",31447 => "10101011",31448 => "01011101",31449 => "01001010",31450 => "11100000",31451 => "10111111",31452 => "11110000",31453 => "11111111",31454 => "00110110",31455 => "01111110",31456 => "00000011",31457 => "01001001",31458 => "01111111",31459 => "10101110",31460 => "11000010",31461 => "01011101",31462 => "10000010",31463 => "11011100",31464 => "00111000",31465 => "00010010",31466 => "00001000",31467 => "00001011",31468 => "00101010",31469 => "00101010",31470 => "01000011",31471 => "01100011",31472 => "11000001",31473 => "11001000",31474 => "01001111",31475 => "11100100",31476 => "00001100",31477 => "10001011",31478 => "11011011",31479 => "10100000",31480 => "10000011",31481 => "10000110",31482 => "00101001",31483 => "00011100",31484 => "01011100",31485 => "10111101",31486 => "01111011",31487 => "10001000",31488 => "10010111",31489 => "00000011",31490 => "00001100",31491 => "01110000",31492 => "10100011",31493 => "01000101",31494 => "01110101",31495 => "11101010",31496 => "01101010",31497 => "10010001",31498 => "10100110",31499 => "00101100",31500 => "01011111",31501 => "01110101",31502 => "10110000",31503 => "10110001",31504 => "01111010",31505 => "01010111",31506 => "00010110",31507 => "10010111",31508 => "00110110",31509 => "10111001",31510 => "10111101",31511 => "11110100",31512 => "10101000",31513 => "11111101",31514 => "01111011",31515 => "01101100",31516 => "00100011",31517 => "11010101",31518 => "11000010",31519 => "00000110",31520 => "10000011",31521 => "10001010",31522 => "01011110",31523 => "00011100",31524 => "11011110",31525 => "10010011",31526 => "01110010",31527 => "10001000",31528 => "00101101",31529 => "00001110",31530 => "11101011",31531 => "11101011",31532 => "11110101",31533 => "10010001",31534 => "10111110",31535 => "11111000",31536 => "00000111",31537 => "10100001",31538 => "00101101",31539 => "00110011",31540 => "11100101",31541 => "10010011",31542 => "00010000",31543 => "00110100",31544 => "01110011",31545 => "10101010",31546 => "11100111",31547 => "11101001",31548 => "11010110",31549 => "00010001",31550 => "10010111",31551 => "01011011",31552 => "01000100",31553 => "10011110",31554 => "11011100",31555 => "11010100",31556 => "01101101",31557 => "11000000",31558 => "10010100",31559 => "00011110",31560 => "00100011",31561 => "00001111",31562 => "10111000",31563 => "11011011",31564 => "11110011",31565 => "10111110",31566 => "01110110",31567 => "01110110",31568 => "00001101",31569 => "00111011",31570 => "10110000",31571 => "11011101",31572 => "01000000",31573 => "01110001",31574 => "11100011",31575 => "00000011",31576 => "10111110",31577 => "00010000",31578 => "01000110",31579 => "11111110",31580 => "00000111",31581 => "11100111",31582 => "10111011",31583 => "01000001",31584 => "00110100",31585 => "11011111",31586 => "00001101",31587 => "10001000",31588 => "10110000",31589 => "10101110",31590 => "11110110",31591 => "10001000",31592 => "11000011",31593 => "00100100",31594 => "10110011",31595 => "01100001",31596 => "00111010",31597 => "01110100",31598 => "10000011",31599 => "11101111",31600 => "01011110",31601 => "10100001",31602 => "00000010",31603 => "01010111",31604 => "11100000",31605 => "00101000",31606 => "10110110",31607 => "10000100",31608 => "00011000",31609 => "11110100",31610 => "11100001",31611 => "01111011",31612 => "00000011",31613 => "11001011",31614 => "00101111",31615 => "00111011",31616 => "01010011",31617 => "10111101",31618 => "00101111",31619 => "01101001",31620 => "10000011",31621 => "01111100",31622 => "11110001",31623 => "00100001",31624 => "01110110",31625 => "10111011",31626 => "00111100",31627 => "11111110",31628 => "00001100",31629 => "00001100",31630 => "11100000",31631 => "10100101",31632 => "00011100",31633 => "11010110",31634 => "01110111",31635 => "01111110",31636 => "00101110",31637 => "11000101",31638 => "11110010",31639 => "00001011",31640 => "11110011",31641 => "11101100",31642 => "00011000",31643 => "11111010",31644 => "01010010",31645 => "11110011",31646 => "10100110",31647 => "00100101",31648 => "00111010",31649 => "01010110",31650 => "00110010",31651 => "10000000",31652 => "01011100",31653 => "10101110",31654 => "01010101",31655 => "10101000",31656 => "01000100",31657 => "00100011",31658 => "00000010",31659 => "10011011",31660 => "10110010",31661 => "11100100",31662 => "01000000",31663 => "10111100",31664 => "00011101",31665 => "11000010",31666 => "00010011",31667 => "10101000",31668 => "01100100",31669 => "11000011",31670 => "11001001",31671 => "00011100",31672 => "11001110",31673 => "10010101",31674 => "01011110",31675 => "00111100",31676 => "00000011",31677 => "00110001",31678 => "00100100",31679 => "10000100",31680 => "01010000",31681 => "00010101",31682 => "11000010",31683 => "11010100",31684 => "10101011",31685 => "01001101",31686 => "00100100",31687 => "11010100",31688 => "10001011",31689 => "10010110",31690 => "01011010",31691 => "00001110",31692 => "01110010",31693 => "10011000",31694 => "11010110",31695 => "00101001",31696 => "11010010",31697 => "11010101",31698 => "00011111",31699 => "10000011",31700 => "00001111",31701 => "01111110",31702 => "01100100",31703 => "01110011",31704 => "01110100",31705 => "01001010",31706 => "01010001",31707 => "00000001",31708 => "01010110",31709 => "10010010",31710 => "11001100",31711 => "10000010",31712 => "00101010",31713 => "00110001",31714 => "01000001",31715 => "10000110",31716 => "11100111",31717 => "10111110",31718 => "00110111",31719 => "00111101",31720 => "11111101",31721 => "00100010",31722 => "00001000",31723 => "01000011",31724 => "01010010",31725 => "01100100",31726 => "11001101",31727 => "01101000",31728 => "00000100",31729 => "10100101",31730 => "10011010",31731 => "11101100",31732 => "00000100",31733 => "10011000",31734 => "01001111",31735 => "10010000",31736 => "10101100",31737 => "01000000",31738 => "00000111",31739 => "11010100",31740 => "00101010",31741 => "00010100",31742 => "01001101",31743 => "00101101",31744 => "00011111",31745 => "00110111",31746 => "00001101",31747 => "00110110",31748 => "10001110",31749 => "10101111",31750 => "11011011",31751 => "00011101",31752 => "10010000",31753 => "10000011",31754 => "01001110",31755 => "11101011",31756 => "00100111",31757 => "11011100",31758 => "00100100",31759 => "11100011",31760 => "00011100",31761 => "11011110",31762 => "11110100",31763 => "10000011",31764 => "11000001",31765 => "01010100",31766 => "11110111",31767 => "01101110",31768 => "00100101",31769 => "11100010",31770 => "01000001",31771 => "11111001",31772 => "11011111",31773 => "11010110",31774 => "11100000",31775 => "00111101",31776 => "00100101",31777 => "11110010",31778 => "01110100",31779 => "11010101",31780 => "00110000",31781 => "10100000",31782 => "11011100",31783 => "11000110",31784 => "00111100",31785 => "10110111",31786 => "01001000",31787 => "11010001",31788 => "10111011",31789 => "10011010",31790 => "10101010",31791 => "00001111",31792 => "01000001",31793 => "11111111",31794 => "00010101",31795 => "01101001",31796 => "11010100",31797 => "11000111",31798 => "01111111",31799 => "00010001",31800 => "10100000",31801 => "00101111",31802 => "01000010",31803 => "11100100",31804 => "01110111",31805 => "01111110",31806 => "01011000",31807 => "10011010",31808 => "11011101",31809 => "10100001",31810 => "01001111",31811 => "01000000",31812 => "10011010",31813 => "11111111",31814 => "01010010",31815 => "10000011",31816 => "00101100",31817 => "01000110",31818 => "10111000",31819 => "01111110",31820 => "11100101",31821 => "01010000",31822 => "00010000",31823 => "11101100",31824 => "01110101",31825 => "10101000",31826 => "01111011",31827 => "00110011",31828 => "10000000",31829 => "00100011",31830 => "01110101",31831 => "10000000",31832 => "01010011",31833 => "10010100",31834 => "00001100",31835 => "10000001",31836 => "10010000",31837 => "01000100",31838 => "10000100",31839 => "10101100",31840 => "10101101",31841 => "11111011",31842 => "01000001",31843 => "11001000",31844 => "10110111",31845 => "00001000",31846 => "01001011",31847 => "01011100",31848 => "10111110",31849 => "00010111",31850 => "10000000",31851 => "00110001",31852 => "01100001",31853 => "11101000",31854 => "00101110",31855 => "00000001",31856 => "01110001",31857 => "11011001",31858 => "00000101",31859 => "01111100",31860 => "00111001",31861 => "11101000",31862 => "00001110",31863 => "10110100",31864 => "01100110",31865 => "01111111",31866 => "10101001",31867 => "01101111",31868 => "11001111",31869 => "00110011",31870 => "10001011",31871 => "01010110",31872 => "11101111",31873 => "11010001",31874 => "11111101",31875 => "10011101",31876 => "00100001",31877 => "00100101",31878 => "00100010",31879 => "10001000",31880 => "01010000",31881 => "10101100",31882 => "10000101",31883 => "01101111",31884 => "00001010",31885 => "10101000",31886 => "01111110",31887 => "01110011",31888 => "01100010",31889 => "01111000",31890 => "10001001",31891 => "11001101",31892 => "00000000",31893 => "10100011",31894 => "11100110",31895 => "11000000",31896 => "01100000",31897 => "01001000",31898 => "10011101",31899 => "11111100",31900 => "01111000",31901 => "10011011",31902 => "10001000",31903 => "00001000",31904 => "10100110",31905 => "00010111",31906 => "10100100",31907 => "01110110",31908 => "11111001",31909 => "01100111",31910 => "00011111",31911 => "01110111",31912 => "01000010",31913 => "01110101",31914 => "11001101",31915 => "01111001",31916 => "11100111",31917 => "01000001",31918 => "00011111",31919 => "11110110",31920 => "11001100",31921 => "11111010",31922 => "10110111",31923 => "10111011",31924 => "11010101",31925 => "11010010",31926 => "11111001",31927 => "00110011",31928 => "11111000",31929 => "10100011",31930 => "11011110",31931 => "00101111",31932 => "00101110",31933 => "01011011",31934 => "00001101",31935 => "11110100",31936 => "01010101",31937 => "01011110",31938 => "10110011",31939 => "00101101",31940 => "00100101",31941 => "01010100",31942 => "10100001",31943 => "00111101",31944 => "10000101",31945 => "11010000",31946 => "11011111",31947 => "10110010",31948 => "11001011",31949 => "11111101",31950 => "00011111",31951 => "00001010",31952 => "11011010",31953 => "11111101",31954 => "01000001",31955 => "01101100",31956 => "01000110",31957 => "11011000",31958 => "10011101",31959 => "01011110",31960 => "10000001",31961 => "11110110",31962 => "10100010",31963 => "00000111",31964 => "01101011",31965 => "10010110",31966 => "01111001",31967 => "01010000",31968 => "11000000",31969 => "10000100",31970 => "01111000",31971 => "01000110",31972 => "10001000",31973 => "00100100",31974 => "11100111",31975 => "00010101",31976 => "01110110",31977 => "00001100",31978 => "10010010",31979 => "10001101",31980 => "10001011",31981 => "00111000",31982 => "10101000",31983 => "01111000",31984 => "01110101",31985 => "00101001",31986 => "00111000",31987 => "00001111",31988 => "00000111",31989 => "01101110",31990 => "00011000",31991 => "10010001",31992 => "00100111",31993 => "01111000",31994 => "00001111",31995 => "00000001",31996 => "00011111",31997 => "10000011",31998 => "00110010",31999 => "00001110",32000 => "11111110",32001 => "01110001",32002 => "01011100",32003 => "01111110",32004 => "00011101",32005 => "00010011",32006 => "00011101",32007 => "01111000",32008 => "10001101",32009 => "01010110",32010 => "01110000",32011 => "10111010",32012 => "10111011",32013 => "00010000",32014 => "01100110",32015 => "11100011",32016 => "00111001",32017 => "11011001",32018 => "01100011",32019 => "01011011",32020 => "01001011",32021 => "01001110",32022 => "11111101",32023 => "11011000",32024 => "01000110",32025 => "00010111",32026 => "01000010",32027 => "00110000",32028 => "10111011",32029 => "11100001",32030 => "00011110",32031 => "01000101",32032 => "11001101",32033 => "01001100",32034 => "11010010",32035 => "11110000",32036 => "11110101",32037 => "10001110",32038 => "00100110",32039 => "01101101",32040 => "00001011",32041 => "11101100",32042 => "10001101",32043 => "00110111",32044 => "01100110",32045 => "01101111",32046 => "10000010",32047 => "01100100",32048 => "11110010",32049 => "10111100",32050 => "00101110",32051 => "00101010",32052 => "10100001",32053 => "01101110",32054 => "00011111",32055 => "00001000",32056 => "01100001",32057 => "10001101",32058 => "00001100",32059 => "11110110",32060 => "11000010",32061 => "01001011",32062 => "00101111",32063 => "10010110",32064 => "00101011",32065 => "00101101",32066 => "00001001",32067 => "00111110",32068 => "01000111",32069 => "11001011",32070 => "00111000",32071 => "10110111",32072 => "00011110",32073 => "00000100",32074 => "11101110",32075 => "11111100",32076 => "10001000",32077 => "10001110",32078 => "01110110",32079 => "01100110",32080 => "01100110",32081 => "00000111",32082 => "01000010",32083 => "00000001",32084 => "01110011",32085 => "10011011",32086 => "00111100",32087 => "01001100",32088 => "01001001",32089 => "00101101",32090 => "00101111",32091 => "00000010",32092 => "00010101",32093 => "01010011",32094 => "10100111",32095 => "10001101",32096 => "00101001",32097 => "11101110",32098 => "00110011",32099 => "11001010",32100 => "11110001",32101 => "01101001",32102 => "11111000",32103 => "10011010",32104 => "00001101",32105 => "01100111",32106 => "01101011",32107 => "10101100",32108 => "10100100",32109 => "01110001",32110 => "11010000",32111 => "01110000",32112 => "10111101",32113 => "11110101",32114 => "11110010",32115 => "00001100",32116 => "00101001",32117 => "01101000",32118 => "00100101",32119 => "00110101",32120 => "01011111",32121 => "11011111",32122 => "11111111",32123 => "01100001",32124 => "11110011",32125 => "11110011",32126 => "01110010",32127 => "00001010",32128 => "10001011",32129 => "11001101",32130 => "01111010",32131 => "11100000",32132 => "10000101",32133 => "01110111",32134 => "11101101",32135 => "10100010",32136 => "01110010",32137 => "11101001",32138 => "10110100",32139 => "00011001",32140 => "11000010",32141 => "11000100",32142 => "00010101",32143 => "01000101",32144 => "00111000",32145 => "00111000",32146 => "00100011",32147 => "11111001",32148 => "01000001",32149 => "01111101",32150 => "01110110",32151 => "10001000",32152 => "10111001",32153 => "10011001",32154 => "10011000",32155 => "00111110",32156 => "11011010",32157 => "00010010",32158 => "01000000",32159 => "11011100",32160 => "11001110",32161 => "10011000",32162 => "11001011",32163 => "01100101",32164 => "10000000",32165 => "00011000",32166 => "01010001",32167 => "01011111",32168 => "00010001",32169 => "11100011",32170 => "00101011",32171 => "11000010",32172 => "11100010",32173 => "00010100",32174 => "01110000",32175 => "01101110",32176 => "01010000",32177 => "10011101",32178 => "00000100",32179 => "00001100",32180 => "11010001",32181 => "10001001",32182 => "10000101",32183 => "10111111",32184 => "11010101",32185 => "00000000",32186 => "10000001",32187 => "00110100",32188 => "11001000",32189 => "10100110",32190 => "01100011",32191 => "01101111",32192 => "01000010",32193 => "01001110",32194 => "00000001",32195 => "00001110",32196 => "10010000",32197 => "10110001",32198 => "11011010",32199 => "10000110",32200 => "11111011",32201 => "11001111",32202 => "01111100",32203 => "00010100",32204 => "11101001",32205 => "01101101",32206 => "01101111",32207 => "10101100",32208 => "00110110",32209 => "01000001",32210 => "00110100",32211 => "11001000",32212 => "10010000",32213 => "00011111",32214 => "10000010",32215 => "01100110",32216 => "00100010",32217 => "11111111",32218 => "01010001",32219 => "00010001",32220 => "10111101",32221 => "10001011",32222 => "10001111",32223 => "11011000",32224 => "11111011",32225 => "11110000",32226 => "01010011",32227 => "10100011",32228 => "10001011",32229 => "11001101",32230 => "01110010",32231 => "00011111",32232 => "01010100",32233 => "11100111",32234 => "00110111",32235 => "00110000",32236 => "11100101",32237 => "11100111",32238 => "11100101",32239 => "00111110",32240 => "00111101",32241 => "00100000",32242 => "01010001",32243 => "11010100",32244 => "10011010",32245 => "10010110",32246 => "10110110",32247 => "11000111",32248 => "00000001",32249 => "11000100",32250 => "11011100",32251 => "00110110",32252 => "01000101",32253 => "00001001",32254 => "01110001",32255 => "01101000",32256 => "00110000",32257 => "10100110",32258 => "11100101",32259 => "00111101",32260 => "10001100",32261 => "11001001",32262 => "11111011",32263 => "11010001",32264 => "01101010",32265 => "01010010",32266 => "10000100",32267 => "10110101",32268 => "00101110",32269 => "01101110",32270 => "01001101",32271 => "10010011",32272 => "11101110",32273 => "01111001",32274 => "11001100",32275 => "01111010",32276 => "10100100",32277 => "11111110",32278 => "00101101",32279 => "01010001",32280 => "01110000",32281 => "01101101",32282 => "00010000",32283 => "01011000",32284 => "01110001",32285 => "00111100",32286 => "10001101",32287 => "00010001",32288 => "11011111",32289 => "10101110",32290 => "00101111",32291 => "11010110",32292 => "01001010",32293 => "11110111",32294 => "11011101",32295 => "11100110",32296 => "10000011",32297 => "00100111",32298 => "01000100",32299 => "00001000",32300 => "11111111",32301 => "00001001",32302 => "01110010",32303 => "00000000",32304 => "01010000",32305 => "00000101",32306 => "11001011",32307 => "11110000",32308 => "10100000",32309 => "01001101",32310 => "00001101",32311 => "01010000",32312 => "11011011",32313 => "11011101",32314 => "00100010",32315 => "11000110",32316 => "00101011",32317 => "10000110",32318 => "10001111",32319 => "11000100",32320 => "01101010",32321 => "00111110",32322 => "10101110",32323 => "01101101",32324 => "00010001",32325 => "10101000",32326 => "00001110",32327 => "11110110",32328 => "10000001",32329 => "11001111",32330 => "00000110",32331 => "01000101",32332 => "11000011",32333 => "01100010",32334 => "00111000",32335 => "00111111",32336 => "11111010",32337 => "10110110",32338 => "10011101",32339 => "00000110",32340 => "01111011",32341 => "00101100",32342 => "00000110",32343 => "10001001",32344 => "01100000",32345 => "10011000",32346 => "00001000",32347 => "00001001",32348 => "01011110",32349 => "11110111",32350 => "00110110",32351 => "01010001",32352 => "11111110",32353 => "10001100",32354 => "01000011",32355 => "10110011",32356 => "01110010",32357 => "00010010",32358 => "01100110",32359 => "01100000",32360 => "10101100",32361 => "11100011",32362 => "01000000",32363 => "00001001",32364 => "00001111",32365 => "00111100",32366 => "10101000",32367 => "10100110",32368 => "11000110",32369 => "11010101",32370 => "11111110",32371 => "00101100",32372 => "11100101",32373 => "01111111",32374 => "01000101",32375 => "11010000",32376 => "01100011",32377 => "01111011",32378 => "00010111",32379 => "11001001",32380 => "01010110",32381 => "11011110",32382 => "00101100",32383 => "01000001",32384 => "10110011",32385 => "11011010",32386 => "11111010",32387 => "00100111",32388 => "00001000",32389 => "00101000",32390 => "11000100",32391 => "01011111",32392 => "00111011",32393 => "00101111",32394 => "01100011",32395 => "10100101",32396 => "10111000",32397 => "11001001",32398 => "11001101",32399 => "11011011",32400 => "10010110",32401 => "01100111",32402 => "10101101",32403 => "10011101",32404 => "11111110",32405 => "11001101",32406 => "11001100",32407 => "00011010",32408 => "01001101",32409 => "01010110",32410 => "01100111",32411 => "10101010",32412 => "11111011",32413 => "11001100",32414 => "10100111",32415 => "10010111",32416 => "11000000",32417 => "10101000",32418 => "10111111",32419 => "01001101",32420 => "00001111",32421 => "10111101",32422 => "00100100",32423 => "10100110",32424 => "10100011",32425 => "01101001",32426 => "11000111",32427 => "11010111",32428 => "01000111",32429 => "10101001",32430 => "01010010",32431 => "11100001",32432 => "10011001",32433 => "10011000",32434 => "01110010",32435 => "11010011",32436 => "01011011",32437 => "00010000",32438 => "10111101",32439 => "10000010",32440 => "00111001",32441 => "01010101",32442 => "11101101",32443 => "11101101",32444 => "01001101",32445 => "01111001",32446 => "00001011",32447 => "10001110",32448 => "11101111",32449 => "01111111",32450 => "10111011",32451 => "01001010",32452 => "11110111",32453 => "00010110",32454 => "00111010",32455 => "01101101",32456 => "10101110",32457 => "11011001",32458 => "01001110",32459 => "10011011",32460 => "10101011",32461 => "00101111",32462 => "00010100",32463 => "01111101",32464 => "11101001",32465 => "10010001",32466 => "10111100",32467 => "10011011",32468 => "11110011",32469 => "11111001",32470 => "00001001",32471 => "00101100",32472 => "01101110",32473 => "01010001",32474 => "00101000",32475 => "01101111",32476 => "10011011",32477 => "01011000",32478 => "00101100",32479 => "01101100",32480 => "00000010",32481 => "00100101",32482 => "00110000",32483 => "11000011",32484 => "01011010",32485 => "10000101",32486 => "10110010",32487 => "00010001",32488 => "00110110",32489 => "01100011",32490 => "11011000",32491 => "11010011",32492 => "11001001",32493 => "00001010",32494 => "10101100",32495 => "11011000",32496 => "11001111",32497 => "11001010",32498 => "11010101",32499 => "11111000",32500 => "01110001",32501 => "00000111",32502 => "11111000",32503 => "10100100",32504 => "10101010",32505 => "11111000",32506 => "01010011",32507 => "00001011",32508 => "00101100",32509 => "01001001",32510 => "01000010",32511 => "01101011",32512 => "10100011",32513 => "00101110",32514 => "10000010",32515 => "00011010",32516 => "01110001",32517 => "01010111",32518 => "11001101",32519 => "11110010",32520 => "01111010",32521 => "11001101",32522 => "00100101",32523 => "11011001",32524 => "00111010",32525 => "10010000",32526 => "10001101",32527 => "11000000",32528 => "11101100",32529 => "10011100",32530 => "10101011",32531 => "10111111",32532 => "10001111",32533 => "00111000",32534 => "01000001",32535 => "10100011",32536 => "11111110",32537 => "10111011",32538 => "01010111",32539 => "00100010",32540 => "11000110",32541 => "10100100",32542 => "01101111",32543 => "00110010",32544 => "10100101",32545 => "01101101",32546 => "11001010",32547 => "01010101",32548 => "10000100",32549 => "01010011",32550 => "10100001",32551 => "01110101",32552 => "10100101",32553 => "01001111",32554 => "10101000",32555 => "10110110",32556 => "01000001",32557 => "10100000",32558 => "10110100",32559 => "00111011",32560 => "10001011",32561 => "00000000",32562 => "10010110",32563 => "11110000",32564 => "00111100",32565 => "11001111",32566 => "10010011",32567 => "11111010",32568 => "01011101",32569 => "00011000",32570 => "10011011",32571 => "01100111",32572 => "01011011",32573 => "11010011",32574 => "10110011",32575 => "01100111",32576 => "11001101",32577 => "01101111",32578 => "10000011",32579 => "00101010",32580 => "11111000",32581 => "01000001",32582 => "01011111",32583 => "10000110",32584 => "01000011",32585 => "11110110",32586 => "10101010",32587 => "10000101",32588 => "01101111",32589 => "01101001",32590 => "10001110",32591 => "11010100",32592 => "01001011",32593 => "00110101",32594 => "10010001",32595 => "10100111",32596 => "10101101",32597 => "00000100",32598 => "11000111",32599 => "00110000",32600 => "01111010",32601 => "00001010",32602 => "00011010",32603 => "01000010",32604 => "11101101",32605 => "01100101",32606 => "00011000",32607 => "00100010",32608 => "00001000",32609 => "01001000",32610 => "10010110",32611 => "01010011",32612 => "00001100",32613 => "01100111",32614 => "11111000",32615 => "01100110",32616 => "10010011",32617 => "00011101",32618 => "10011000",32619 => "01100111",32620 => "00001101",32621 => "11100110",32622 => "01010110",32623 => "00100101",32624 => "10000001",32625 => "11111111",32626 => "10100101",32627 => "01110010",32628 => "01110011",32629 => "01100010",32630 => "01111101",32631 => "00100000",32632 => "11111011",32633 => "01110011",32634 => "01110000",32635 => "11000111",32636 => "01000100",32637 => "11001011",32638 => "11000111",32639 => "10000000",32640 => "01111100",32641 => "10010011",32642 => "10100000",32643 => "00001010",32644 => "00110001",32645 => "11010101",32646 => "00101110",32647 => "01111111",32648 => "01011000",32649 => "00011100",32650 => "11001010",32651 => "11100010",32652 => "10011001",32653 => "10101011",32654 => "11111010",32655 => "10110000",32656 => "10111111",32657 => "10010100",32658 => "00100001",32659 => "10100111",32660 => "00000110",32661 => "10111011",32662 => "01111111",32663 => "10001101",32664 => "10111000",32665 => "01010000",32666 => "00000100",32667 => "00010001",32668 => "01001000",32669 => "01111110",32670 => "11011111",32671 => "10110011",32672 => "00001100",32673 => "00001110",32674 => "00101110",32675 => "10101001",32676 => "00001101",32677 => "11011110",32678 => "00111110",32679 => "10110010",32680 => "01100001",32681 => "01010110",32682 => "10001101",32683 => "00110111",32684 => "10110101",32685 => "00100000",32686 => "11011110",32687 => "00010101",32688 => "10001010",32689 => "10000101",32690 => "11100001",32691 => "01011010",32692 => "11001010",32693 => "01100010",32694 => "00011000",32695 => "00100101",32696 => "11111111",32697 => "10100101",32698 => "01011010",32699 => "00100011",32700 => "00001011",32701 => "00010000",32702 => "11110011",32703 => "00010111",32704 => "10010101",32705 => "00010000",32706 => "10010001",32707 => "00011010",32708 => "10100001",32709 => "10110000",32710 => "00101100",32711 => "01101100",32712 => "10110101",32713 => "11101110",32714 => "00000001",32715 => "11001110",32716 => "00110011",32717 => "11010010",32718 => "01011011",32719 => "00000000",32720 => "00110010",32721 => "00111010",32722 => "00000101",32723 => "00010001",32724 => "10110010",32725 => "11110011",32726 => "01110010",32727 => "10010101",32728 => "10100111",32729 => "10010100",32730 => "01001110",32731 => "00000111",32732 => "01010100",32733 => "11101000",32734 => "10010111",32735 => "10001110",32736 => "00010110",32737 => "01010000",32738 => "11000110",32739 => "10111000",32740 => "10001100",32741 => "10001111",32742 => "11000100",32743 => "10001100",32744 => "01100011",32745 => "01101101",32746 => "10110000",32747 => "01001101",32748 => "11100101",32749 => "10011101",32750 => "00110110",32751 => "10100111",32752 => "01000011",32753 => "11010110",32754 => "10001010",32755 => "11011010",32756 => "11111001",32757 => "11110001",32758 => "01110010",32759 => "00010010",32760 => "10111010",32761 => "11011111",32762 => "00011000",32763 => "10001011",32764 => "10111101",32765 => "01111111",32766 => "00000000",32767 => "00011100",32768 => "01011001",32769 => "00101011",32770 => "11101110",32771 => "11100000",32772 => "01001001",32773 => "00101100",32774 => "10001000",32775 => "11000101",32776 => "01010101",32777 => "00001111",32778 => "11100110",32779 => "11111100",32780 => "11000100",32781 => "00010010",32782 => "10101001",32783 => "01100110",32784 => "00001100",32785 => "11101100",32786 => "10001100",32787 => "11100011",32788 => "00100100",32789 => "11010011",32790 => "01101100",32791 => "01111111",32792 => "01001011",32793 => "01100010",32794 => "10000100",32795 => "01011101",32796 => "00101111",32797 => "10000010",32798 => "01111001",32799 => "01011000",32800 => "11101100",32801 => "10111001",32802 => "10011001",32803 => "01000101",32804 => "00000011",32805 => "01111110",32806 => "01000011",32807 => "00011100",32808 => "01101110",32809 => "00001101",32810 => "00111011",32811 => "10011100",32812 => "00110011",32813 => "00111000",32814 => "11000110",32815 => "11110001",32816 => "01011010",32817 => "01001111",32818 => "10111111",32819 => "11000111",32820 => "11000100",32821 => "00011001",32822 => "10100100",32823 => "11011110",32824 => "01101011",32825 => "11110001",32826 => "01011001",32827 => "00001000",32828 => "00011000",32829 => "01011101",32830 => "01010010",32831 => "10110101",32832 => "00110101",32833 => "01111010",32834 => "01011111",32835 => "01101000",32836 => "01010111",32837 => "11010111",32838 => "01010000",32839 => "11000111",32840 => "00111011",32841 => "01110000",32842 => "00100101",32843 => "01100010",32844 => "01001110",32845 => "11101001",32846 => "11010011",32847 => "00001011",32848 => "00100010",32849 => "00001110",32850 => "11110101",32851 => "10111111",32852 => "10110110",32853 => "10001101",32854 => "00011111",32855 => "00001110",32856 => "01101011",32857 => "00000010",32858 => "10010011",32859 => "10011010",32860 => "00110010",32861 => "10101011",32862 => "11110101",32863 => "11000101",32864 => "10011010",32865 => "11001110",32866 => "00010000",32867 => "01101111",32868 => "11001000",32869 => "11101111",32870 => "00000110",32871 => "01010000",32872 => "01001100",32873 => "00011011",32874 => "10101011",32875 => "11001000",32876 => "11111111",32877 => "11100110",32878 => "11011110",32879 => "10111011",32880 => "01001000",32881 => "10101010",32882 => "00101111",32883 => "00011001",32884 => "00100110",32885 => "10111111",32886 => "11000011",32887 => "10001010",32888 => "01000100",32889 => "00000111",32890 => "10111110",32891 => "11010001",32892 => "11010100",32893 => "10101011",32894 => "01101100",32895 => "10000101",32896 => "01000000",32897 => "10111100",32898 => "10000101",32899 => "11001010",32900 => "11011111",32901 => "00010010",32902 => "10110000",32903 => "11000101",32904 => "10011010",32905 => "01111000",32906 => "01111111",32907 => "01010110",32908 => "11001111",32909 => "00110111",32910 => "11011110",32911 => "00001011",32912 => "00011111",32913 => "10101100",32914 => "11011110",32915 => "00000101",32916 => "01011111",32917 => "00100111",32918 => "11111100",32919 => "00000000",32920 => "10011000",32921 => "11100111",32922 => "01111010",32923 => "01010101",32924 => "10101101",32925 => "01101111",32926 => "01000000",32927 => "10010100",32928 => "00000010",32929 => "10100100",32930 => "01110011",32931 => "11110000",32932 => "00000100",32933 => "11010000",32934 => "10110111",32935 => "11100110",32936 => "01011111",32937 => "01100000",32938 => "10010001",32939 => "11011110",32940 => "01111010",32941 => "10111010",32942 => "10000110",32943 => "10101101",32944 => "11010001",32945 => "10100000",32946 => "01001111",32947 => "11101111",32948 => "10010111",32949 => "11101110",32950 => "11011100",32951 => "01001000",32952 => "11001000",32953 => "11010100",32954 => "11011001",32955 => "10000111",32956 => "00101010",32957 => "10011101",32958 => "10111000",32959 => "00001001",32960 => "01010111",32961 => "10100100",32962 => "10000101",32963 => "01100010",32964 => "01101111",32965 => "11101001",32966 => "11010111",32967 => "10101010",32968 => "10100111",32969 => "10100100",32970 => "01011011",32971 => "11011010",32972 => "11000001",32973 => "10100111",32974 => "01011000",32975 => "01110011",32976 => "11011011",32977 => "11110101",32978 => "10011001",32979 => "00010001",32980 => "10001101",32981 => "00101001",32982 => "10001001",32983 => "10000001",32984 => "10001111",32985 => "01100100",32986 => "10000001",32987 => "10111101",32988 => "11101000",32989 => "01110000",32990 => "00010001",32991 => "00111101",32992 => "01101101",32993 => "11101010",32994 => "11100010",32995 => "01111111",32996 => "01111001",32997 => "00010000",32998 => "11111010",32999 => "00111000",33000 => "00110101",33001 => "00101101",33002 => "00111110",33003 => "01100011",33004 => "10100000",33005 => "00101110",33006 => "00101001",33007 => "11100011",33008 => "10000110",33009 => "10011001",33010 => "10111100",33011 => "10110001",33012 => "11100100",33013 => "00010111",33014 => "11100110",33015 => "10011010",33016 => "11111010",33017 => "10011010",33018 => "01010110",33019 => "01010101",33020 => "11100011",33021 => "01010100",33022 => "10110111",33023 => "00101000",33024 => "10000000",33025 => "00000000",33026 => "01000101",33027 => "00100010",33028 => "00111010",33029 => "11000010",33030 => "11011110",33031 => "00111010",33032 => "11000001",33033 => "10011101",33034 => "00011101",33035 => "00101001",33036 => "01010111",33037 => "11110011",33038 => "10001110",33039 => "10101110",33040 => "10010111",33041 => "10110010",33042 => "11011100",33043 => "10111100",33044 => "10110000",33045 => "10001000",33046 => "10001111",33047 => "10110110",33048 => "11001000",33049 => "00011001",33050 => "10010011",33051 => "00001110",33052 => "01110000",33053 => "11111000",33054 => "11000111",33055 => "10000100",33056 => "11000000",33057 => "01110100",33058 => "10011011",33059 => "01011101",33060 => "00110001",33061 => "00101001",33062 => "10010101",33063 => "01010110",33064 => "00011100",33065 => "11000000",33066 => "00101100",33067 => "10001001",33068 => "11101001",33069 => "10101101",33070 => "00100001",33071 => "11111010",33072 => "10011001",33073 => "10011010",33074 => "11010000",33075 => "10000110",33076 => "01111100",33077 => "00011110",33078 => "11110010",33079 => "10100001",33080 => "10100100",33081 => "11111100",33082 => "11000110",33083 => "11011000",33084 => "10011011",33085 => "10001000",33086 => "11110011",33087 => "10111101",33088 => "10011111",33089 => "10001011",33090 => "11011011",33091 => "00111100",33092 => "10111111",33093 => "11101111",33094 => "10101010",33095 => "10010000",33096 => "11001001",33097 => "11101100",33098 => "11011010",33099 => "00001000",33100 => "11100110",33101 => "10101100",33102 => "11000001",33103 => "00111001",33104 => "10000111",33105 => "11000101",33106 => "11010111",33107 => "00011101",33108 => "00010000",33109 => "10101101",33110 => "11001100",33111 => "11011101",33112 => "10000010",33113 => "11000000",33114 => "10011010",33115 => "00110101",33116 => "01110100",33117 => "01100100",33118 => "10011001",33119 => "00010101",33120 => "01100101",33121 => "01111000",33122 => "11101011",33123 => "10000010",33124 => "11001110",33125 => "11001110",33126 => "01100000",33127 => "11101110",33128 => "11011110",33129 => "00000101",33130 => "01011010",33131 => "01011101",33132 => "10011101",33133 => "10110110",33134 => "10101010",33135 => "11110101",33136 => "11010011",33137 => "10110001",33138 => "00110110",33139 => "01111010",33140 => "01000011",33141 => "11100101",33142 => "10110000",33143 => "10100011",33144 => "11010100",33145 => "10111101",33146 => "01001111",33147 => "11001011",33148 => "10010100",33149 => "11111101",33150 => "11001111",33151 => "00000000",33152 => "00010111",33153 => "00011100",33154 => "01100111",33155 => "10000110",33156 => "10110010",33157 => "01010001",33158 => "00111101",33159 => "10010000",33160 => "01110001",33161 => "11111000",33162 => "10010100",33163 => "01110111",33164 => "11011001",33165 => "11000001",33166 => "01111101",33167 => "11100010",33168 => "01111011",33169 => "10011100",33170 => "10000100",33171 => "11001100",33172 => "00011010",33173 => "00001010",33174 => "11000010",33175 => "01001100",33176 => "00010100",33177 => "00101101",33178 => "11100111",33179 => "10101101",33180 => "11100010",33181 => "10111111",33182 => "11001111",33183 => "10000110",33184 => "11001000",33185 => "01010011",33186 => "11110111",33187 => "10111111",33188 => "11011001",33189 => "01100100",33190 => "11000101",33191 => "11011111",33192 => "00011011",33193 => "10111101",33194 => "01000111",33195 => "10110101",33196 => "00100010",33197 => "11101010",33198 => "01001011",33199 => "01101010",33200 => "01011111",33201 => "11101001",33202 => "10101011",33203 => "10001010",33204 => "11011111",33205 => "00101110",33206 => "00110001",33207 => "01001000",33208 => "11110000",33209 => "11001111",33210 => "01001111",33211 => "10000110",33212 => "01010000",33213 => "00110100",33214 => "01000000",33215 => "11101110",33216 => "10101110",33217 => "00000101",33218 => "01000100",33219 => "01100011",33220 => "10001000",33221 => "00011101",33222 => "01110001",33223 => "01000110",33224 => "01100011",33225 => "11110100",33226 => "00001001",33227 => "11111011",33228 => "10000110",33229 => "00110001",33230 => "11110000",33231 => "01111101",33232 => "11000111",33233 => "11100000",33234 => "11111011",33235 => "00110010",33236 => "11100000",33237 => "11000011",33238 => "10110111",33239 => "10101010",33240 => "10011000",33241 => "00101101",33242 => "00101000",33243 => "01001001",33244 => "11010000",33245 => "10111100",33246 => "11110110",33247 => "00111101",33248 => "00011010",33249 => "00001100",33250 => "01111010",33251 => "00000110",33252 => "00001101",33253 => "10100101",33254 => "00010110",33255 => "10110010",33256 => "10110101",33257 => "00001110",33258 => "00111001",33259 => "10101110",33260 => "10000110",33261 => "11100001",33262 => "01111111",33263 => "10100000",33264 => "11111111",33265 => "11001110",33266 => "00000010",33267 => "01100001",33268 => "00010111",33269 => "00101110",33270 => "01010110",33271 => "01011001",33272 => "01000011",33273 => "00000000",33274 => "01011101",33275 => "00001001",33276 => "00101011",33277 => "11111101",33278 => "00111101",33279 => "10011010",33280 => "11101110",33281 => "01010010",33282 => "00110111",33283 => "11100011",33284 => "10001000",33285 => "10111010",33286 => "01010111",33287 => "11001101",33288 => "10000111",33289 => "00001110",33290 => "10011101",33291 => "01110101",33292 => "01100000",33293 => "10010101",33294 => "11111100",33295 => "01101010",33296 => "01111101",33297 => "10001110",33298 => "00011111",33299 => "01010110",33300 => "11111101",33301 => "00110111",33302 => "01100010",33303 => "10110011",33304 => "10101010",33305 => "11110110",33306 => "11111110",33307 => "10111010",33308 => "00000111",33309 => "11100100",33310 => "01101101",33311 => "01100000",33312 => "01101101",33313 => "01111111",33314 => "11010001",33315 => "11001110",33316 => "01101010",33317 => "00011110",33318 => "01110000",33319 => "10111001",33320 => "01111101",33321 => "01100011",33322 => "10100110",33323 => "01111010",33324 => "11101100",33325 => "01011110",33326 => "00111100",33327 => "01111110",33328 => "11101000",33329 => "01110110",33330 => "01011111",33331 => "00000111",33332 => "10011000",33333 => "00010111",33334 => "10010001",33335 => "00110100",33336 => "10111011",33337 => "01111101",33338 => "00100001",33339 => "00101111",33340 => "11001100",33341 => "10100010",33342 => "01010111",33343 => "11100111",33344 => "01110000",33345 => "00000010",33346 => "01001110",33347 => "00010010",33348 => "11101001",33349 => "10011001",33350 => "10011100",33351 => "11100000",33352 => "11111001",33353 => "10100011",33354 => "11101111",33355 => "11011001",33356 => "00101001",33357 => "00110110",33358 => "10111110",33359 => "00010011",33360 => "10011000",33361 => "01100000",33362 => "10010001",33363 => "10111011",33364 => "01010011",33365 => "11001100",33366 => "10011011",33367 => "11011000",33368 => "00010000",33369 => "00011011",33370 => "00000010",33371 => "11001111",33372 => "11100101",33373 => "00101000",33374 => "00101111",33375 => "00010100",33376 => "11010001",33377 => "00111110",33378 => "10100001",33379 => "00101000",33380 => "00101100",33381 => "01111001",33382 => "10000000",33383 => "00010110",33384 => "10001001",33385 => "11001001",33386 => "00110001",33387 => "00000110",33388 => "10010001",33389 => "10110100",33390 => "00011110",33391 => "00110100",33392 => "11110110",33393 => "01110011",33394 => "11110110",33395 => "11111100",33396 => "10100101",33397 => "11101000",33398 => "00011101",33399 => "00001101",33400 => "01010110",33401 => "11110010",33402 => "11011010",33403 => "01110100",33404 => "10101001",33405 => "01100111",33406 => "11110110",33407 => "01001001",33408 => "10100101",33409 => "01010000",33410 => "01000101",33411 => "01000110",33412 => "11011110",33413 => "00011100",33414 => "10011101",33415 => "10010110",33416 => "01111100",33417 => "10101010",33418 => "10000101",33419 => "00100101",33420 => "11011110",33421 => "10101111",33422 => "10011010",33423 => "10011111",33424 => "00101101",33425 => "00001000",33426 => "01110000",33427 => "10000010",33428 => "11111000",33429 => "00001010",33430 => "10001010",33431 => "01110000",33432 => "11011110",33433 => "01001111",33434 => "10111111",33435 => "01001101",33436 => "11110111",33437 => "01000110",33438 => "01100000",33439 => "01011010",33440 => "11100111",33441 => "11010110",33442 => "00000000",33443 => "11100000",33444 => "10110011",33445 => "10001011",33446 => "01100110",33447 => "01001100",33448 => "00010000",33449 => "10110011",33450 => "11101000",33451 => "01110010",33452 => "01101100",33453 => "10111011",33454 => "10100111",33455 => "10100011",33456 => "00101110",33457 => "10110000",33458 => "11100010",33459 => "01110010",33460 => "10110110",33461 => "11101010",33462 => "01011000",33463 => "11111111",33464 => "01001101",33465 => "10000011",33466 => "11011111",33467 => "00100001",33468 => "01101100",33469 => "11100111",33470 => "11111110",33471 => "10110011",33472 => "11111000",33473 => "00110111",33474 => "11011110",33475 => "00111100",33476 => "10000101",33477 => "00110111",33478 => "01100100",33479 => "11111101",33480 => "11001110",33481 => "10111011",33482 => "01110101",33483 => "00011110",33484 => "01001001",33485 => "01101101",33486 => "00111100",33487 => "10000010",33488 => "00001100",33489 => "10001000",33490 => "00110101",33491 => "10000001",33492 => "00101011",33493 => "01011100",33494 => "10001001",33495 => "10001100",33496 => "11111111",33497 => "11100100",33498 => "01100111",33499 => "11001001",33500 => "00001110",33501 => "10101000",33502 => "10110010",33503 => "11000111",33504 => "01111111",33505 => "10100111",33506 => "01111100",33507 => "11101110",33508 => "00010101",33509 => "11010010",33510 => "11100110",33511 => "01000101",33512 => "00000011",33513 => "00010110",33514 => "10000011",33515 => "01011101",33516 => "01000001",33517 => "11101000",33518 => "11101011",33519 => "01111000",33520 => "10010000",33521 => "11101001",33522 => "00011011",33523 => "00011100",33524 => "00010111",33525 => "11111001",33526 => "10110101",33527 => "11110111",33528 => "01000000",33529 => "00000001",33530 => "01111101",33531 => "11101100",33532 => "10000110",33533 => "01011010",33534 => "11100001",33535 => "01000100",33536 => "10001111",33537 => "00011101",33538 => "01100010",33539 => "11110011",33540 => "11111100",33541 => "00100011",33542 => "10000000",33543 => "11010100",33544 => "01101101",33545 => "01001110",33546 => "01001110",33547 => "00011111",33548 => "10000001",33549 => "10000000",33550 => "01101110",33551 => "01011000",33552 => "01010011",33553 => "01101010",33554 => "01001000",33555 => "00000101",33556 => "10000000",33557 => "01010001",33558 => "11100011",33559 => "11001011",33560 => "11111111",33561 => "10111010",33562 => "11100001",33563 => "11110001",33564 => "11111110",33565 => "10100100",33566 => "10001011",33567 => "11110101",33568 => "10000011",33569 => "10100101",33570 => "11000101",33571 => "11001110",33572 => "01000100",33573 => "11011101",33574 => "00011110",33575 => "00101001",33576 => "11010010",33577 => "01110001",33578 => "00000011",33579 => "01101101",33580 => "01011111",33581 => "10101010",33582 => "10001111",33583 => "10011010",33584 => "01000110",33585 => "00100110",33586 => "00101000",33587 => "10101100",33588 => "01011111",33589 => "01110111",33590 => "01001101",33591 => "01000110",33592 => "11101100",33593 => "10001110",33594 => "01101101",33595 => "11011000",33596 => "10101011",33597 => "10011111",33598 => "11111000",33599 => "11101110",33600 => "00110101",33601 => "11100000",33602 => "01010100",33603 => "01001110",33604 => "01010001",33605 => "10101011",33606 => "01010000",33607 => "01010000",33608 => "00001011",33609 => "10010111",33610 => "00101001",33611 => "00100001",33612 => "11101101",33613 => "10110001",33614 => "11011110",33615 => "00111100",33616 => "01111111",33617 => "00001110",33618 => "01000110",33619 => "00100110",33620 => "01111100",33621 => "00110011",33622 => "00111010",33623 => "11011111",33624 => "10111101",33625 => "10110001",33626 => "00111111",33627 => "01011110",33628 => "10111011",33629 => "11100110",33630 => "11000010",33631 => "00001010",33632 => "11110111",33633 => "01111010",33634 => "11100111",33635 => "10101100",33636 => "11110011",33637 => "00010111",33638 => "01111000",33639 => "00000110",33640 => "11100001",33641 => "01000000",33642 => "00110000",33643 => "01011101",33644 => "01100010",33645 => "11001011",33646 => "11010000",33647 => "00011101",33648 => "01010100",33649 => "00010110",33650 => "11010101",33651 => "11001001",33652 => "00100001",33653 => "01110100",33654 => "10011100",33655 => "10011010",33656 => "11001111",33657 => "11100110",33658 => "01001010",33659 => "10000010",33660 => "11101101",33661 => "01000101",33662 => "01000010",33663 => "10010010",33664 => "01010100",33665 => "11110000",33666 => "00111110",33667 => "10010011",33668 => "01000111",33669 => "01110000",33670 => "00011011",33671 => "01010111",33672 => "10010101",33673 => "01010100",33674 => "00110011",33675 => "10101100",33676 => "01110001",33677 => "11110111",33678 => "00110101",33679 => "10011100",33680 => "10111111",33681 => "00111001",33682 => "11001011",33683 => "00010001",33684 => "10000010",33685 => "11011001",33686 => "00111010",33687 => "00000001",33688 => "10111000",33689 => "11011001",33690 => "00001111",33691 => "11110000",33692 => "10100100",33693 => "11111110",33694 => "10011011",33695 => "10100111",33696 => "11101100",33697 => "10001011",33698 => "10110000",33699 => "01110101",33700 => "00101011",33701 => "01000100",33702 => "01110000",33703 => "01100001",33704 => "10000110",33705 => "01111100",33706 => "10111000",33707 => "11000110",33708 => "01010110",33709 => "01010000",33710 => "00010101",33711 => "10110110",33712 => "11100001",33713 => "11000011",33714 => "11110111",33715 => "11100001",33716 => "10100000",33717 => "01001101",33718 => "10010101",33719 => "01011110",33720 => "01011111",33721 => "01101101",33722 => "01010000",33723 => "00011010",33724 => "01001100",33725 => "00000110",33726 => "10001010",33727 => "00010111",33728 => "10010100",33729 => "01010000",33730 => "01001101",33731 => "01010110",33732 => "10001001",33733 => "10100101",33734 => "01010110",33735 => "11001001",33736 => "00110011",33737 => "01100100",33738 => "11000100",33739 => "10100100",33740 => "11001101",33741 => "10101101",33742 => "01110010",33743 => "11011011",33744 => "10010001",33745 => "01000101",33746 => "00100010",33747 => "11011011",33748 => "00011100",33749 => "10011100",33750 => "10110011",33751 => "11100101",33752 => "10000101",33753 => "01100111",33754 => "01111100",33755 => "10010100",33756 => "01111011",33757 => "10011100",33758 => "11011011",33759 => "11111010",33760 => "10111011",33761 => "01011100",33762 => "00011000",33763 => "01000001",33764 => "11001000",33765 => "01111001",33766 => "10001000",33767 => "10101100",33768 => "10101001",33769 => "00001001",33770 => "10101100",33771 => "01001101",33772 => "10110001",33773 => "01110110",33774 => "10100111",33775 => "10111010",33776 => "00011001",33777 => "10010000",33778 => "01110100",33779 => "11101011",33780 => "00111100",33781 => "10010001",33782 => "11110101",33783 => "01000001",33784 => "01000110",33785 => "11001000",33786 => "01010001",33787 => "00010100",33788 => "10011010",33789 => "01110001",33790 => "11001000",33791 => "00100011",33792 => "00011110",33793 => "10010110",33794 => "00001000",33795 => "01111001",33796 => "11111001",33797 => "11001000",33798 => "11010001",33799 => "00011101",33800 => "10000101",33801 => "11101100",33802 => "00001101",33803 => "00010000",33804 => "01001111",33805 => "01110001",33806 => "00011001",33807 => "01001100",33808 => "00010101",33809 => "11011111",33810 => "11011001",33811 => "01001100",33812 => "10010011",33813 => "10111010",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "10000100" report "FAIL high bits" severity failure;
assert RAM(0) = "00010101" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
