 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01111100",3 => "10000010",4 => "01100000",5 => "01110001",6 => "01010101",7 => "10011101",8 => "11101110",9 => "01011011",10 => "01101000",11 => "10001110",12 => "00111011",13 => "11010000",14 => "10101100",15 => "11000010",16 => "11100111",17 => "01111011",18 => "00001111",19 => "00000010",20 => "01001111",21 => "10111110",22 => "01011010",23 => "11010110",24 => "01011010",25 => "01110001",26 => "01000001",27 => "10000101",28 => "01111011",29 => "00011101",30 => "00010101",31 => "00101110",32 => "11000010",33 => "01111110",34 => "01110001",35 => "11110110",36 => "10011111",37 => "10011011",38 => "01001001",39 => "11011001",40 => "01001001",41 => "11010001",42 => "01100110",43 => "11110011",44 => "10001110",45 => "00010101",46 => "01100111",47 => "10110010",48 => "10000010",49 => "11101000",50 => "10111100",51 => "00011100",52 => "00001011",53 => "10011001",54 => "00101100",55 => "10111100",56 => "10100110",57 => "01010101",58 => "01111100",59 => "10101101",60 => "10101110",61 => "00010110",62 => "11110100",63 => "00110010",64 => "01100001",65 => "00111100",66 => "00010101",67 => "00111110",68 => "10011110",69 => "01001000",70 => "01011011",71 => "01111001",72 => "01111111",73 => "10111101",74 => "10010001",75 => "01100010",76 => "01101101",77 => "11000011",78 => "01111110",79 => "01111100",80 => "00011000",81 => "10011001",82 => "01100101",83 => "01100111",84 => "01101011",85 => "01000000",86 => "00010101",87 => "11010011",88 => "00110101",89 => "00010100",90 => "11000101",91 => "11000111",92 => "11000100",93 => "01100011",94 => "10101100",95 => "01000001",96 => "10010111",97 => "11011011",98 => "01010000",99 => "11000101",100 => "01011100",101 => "11000100",102 => "10000100",103 => "01101110",104 => "10111101",105 => "11111101",106 => "01110000",107 => "00100010",108 => "10001110",109 => "11010011",110 => "10010100",111 => "10101010",112 => "11001010",113 => "01111110",114 => "11111011",115 => "11000000",116 => "10101011",117 => "00101101",118 => "11010010",119 => "11110011",120 => "10001101",121 => "10000111",122 => "11010000",123 => "10001111",124 => "01010001",125 => "01111101",126 => "10100010",127 => "01100111",128 => "00010011",129 => "11100111",130 => "01100101",131 => "00011001",132 => "10001000",133 => "01110111",134 => "11000101",135 => "11001000",136 => "00011001",137 => "01111100",138 => "10001101",139 => "01000100",140 => "11101001",141 => "01101011",142 => "10101101",143 => "11011001",144 => "11100001",145 => "00100110",146 => "01101011",147 => "10100001",148 => "10000010",149 => "01001000",150 => "00010010",151 => "10000001",152 => "10101000",153 => "10110001",154 => "01101100",155 => "10100010",156 => "11110010",157 => "01110010",158 => "00101000",159 => "10010111",160 => "11110111",161 => "00001000",162 => "11001011",163 => "11111101",164 => "11111001",165 => "01100101",166 => "01001101",167 => "00010110",168 => "01010100",169 => "01001011",170 => "10111010",171 => "10001111",172 => "01111110",173 => "10100001",174 => "10100101",175 => "00001001",176 => "11001111",177 => "01101011",178 => "10001001",179 => "10100101",180 => "01110111",181 => "00011010",182 => "01110011",183 => "00010010",184 => "00100100",185 => "11010111",186 => "10001101",187 => "10000010",188 => "10111000",189 => "00101101",190 => "00010011",191 => "10000000",192 => "00001011",193 => "10001000",194 => "11001100",195 => "11010000",196 => "01100011",197 => "01110110",198 => "10111111",199 => "10011011",200 => "00110000",201 => "11011001",202 => "01000000",203 => "11100011",204 => "01111001",205 => "01101110",206 => "01100010",207 => "11101101",208 => "10100100",209 => "10001000",210 => "11111000",211 => "00001010",212 => "01101000",213 => "11111111",214 => "10000110",215 => "10010101",216 => "00111011",217 => "01001110",218 => "01001101",219 => "01001100",220 => "10100001",221 => "01110101",222 => "00010000",223 => "10010001",224 => "10111000",225 => "10000100",226 => "01111000",227 => "00100100",228 => "10000011",229 => "10111111",230 => "10110100",231 => "11010001",232 => "01100101",233 => "10111011",234 => "00011100",235 => "11010111",236 => "10110110",237 => "10000110",238 => "00001100",239 => "01000000",240 => "01100011",241 => "01111001",242 => "00000101",243 => "01010111",244 => "00001100",245 => "01101011",246 => "11111010",247 => "01101110",248 => "01100101",249 => "01101101",250 => "11010100",251 => "01101000",252 => "01100100",253 => "11001000",254 => "00110111",255 => "11000000",256 => "10010000",257 => "10000110",258 => "10000100",259 => "01000001",260 => "11111101",261 => "01000001",262 => "01100000",263 => "10000010",264 => "00101000",265 => "00110111",266 => "10001100",267 => "01110000",268 => "10110000",269 => "11100100",270 => "11111111",271 => "01010000",272 => "00111011",273 => "00001110",274 => "00111000",275 => "10101010",276 => "11000011",277 => "00010000",278 => "00101111",279 => "00111011",280 => "00010111",281 => "01100011",282 => "10101011",283 => "00001101",284 => "00111010",285 => "01111111",286 => "11011010",287 => "10101111",288 => "00011110",289 => "10111110",290 => "01111000",291 => "10000000",292 => "01000010",293 => "10111000",294 => "00010110",295 => "10110101",296 => "11010101",297 => "10101011",298 => "10100010",299 => "11011110",300 => "00000111",301 => "11010001",302 => "00100000",303 => "10111100",304 => "11001000",305 => "00001010",306 => "00111111",307 => "00010100",308 => "00000010",309 => "11000000",310 => "10011001",311 => "11100111",312 => "00010111",313 => "00101001",314 => "00101000",315 => "10101101",316 => "00100110",317 => "01010100",318 => "10110001",319 => "10011001",320 => "11100101",321 => "10000110",322 => "00000010",323 => "00101011",324 => "11110001",325 => "00110111",326 => "01111001",327 => "01111010",328 => "10110110",329 => "01010101",330 => "00100010",331 => "10101110",332 => "01111101",333 => "11101101",334 => "00111000",335 => "01101100",336 => "01000000",337 => "01110001",338 => "11111110",339 => "01100001",340 => "00001000",341 => "11001000",342 => "01101011",343 => "10100001",344 => "11101100",345 => "00010011",346 => "11111000",347 => "10110010",348 => "11101000",349 => "11100100",350 => "10001111",351 => "00000111",352 => "01011100",353 => "00010011",354 => "01111111",355 => "00110011",356 => "11001000",357 => "01101101",358 => "01001000",359 => "10011001",360 => "10101111",361 => "11000011",362 => "00010010",363 => "11110001",364 => "11110101",365 => "01101101",366 => "00001000",367 => "11111110",368 => "00010000",369 => "01100010",370 => "10100100",371 => "01010010",372 => "01100011",373 => "01110101",374 => "10010100",375 => "01100001",376 => "10101100",377 => "01011100",378 => "01010010",379 => "00100111",380 => "11110100",381 => "11111100",382 => "10110100",383 => "10010010",384 => "01100111",385 => "11010011",386 => "10111100",387 => "10011110",388 => "01010111",389 => "01100111",390 => "01101011",391 => "10100010",392 => "11011010",393 => "10010110",394 => "10101101",395 => "10000001",396 => "00000010",397 => "01011101",398 => "01101111",399 => "01100111",400 => "11100111",401 => "11101010",402 => "11111110",403 => "01110111",404 => "00100000",405 => "00011101",406 => "01111000",407 => "00111111",408 => "11111011",409 => "00100101",410 => "01000010",411 => "10111110",412 => "01100101",413 => "00101111",414 => "10100000",415 => "01111111",416 => "01000100",417 => "10111101",418 => "10100110",419 => "00001010",420 => "00100101",421 => "10000001",422 => "10110010",423 => "11010000",424 => "10010001",425 => "01010111",426 => "01100110",427 => "00101001",428 => "00100101",429 => "00011111",430 => "11101011",431 => "01010000",432 => "11011111",433 => "10010111",434 => "11011101",435 => "10010110",436 => "10000100",437 => "01110110",438 => "10000111",439 => "11011110",440 => "00001011",441 => "01110011",442 => "00001100",443 => "01010100",444 => "00001011",445 => "00111001",446 => "11110110",447 => "01011111",448 => "10011000",449 => "00111011",450 => "10001110",451 => "10000111",452 => "00010010",453 => "10001010",454 => "11001000",455 => "00100100",456 => "01101101",457 => "10111011",458 => "00100001",459 => "00110000",460 => "10001010",461 => "01101110",462 => "00111100",463 => "11001001",464 => "10011000",465 => "11100001",466 => "11011011",467 => "01100110",468 => "00110011",469 => "10110111",470 => "01100110",471 => "11010111",472 => "11000010",473 => "10010001",474 => "00100011",475 => "10101011",476 => "10110100",477 => "11001010",478 => "10101000",479 => "11001110",480 => "11010001",481 => "01011010",482 => "00010011",483 => "11001000",484 => "00000010",485 => "11000010",486 => "11011011",487 => "10011011",488 => "01010000",489 => "10110110",490 => "01110100",491 => "00111111",492 => "00100110",493 => "11101000",494 => "10011000",495 => "11000000",496 => "01000100",497 => "01111111",498 => "10010110",499 => "10001001",500 => "01000011",501 => "11111001",502 => "10100110",503 => "10011010",504 => "00100111",505 => "11110111",506 => "10101100",507 => "11111001",508 => "11110111",509 => "11011011",510 => "10010110",511 => "01111111",512 => "00000111",513 => "10110101",514 => "10110110",515 => "00111000",516 => "11110011",517 => "01110110",518 => "00101011",519 => "10000110",520 => "11011101",521 => "01001001",522 => "00100010",523 => "11111010",524 => "11001101",525 => "10110001",526 => "00011110",527 => "11110100",528 => "11000011",529 => "10000100",530 => "00010001",531 => "10101001",532 => "01100101",533 => "01010001",534 => "00111001",535 => "01101111",536 => "01100000",537 => "01111110",538 => "11010001",539 => "10011101",540 => "01010010",541 => "10000001",542 => "11010001",543 => "01000101",544 => "01000101",545 => "10011011",546 => "00101110",547 => "11101001",548 => "10000011",549 => "11101111",550 => "00001001",551 => "00011110",552 => "11001001",553 => "10111000",554 => "00010011",555 => "01110100",556 => "00101001",557 => "10010101",558 => "10110100",559 => "00100111",560 => "11011100",561 => "11101000",562 => "11001010",563 => "00100010",564 => "01110100",565 => "00010001",566 => "10000110",567 => "00101010",568 => "00110010",569 => "01110010",570 => "11001101",571 => "00110101",572 => "11101110",573 => "10100000",574 => "01100000",575 => "10000101",576 => "11101000",577 => "10010101",578 => "01100110",579 => "11110010",580 => "10010000",581 => "11010100",582 => "01110000",583 => "00110100",584 => "11100001",585 => "00011101",586 => "10110111",587 => "10111111",588 => "01010100",589 => "11000001",590 => "11100101",591 => "10000000",592 => "11111100",593 => "11010010",594 => "01100111",595 => "10010001",596 => "00110111",597 => "01110100",598 => "01101011",599 => "11110010",600 => "01101000",601 => "00000111",602 => "11100010",603 => "11110111",604 => "11100111",605 => "11101101",606 => "00110010",607 => "00111100",608 => "10111011",609 => "11110111",610 => "00011011",611 => "01110110",612 => "00101000",613 => "01011010",614 => "10011100",615 => "01010100",616 => "10010101",617 => "00011110",618 => "01000101",619 => "10100011",620 => "11110101",621 => "10000111",622 => "00101100",623 => "11111010",624 => "10001100",625 => "11011110",626 => "11000000",627 => "10011010",628 => "10101111",629 => "00110000",630 => "11010001",631 => "11011010",632 => "01011110",633 => "10001010",634 => "10110011",635 => "00101010",636 => "01100111",637 => "00011110",638 => "01010011",639 => "00010111",640 => "00111110",641 => "10110000",642 => "01101011",643 => "00001111",644 => "00111110",645 => "10111111",646 => "01100101",647 => "10100111",648 => "10010111",649 => "00110111",650 => "00000010",651 => "01000101",652 => "10000100",653 => "01110000",654 => "10101101",655 => "00110101",656 => "11000000",657 => "10000001",658 => "01000110",659 => "10000010",660 => "01100001",661 => "10000100",662 => "01111010",663 => "01010100",664 => "11100001",665 => "11101001",666 => "10111010",667 => "11000100",668 => "01100110",669 => "01100000",670 => "11110100",671 => "00000101",672 => "10100000",673 => "01001111",674 => "01011000",675 => "01000011",676 => "10101110",677 => "11010101",678 => "01000001",679 => "00100001",680 => "01011110",681 => "01011100",682 => "10101000",683 => "01010010",684 => "01101101",685 => "10011001",686 => "11100001",687 => "11110001",688 => "11010000",689 => "01000111",690 => "10101101",691 => "11101001",692 => "01100111",693 => "01101000",694 => "01101111",695 => "00110101",696 => "10100100",697 => "01100000",698 => "10101101",699 => "10100110",700 => "10001001",701 => "01010110",702 => "00011000",703 => "10100011",704 => "10001000",705 => "01110000",706 => "10101100",707 => "00001110",708 => "11010110",709 => "11100000",710 => "10000001",711 => "00111101",712 => "01111101",713 => "11001010",714 => "01001101",715 => "11011010",716 => "11001010",717 => "11010100",718 => "00101100",719 => "10011101",720 => "00111000",721 => "01110110",722 => "00000111",723 => "00111001",724 => "00111111",725 => "11101010",726 => "01101001",727 => "11000011",728 => "00111111",729 => "01010111",730 => "10111101",731 => "10101000",732 => "10110010",733 => "00110001",734 => "01101100",735 => "01101001",736 => "10111000",737 => "11110000",738 => "01100110",739 => "10010011",740 => "01110100",741 => "00011011",742 => "00100110",743 => "01101101",744 => "00000111",745 => "00000010",746 => "01101101",747 => "00011111",748 => "00101101",749 => "10100111",750 => "00101010",751 => "11001000",752 => "00101101",753 => "00100100",754 => "01110010",755 => "01100110",756 => "10111100",757 => "01000100",758 => "11010111",759 => "11100110",760 => "11111101",761 => "00101101",762 => "10110000",763 => "11111011",764 => "00111100",765 => "00100000",766 => "00011111",767 => "10111111",768 => "01011100",769 => "01101000",770 => "01101111",771 => "00001111",772 => "00010101",773 => "11000111",774 => "10100000",775 => "10101111",776 => "10000001",777 => "00110000",778 => "00111101",779 => "10011010",780 => "10001000",781 => "00011100",782 => "10111101",783 => "01011001",784 => "11010111",785 => "00110011",786 => "01101000",787 => "10001101",788 => "11010110",789 => "11000000",790 => "11110100",791 => "11100101",792 => "00011000",793 => "10100110",794 => "10111110",795 => "10001101",796 => "10100010",797 => "01000111",798 => "01000100",799 => "00000001",800 => "00011111",801 => "10000100",802 => "01000111",803 => "10001010",804 => "01110101",805 => "10101101",806 => "00110100",807 => "11111111",808 => "10000110",809 => "11111101",810 => "00010010",811 => "10011111",812 => "10010011",813 => "10011100",814 => "00100100",815 => "00110111",816 => "10000111",817 => "10001001",818 => "11001001",819 => "10010101",820 => "11111110",821 => "10100010",822 => "11100110",823 => "10110000",824 => "01011000",825 => "00100000",826 => "00000101",827 => "01110001",828 => "10001001",829 => "11100101",830 => "01001000",831 => "01001110",832 => "01011100",833 => "00010101",834 => "10100000",835 => "11010100",836 => "10101011",837 => "11010011",838 => "01011111",839 => "11000111",840 => "11001000",841 => "10001011",842 => "10111110",843 => "00110100",844 => "11010110",845 => "00001100",846 => "11100001",847 => "10011101",848 => "00001011",849 => "01010100",850 => "11010011",851 => "01111111",852 => "01100011",853 => "00111011",854 => "00110000",855 => "01100000",856 => "00110011",857 => "10011101",858 => "00000000",859 => "00101010",860 => "01110100",861 => "00101010",862 => "11000110",863 => "10100100",864 => "01000010",865 => "10110001",866 => "00011011",867 => "10101101",868 => "00101000",869 => "01100101",870 => "10001001",871 => "11001010",872 => "10101110",873 => "01011101",874 => "10101100",875 => "01111110",876 => "01001110",877 => "11000010",878 => "11000010",879 => "01100010",880 => "00010000",881 => "01101000",882 => "00100001",883 => "11001011",884 => "11101110",885 => "10011100",886 => "11000000",887 => "01101011",888 => "00111111",889 => "00100100",890 => "01100100",891 => "10111110",892 => "00111111",893 => "01110101",894 => "10011010",895 => "00110000",896 => "11110110",897 => "11100100",898 => "01010101",899 => "01010010",900 => "01001111",901 => "11011000",902 => "11000001",903 => "11111011",904 => "11111000",905 => "00110100",906 => "11000010",907 => "10101111",908 => "00101110",909 => "00101010",910 => "11101110",911 => "10111111",912 => "10000100",913 => "00100001",914 => "11000010",915 => "00101000",916 => "00001010",917 => "10000000",918 => "01111111",919 => "00010011",920 => "11110110",921 => "11110100",922 => "10010000",923 => "00000010",924 => "11000001",925 => "00100011",926 => "00010110",927 => "01010001",928 => "11100001",929 => "11011110",930 => "01011111",931 => "11001111",932 => "10100010",933 => "10100011",934 => "10011001",935 => "00111000",936 => "10000000",937 => "11101000",938 => "10000001",939 => "00010111",940 => "01010010",941 => "11011111",942 => "00100101",943 => "10111010",944 => "01110110",945 => "00110111",946 => "01000010",947 => "11110001",948 => "10000000",949 => "11101010",950 => "11110101",951 => "01001101",952 => "10111010",953 => "11100110",954 => "11000111",955 => "01011111",956 => "01000111",957 => "01101000",958 => "01101001",959 => "11001101",960 => "11011100",961 => "01101110",962 => "10110011",963 => "10011110",964 => "00101101",965 => "10111111",966 => "11000100",967 => "10010100",968 => "01000010",969 => "10110110",970 => "01011110",971 => "01000100",972 => "00101000",973 => "00110111",974 => "10100000",975 => "01110111",976 => "01101101",977 => "01011110",978 => "00111001",979 => "10000111",980 => "00010010",981 => "00100001",982 => "11011001",983 => "10110010",984 => "00000111",985 => "01000111",986 => "11110010",987 => "00100000",988 => "10111111",989 => "11011101",990 => "10010100",991 => "11111011",992 => "01011001",993 => "11001000",994 => "01100111",995 => "11010000",996 => "01001110",997 => "01001101",998 => "01101111",999 => "00110001",1000 => "00010111",1001 => "11010101",1002 => "11010100",1003 => "10010000",1004 => "00000010",1005 => "01110101",1006 => "11000001",1007 => "01001101",1008 => "00010101",1009 => "01001111",1010 => "01011000",1011 => "01111001",1012 => "00010011",1013 => "01001101",1014 => "01000110",1015 => "11101101",1016 => "11100001",1017 => "01100001",1018 => "01000011",1019 => "01100001",1020 => "00010100",1021 => "10110101",1022 => "00011100",1023 => "01010010",1024 => "00011110",1025 => "01010101",1026 => "01001011",1027 => "11001100",1028 => "11000011",1029 => "11010010",1030 => "00100010",1031 => "10001100",1032 => "01101011",1033 => "11000001",1034 => "00011110",1035 => "01100101",1036 => "00101110",1037 => "11101010",1038 => "11010000",1039 => "11110111",1040 => "00000001",1041 => "10111011",1042 => "11011110",1043 => "01001010",1044 => "00111111",1045 => "01000101",1046 => "01111100",1047 => "11010010",1048 => "01001001",1049 => "00110101",1050 => "11001011",1051 => "10011110",1052 => "00111101",1053 => "00011000",1054 => "01011010",1055 => "11101100",1056 => "01001100",1057 => "11100010",1058 => "00001100",1059 => "01100101",1060 => "10111100",1061 => "11010010",1062 => "01001100",1063 => "01011100",1064 => "01000011",1065 => "01011001",1066 => "00010101",1067 => "00101110",1068 => "01011101",1069 => "01110011",1070 => "11001101",1071 => "00001110",1072 => "11101101",1073 => "10110001",1074 => "01101011",1075 => "11011100",1076 => "10011101",1077 => "00110011",1078 => "01110100",1079 => "11010000",1080 => "00101100",1081 => "01010011",1082 => "10010010",1083 => "00011100",1084 => "10001101",1085 => "00000110",1086 => "10111000",1087 => "10100100",1088 => "01000000",1089 => "00101010",1090 => "10011001",1091 => "11100110",1092 => "10101001",1093 => "11011100",1094 => "10101000",1095 => "11110100",1096 => "10011001",1097 => "01110100",1098 => "01110111",1099 => "00111001",1100 => "00101010",1101 => "11110000",1102 => "01001000",1103 => "01100100",1104 => "01001000",1105 => "10000001",1106 => "10010011",1107 => "00110001",1108 => "11101100",1109 => "10110001",1110 => "01101001",1111 => "11000011",1112 => "00100110",1113 => "01011000",1114 => "00111101",1115 => "01100111",1116 => "01001100",1117 => "01100100",1118 => "11110100",1119 => "00111011",1120 => "00000101",1121 => "01110100",1122 => "10011101",1123 => "10010011",1124 => "00011001",1125 => "00010010",1126 => "10101101",1127 => "10011111",1128 => "11111110",1129 => "10010011",1130 => "11011100",1131 => "10111011",1132 => "10010001",1133 => "10010111",1134 => "01111011",1135 => "00011001",1136 => "10010111",1137 => "01100101",1138 => "01101001",1139 => "01000000",1140 => "10111011",1141 => "01100100",1142 => "11110001",1143 => "01000111",1144 => "01110110",1145 => "01101010",1146 => "00010100",1147 => "01000111",1148 => "00010100",1149 => "01010000",1150 => "01000001",1151 => "01100110",1152 => "00010000",1153 => "01100001",1154 => "11000000",1155 => "11011010",1156 => "11110011",1157 => "10111001",1158 => "00101000",1159 => "10110000",1160 => "01101000",1161 => "10001001",1162 => "01101110",1163 => "11101100",1164 => "11100010",1165 => "10110111",1166 => "10001100",1167 => "01010111",1168 => "00000101",1169 => "00101110",1170 => "10111001",1171 => "10100000",1172 => "01111011",1173 => "10011101",1174 => "11110000",1175 => "11101010",1176 => "11111011",1177 => "11111100",1178 => "00111000",1179 => "00000000",1180 => "01011100",1181 => "11101101",1182 => "01001110",1183 => "10011110",1184 => "01000101",1185 => "00011111",1186 => "10011101",1187 => "10101111",1188 => "01001010",1189 => "11100111",1190 => "11010101",1191 => "01011111",1192 => "00100100",1193 => "11000100",1194 => "00110110",1195 => "01110010",1196 => "11010011",1197 => "01100101",1198 => "10000011",1199 => "00000101",1200 => "01110100",1201 => "10111101",1202 => "11011011",1203 => "11111100",1204 => "10111111",1205 => "00101101",1206 => "11100111",1207 => "00001001",1208 => "01000111",1209 => "01000101",1210 => "11011000",1211 => "00100111",1212 => "00001000",1213 => "11111011",1214 => "01011011",1215 => "10100000",1216 => "11101111",1217 => "00101110",1218 => "00001010",1219 => "01100110",1220 => "11101000",1221 => "11001111",1222 => "01010011",1223 => "00010000",1224 => "10011101",1225 => "01100001",1226 => "10100110",1227 => "00010100",1228 => "11000111",1229 => "10000010",1230 => "01100001",1231 => "00100011",1232 => "00011110",1233 => "00001010",1234 => "01001001",1235 => "01110110",1236 => "10100011",1237 => "11111100",1238 => "11001010",1239 => "00010110",1240 => "11110100",1241 => "11111011",1242 => "00011001",1243 => "10111111",1244 => "11001100",1245 => "10110010",1246 => "01000111",1247 => "10001101",1248 => "01110011",1249 => "00010101",1250 => "00000110",1251 => "10111100",1252 => "11100010",1253 => "00011001",1254 => "01001100",1255 => "01110101",1256 => "01111000",1257 => "11111010",1258 => "01010101",1259 => "01101001",1260 => "00001101",1261 => "01111111",1262 => "11010111",1263 => "00101000",1264 => "11111000",1265 => "10010011",1266 => "00100111",1267 => "01100011",1268 => "10111010",1269 => "00110101",1270 => "00110110",1271 => "00001100",1272 => "01100110",1273 => "11101111",1274 => "01111000",1275 => "11000111",1276 => "10100111",1277 => "01011111",1278 => "01000000",1279 => "11000100",1280 => "10100110",1281 => "00011011",1282 => "11010101",1283 => "00001010",1284 => "10011111",1285 => "11110100",1286 => "11010111",1287 => "10001011",1288 => "11000000",1289 => "11011010",1290 => "00111110",1291 => "11111001",1292 => "10100111",1293 => "00100011",1294 => "00001001",1295 => "11010010",1296 => "01100101",1297 => "01101000",1298 => "01010111",1299 => "10011001",1300 => "11110001",1301 => "01000101",1302 => "00100110",1303 => "10000001",1304 => "10110101",1305 => "00000110",1306 => "00110011",1307 => "00110000",1308 => "01110110",1309 => "10000000",1310 => "10111011",1311 => "01001000",1312 => "11001101",1313 => "10110111",1314 => "10101010",1315 => "00111101",1316 => "01011011",1317 => "01010101",1318 => "01100100",1319 => "10100001",1320 => "01100111",1321 => "01101111",1322 => "10100111",1323 => "01001100",1324 => "01110101",1325 => "10000111",1326 => "01000111",1327 => "11100100",1328 => "00000001",1329 => "11100101",1330 => "00000110",1331 => "10011110",1332 => "01010010",1333 => "01111111",1334 => "00101100",1335 => "10011110",1336 => "01110110",1337 => "11011110",1338 => "00010011",1339 => "11011011",1340 => "10001100",1341 => "00110011",1342 => "00000010",1343 => "01010110",1344 => "00101010",1345 => "11000010",1346 => "01001111",1347 => "00111011",1348 => "01011001",1349 => "10111000",1350 => "00010001",1351 => "00010110",1352 => "11010001",1353 => "11101001",1354 => "01011001",1355 => "01110000",1356 => "01010111",1357 => "11111110",1358 => "00011010",1359 => "01011001",1360 => "10010100",1361 => "01111000",1362 => "11000100",1363 => "11010011",1364 => "11011011",1365 => "11001101",1366 => "00101000",1367 => "10111101",1368 => "11010010",1369 => "00111001",1370 => "11110000",1371 => "10101111",1372 => "11010001",1373 => "00100010",1374 => "01111011",1375 => "00101111",1376 => "11000100",1377 => "01100110",1378 => "00111111",1379 => "10110100",1380 => "10100001",1381 => "01010011",1382 => "11111000",1383 => "00000011",1384 => "10100100",1385 => "10010010",1386 => "11000011",1387 => "11000001",1388 => "00110101",1389 => "00010110",1390 => "01011011",1391 => "11111000",1392 => "00010111",1393 => "01001100",1394 => "00111011",1395 => "01110000",1396 => "11010111",1397 => "10100000",1398 => "01000011",1399 => "00110000",1400 => "01010010",1401 => "10100010",1402 => "01001101",1403 => "00100101",1404 => "10011010",1405 => "11111011",1406 => "10100000",1407 => "10000000",1408 => "01000111",1409 => "11110111",1410 => "11111000",1411 => "01001000",1412 => "10101010",1413 => "11100111",1414 => "10010100",1415 => "11111001",1416 => "01110100",1417 => "00001010",1418 => "01001010",1419 => "01100000",1420 => "00110010",1421 => "00101011",1422 => "00011000",1423 => "00011101",1424 => "10001101",1425 => "01010100",1426 => "01001010",1427 => "10110010",1428 => "00110100",1429 => "00111010",1430 => "11100100",1431 => "00000101",1432 => "11101010",1433 => "11100010",1434 => "01011011",1435 => "11111000",1436 => "00110111",1437 => "00011110",1438 => "01111000",1439 => "01010111",1440 => "11100011",1441 => "01001111",1442 => "11001110",1443 => "00111101",1444 => "10011100",1445 => "00101011",1446 => "00000111",1447 => "01000110",1448 => "01110000",1449 => "00101101",1450 => "11101111",1451 => "11000100",1452 => "01100110",1453 => "01101111",1454 => "01011000",1455 => "01010001",1456 => "00000100",1457 => "10010101",1458 => "11000110",1459 => "11111011",1460 => "01000111",1461 => "00011001",1462 => "00110001",1463 => "01010000",1464 => "00111010",1465 => "11111011",1466 => "11001101",1467 => "01111000",1468 => "00000100",1469 => "10110010",1470 => "00100101",1471 => "00111010",1472 => "01100111",1473 => "10111001",1474 => "10101110",1475 => "11000001",1476 => "00110110",1477 => "11100000",1478 => "01000110",1479 => "11101010",1480 => "11001011",1481 => "10110111",1482 => "10110010",1483 => "11110101",1484 => "00110101",1485 => "00011100",1486 => "01100010",1487 => "10111101",1488 => "00101100",1489 => "10111110",1490 => "11111101",1491 => "00011101",1492 => "11010010",1493 => "00001010",1494 => "10010000",1495 => "00110101",1496 => "10010100",1497 => "11110111",1498 => "00111010",1499 => "11010000",1500 => "11000001",1501 => "01101101",1502 => "11100110",1503 => "00111111",1504 => "11000010",1505 => "11111001",1506 => "10101000",1507 => "00110101",1508 => "01101000",1509 => "00110110",1510 => "01101000",1511 => "01100111",1512 => "10100100",1513 => "01111111",1514 => "00001111",1515 => "10110000",1516 => "10010100",1517 => "01010010",1518 => "11010101",1519 => "10110010",1520 => "10111010",1521 => "00011000",1522 => "01110100",1523 => "00110000",1524 => "00110011",1525 => "01000001",1526 => "11010000",1527 => "11100010",1528 => "01001111",1529 => "11010001",1530 => "10000011",1531 => "11010010",1532 => "10000100",1533 => "00111010",1534 => "01110001",1535 => "10100011",1536 => "01001010",1537 => "00011101",1538 => "11111000",1539 => "11001110",1540 => "00101000",1541 => "01010011",1542 => "11000110",1543 => "01000010",1544 => "11000011",1545 => "10001010",1546 => "00000011",1547 => "00100110",1548 => "11101100",1549 => "01100100",1550 => "00110010",1551 => "11011011",1552 => "01001000",1553 => "11010110",1554 => "10101101",1555 => "00000101",1556 => "01110000",1557 => "00000011",1558 => "00011000",1559 => "11100100",1560 => "10101001",1561 => "10110000",1562 => "01000000",1563 => "11101101",1564 => "11001101",1565 => "10101100",1566 => "00111100",1567 => "11101001",1568 => "00100101",1569 => "01100110",1570 => "11111100",1571 => "00000101",1572 => "01111110",1573 => "00001111",1574 => "01101110",1575 => "11010010",1576 => "10001100",1577 => "00110101",1578 => "11101000",1579 => "10011110",1580 => "00010000",1581 => "00010110",1582 => "10000001",1583 => "01111010",1584 => "01010100",1585 => "11111110",1586 => "10001000",1587 => "00011000",1588 => "00001100",1589 => "11001111",1590 => "01111011",1591 => "10110010",1592 => "11111010",1593 => "00100101",1594 => "11010010",1595 => "00000000",1596 => "11001101",1597 => "11110110",1598 => "01000000",1599 => "11010010",1600 => "00011011",1601 => "01101000",1602 => "00000110",1603 => "11000011",1604 => "00101010",1605 => "11110000",1606 => "10001110",1607 => "10101010",1608 => "11010001",1609 => "01101100",1610 => "11001111",1611 => "01011110",1612 => "10011111",1613 => "10100111",1614 => "10010001",1615 => "10110000",1616 => "00010001",1617 => "10000111",1618 => "11000100",1619 => "01110000",1620 => "00101110",1621 => "11000011",1622 => "00101000",1623 => "01011011",1624 => "10011010",1625 => "10110001",1626 => "01100010",1627 => "01001011",1628 => "00111001",1629 => "10011010",1630 => "01000100",1631 => "11101100",1632 => "10001101",1633 => "01001010",1634 => "11011101",1635 => "00111111",1636 => "11011011",1637 => "00001000",1638 => "01010000",1639 => "01110100",1640 => "10101000",1641 => "01111100",1642 => "01011000",1643 => "01010110",1644 => "11100001",1645 => "11110110",1646 => "11100011",1647 => "01110100",1648 => "11001111",1649 => "11111000",1650 => "01000011",1651 => "10001100",1652 => "01001010",1653 => "01100001",1654 => "11111001",1655 => "01101010",1656 => "01000110",1657 => "00010010",1658 => "01100010",1659 => "10100001",1660 => "10111101",1661 => "10011010",1662 => "11000111",1663 => "00001011",1664 => "11010111",1665 => "00100010",1666 => "01101101",1667 => "11000101",1668 => "11000111",1669 => "00010100",1670 => "00000000",1671 => "00001110",1672 => "01000010",1673 => "00000100",1674 => "01011101",1675 => "01000000",1676 => "00110000",1677 => "01010011",1678 => "10110001",1679 => "01111010",1680 => "10101100",1681 => "00111111",1682 => "10110010",1683 => "10101000",1684 => "00010100",1685 => "11100101",1686 => "00111110",1687 => "11110111",1688 => "11101110",1689 => "01011010",1690 => "00111010",1691 => "11110000",1692 => "11000011",1693 => "10010000",1694 => "10110110",1695 => "10001101",1696 => "11110111",1697 => "00110010",1698 => "11110111",1699 => "01101011",1700 => "00010101",1701 => "10101100",1702 => "01011001",1703 => "10111101",1704 => "01010010",1705 => "11100100",1706 => "01111100",1707 => "00101101",1708 => "01011010",1709 => "11111000",1710 => "01010011",1711 => "01110111",1712 => "11001111",1713 => "00011010",1714 => "00010001",1715 => "00000110",1716 => "11110011",1717 => "01111000",1718 => "10100100",1719 => "10010010",1720 => "10000101",1721 => "00110011",1722 => "00101010",1723 => "00000100",1724 => "10101011",1725 => "00010011",1726 => "10000111",1727 => "01001111",1728 => "11110010",1729 => "11010110",1730 => "00100111",1731 => "00101101",1732 => "00100000",1733 => "11001001",1734 => "10100101",1735 => "11100010",1736 => "10100100",1737 => "10001000",1738 => "11111110",1739 => "10110010",1740 => "01101110",1741 => "10111101",1742 => "11001010",1743 => "01100111",1744 => "01101101",1745 => "10000001",1746 => "01100101",1747 => "10000000",1748 => "01011101",1749 => "10101000",1750 => "10011010",1751 => "00111001",1752 => "01001011",1753 => "10110000",1754 => "10011100",1755 => "10111001",1756 => "01101111",1757 => "11101101",1758 => "11111111",1759 => "01000111",1760 => "00011111",1761 => "10000011",1762 => "01100010",1763 => "01100000",1764 => "10000000",1765 => "00100101",1766 => "11001101",1767 => "00001111",1768 => "11001001",1769 => "10000101",1770 => "11000001",1771 => "00011100",1772 => "11110011",1773 => "01011101",1774 => "11010100",1775 => "10101111",1776 => "01100011",1777 => "11110100",1778 => "01100111",1779 => "00011101",1780 => "10101000",1781 => "01011000",1782 => "11110100",1783 => "11001010",1784 => "01001100",1785 => "11110111",1786 => "11111000",1787 => "10100000",1788 => "00010001",1789 => "01001110",1790 => "11001000",1791 => "11111100",1792 => "01011110",1793 => "01000011",1794 => "10010100",1795 => "01110100",1796 => "10101100",1797 => "00011100",1798 => "00111111",1799 => "10110000",1800 => "01011111",1801 => "00101000",1802 => "10001101",1803 => "10110001",1804 => "10010111",1805 => "00101000",1806 => "01111011",1807 => "11010111",1808 => "11010100",1809 => "11111110",1810 => "00010100",1811 => "00101110",1812 => "11101101",1813 => "11111110",1814 => "11110001",1815 => "11101110",1816 => "01110011",1817 => "10111111",1818 => "10101111",1819 => "10001000",1820 => "01011110",1821 => "01011011",1822 => "01100011",1823 => "11001001",1824 => "01001010",1825 => "01111010",1826 => "01011000",1827 => "00010100",1828 => "11001001",1829 => "11000001",1830 => "01101101",1831 => "00101000",1832 => "00101101",1833 => "10100010",1834 => "11001000",1835 => "11101101",1836 => "01100100",1837 => "11100001",1838 => "11001011",1839 => "01100100",1840 => "11111101",1841 => "00000100",1842 => "10110001",1843 => "00011100",1844 => "11011110",1845 => "00000011",1846 => "01110010",1847 => "01000101",1848 => "01010111",1849 => "11100010",1850 => "01000011",1851 => "11010101",1852 => "00100000",1853 => "01011010",1854 => "00000101",1855 => "11110110",1856 => "11110110",1857 => "11100100",1858 => "10001011",1859 => "01011000",1860 => "00001110",1861 => "11100101",1862 => "11111011",1863 => "01011110",1864 => "11010110",1865 => "11000101",1866 => "01111101",1867 => "01110111",1868 => "00010111",1869 => "00010110",1870 => "01001100",1871 => "10001000",1872 => "01001001",1873 => "11100110",1874 => "00101011",1875 => "10110001",1876 => "01101001",1877 => "10111011",1878 => "10011110",1879 => "10101011",1880 => "00100110",1881 => "11010110",1882 => "10011111",1883 => "10101110",1884 => "00000100",1885 => "00111011",1886 => "11010110",1887 => "00010100",1888 => "00011000",1889 => "11111001",1890 => "10100001",1891 => "10101010",1892 => "10110101",1893 => "00000111",1894 => "01101001",1895 => "11111100",1896 => "00111100",1897 => "11001011",1898 => "00010100",1899 => "10110101",1900 => "10101000",1901 => "01110101",1902 => "11101101",1903 => "00000111",1904 => "00110011",1905 => "01110100",1906 => "00011111",1907 => "10110101",1908 => "10111101",1909 => "00011101",1910 => "10011101",1911 => "01001000",1912 => "10101111",1913 => "11001011",1914 => "11101001",1915 => "01010111",1916 => "00111100",1917 => "00100111",1918 => "10001111",1919 => "01011000",1920 => "01100101",1921 => "10100101",1922 => "00110100",1923 => "11000110",1924 => "11011100",1925 => "10010100",1926 => "11100000",1927 => "00000011",1928 => "01100110",1929 => "01100101",1930 => "10001010",1931 => "10111101",1932 => "00011010",1933 => "11010010",1934 => "01011000",1935 => "00010010",1936 => "01111110",1937 => "01110110",1938 => "11111011",1939 => "10000011",1940 => "11011001",1941 => "01000101",1942 => "00001001",1943 => "11001100",1944 => "01001111",1945 => "11011101",1946 => "01100000",1947 => "10011010",1948 => "11000010",1949 => "01100011",1950 => "10000111",1951 => "11101101",1952 => "10011000",1953 => "11010101",1954 => "00001110",1955 => "11010010",1956 => "10001110",1957 => "01000101",1958 => "10110101",1959 => "10000001",1960 => "11001010",1961 => "00100011",1962 => "10101101",1963 => "11011001",1964 => "10111010",1965 => "10110010",1966 => "10100101",1967 => "10010111",1968 => "11010010",1969 => "01011101",1970 => "01100101",1971 => "01101110",1972 => "01100011",1973 => "00110010",1974 => "11101111",1975 => "10101001",1976 => "00100110",1977 => "01100100",1978 => "11111000",1979 => "10110010",1980 => "11110101",1981 => "11101000",1982 => "10100101",1983 => "00101000",1984 => "01011011",1985 => "11111000",1986 => "11000101",1987 => "10001000",1988 => "00110001",1989 => "11010111",1990 => "01001101",1991 => "01000011",1992 => "01101001",1993 => "10111100",1994 => "10011101",1995 => "00110101",1996 => "11101001",1997 => "00011010",1998 => "11101111",1999 => "11101101",2000 => "01000111",2001 => "10001011",2002 => "01110100",2003 => "00110001",2004 => "00000110",2005 => "10101010",2006 => "11111110",2007 => "01011110",2008 => "00100001",2009 => "00111101",2010 => "10010011",2011 => "10101001",2012 => "00111110",2013 => "01100000",2014 => "10010001",2015 => "11011010",2016 => "11110111",2017 => "10111101",2018 => "00001111",2019 => "00100011",2020 => "11111011",2021 => "00100111",2022 => "10001010",2023 => "10011101",2024 => "10010111",2025 => "01000000",2026 => "11110000",2027 => "11101000",2028 => "01011001",2029 => "00001010",2030 => "01001101",2031 => "00100011",2032 => "11001000",2033 => "11000010",2034 => "00000110",2035 => "10101010",2036 => "00100000",2037 => "10010000",2038 => "01011110",2039 => "11110100",2040 => "01101001",2041 => "00110111",2042 => "01101011",2043 => "00010101",2044 => "10001100",2045 => "00101100",2046 => "10010111",2047 => "11110001",2048 => "00110001",2049 => "01110110",2050 => "10100110",2051 => "10010100",2052 => "00101010",2053 => "00111110",2054 => "11100010",2055 => "01000011",2056 => "00110011",2057 => "10001010",2058 => "10000000",2059 => "00000110",2060 => "01110101",2061 => "01001000",2062 => "01001011",2063 => "00001001",2064 => "01011000",2065 => "11100111",2066 => "00001110",2067 => "10000011",2068 => "11010001",2069 => "10101100",2070 => "01010110",2071 => "11111000",2072 => "11010000",2073 => "01100111",2074 => "11110111",2075 => "00111001",2076 => "10101110",2077 => "00111000",2078 => "11110001",2079 => "01010000",2080 => "11011100",2081 => "11001000",2082 => "01001001",2083 => "11111110",2084 => "10000001",2085 => "10001101",2086 => "01111100",2087 => "01001010",2088 => "01100100",2089 => "10111011",2090 => "11111010",2091 => "01111110",2092 => "11101010",2093 => "10000110",2094 => "00010101",2095 => "11110111",2096 => "00110100",2097 => "00111011",2098 => "00000010",2099 => "10100101",2100 => "00010101",2101 => "01100101",2102 => "11011111",2103 => "00111111",2104 => "11000111",2105 => "11101111",2106 => "11001010",2107 => "10000100",2108 => "11000001",2109 => "11110001",2110 => "11101000",2111 => "10110001",2112 => "01000010",2113 => "00110001",2114 => "01001000",2115 => "01110011",2116 => "00110010",2117 => "01010111",2118 => "00011001",2119 => "10110000",2120 => "10111001",2121 => "11001001",2122 => "01111100",2123 => "11110100",2124 => "00111011",2125 => "01000111",2126 => "01000011",2127 => "00011011",2128 => "00011111",2129 => "10110010",2130 => "01110010",2131 => "11100010",2132 => "00111110",2133 => "11100101",2134 => "00011110",2135 => "01111000",2136 => "00100010",2137 => "00001000",2138 => "11101101",2139 => "10001001",2140 => "01011101",2141 => "00010100",2142 => "11001110",2143 => "11001110",2144 => "00100001",2145 => "01011011",2146 => "00000010",2147 => "01111001",2148 => "10001111",2149 => "01001100",2150 => "11111011",2151 => "10101100",2152 => "10011000",2153 => "11010011",2154 => "01100101",2155 => "10001101",2156 => "00111011",2157 => "11111100",2158 => "00011000",2159 => "01011110",2160 => "11001111",2161 => "00011011",2162 => "11011111",2163 => "11010101",2164 => "11111111",2165 => "01001101",2166 => "01110010",2167 => "11110011",2168 => "01011101",2169 => "00011110",2170 => "11111111",2171 => "11110000",2172 => "10111110",2173 => "10110111",2174 => "11100001",2175 => "10100010",2176 => "10000100",2177 => "11000100",2178 => "10001110",2179 => "01000101",2180 => "01001110",2181 => "00100010",2182 => "00001000",2183 => "01011101",2184 => "01001110",2185 => "10000110",2186 => "10110111",2187 => "01110100",2188 => "11001000",2189 => "10101110",2190 => "10001110",2191 => "11010001",2192 => "11110100",2193 => "10010000",2194 => "01100101",2195 => "01110000",2196 => "01000111",2197 => "01101111",2198 => "10101101",2199 => "00110011",2200 => "01011001",2201 => "01100101",2202 => "10001110",2203 => "11100100",2204 => "00111000",2205 => "10011100",2206 => "11101010",2207 => "11001111",2208 => "10110010",2209 => "11010101",2210 => "11111110",2211 => "10000000",2212 => "10001000",2213 => "01010000",2214 => "11100100",2215 => "10101110",2216 => "00110010",2217 => "11011001",2218 => "11011101",2219 => "10110110",2220 => "01010110",2221 => "11011100",2222 => "11100011",2223 => "10001000",2224 => "01011011",2225 => "10001100",2226 => "10111110",2227 => "00000000",2228 => "10111100",2229 => "00001101",2230 => "00101111",2231 => "01010111",2232 => "01101100",2233 => "11101100",2234 => "11011100",2235 => "10100001",2236 => "00100011",2237 => "10011100",2238 => "10110100",2239 => "10011100",2240 => "10011010",2241 => "11101010",2242 => "11101101",2243 => "01100101",2244 => "11010000",2245 => "11011111",2246 => "01101000",2247 => "01010001",2248 => "01000010",2249 => "01111111",2250 => "11110001",2251 => "00001010",2252 => "11100100",2253 => "10101001",2254 => "00111000",2255 => "11100100",2256 => "00000010",2257 => "01011101",2258 => "11010011",2259 => "01011101",2260 => "10001011",2261 => "00110000",2262 => "00100100",2263 => "00010111",2264 => "00010011",2265 => "01110011",2266 => "11111011",2267 => "01010011",2268 => "00001011",2269 => "00001100",2270 => "11101010",2271 => "11000111",2272 => "11100111",2273 => "11000110",2274 => "01000100",2275 => "10010001",2276 => "10110110",2277 => "00111101",2278 => "01100100",2279 => "10110011",2280 => "11111010",2281 => "10110010",2282 => "01011001",2283 => "10101000",2284 => "01011111",2285 => "01100011",2286 => "01110110",2287 => "10100110",2288 => "01000100",2289 => "00101000",2290 => "11101010",2291 => "11000111",2292 => "00100111",2293 => "11110011",2294 => "10101011",2295 => "11001100",2296 => "11110001",2297 => "01001000",2298 => "01111001",2299 => "10101011",2300 => "01100110",2301 => "10101011",2302 => "00011101",2303 => "10010010",2304 => "11111010",2305 => "11101011",2306 => "10010001",2307 => "10010100",2308 => "01111111",2309 => "11000101",2310 => "11000101",2311 => "10001101",2312 => "10110101",2313 => "00000011",2314 => "10001100",2315 => "00110011",2316 => "00011100",2317 => "11000111",2318 => "11100110",2319 => "00011000",2320 => "00101011",2321 => "11001000",2322 => "01101101",2323 => "01010010",2324 => "11001100",2325 => "01000100",2326 => "01000000",2327 => "01011010",2328 => "10111000",2329 => "00000100",2330 => "00100111",2331 => "11011001",2332 => "01011011",2333 => "00011011",2334 => "01101000",2335 => "10001111",2336 => "01101001",2337 => "11011100",2338 => "00101110",2339 => "01001111",2340 => "10000011",2341 => "11010101",2342 => "00101000",2343 => "01111010",2344 => "11001010",2345 => "10111011",2346 => "01111000",2347 => "11010111",2348 => "10001111",2349 => "00101010",2350 => "00011110",2351 => "00101000",2352 => "01100101",2353 => "10111101",2354 => "11001111",2355 => "10001001",2356 => "10111101",2357 => "10010100",2358 => "00110010",2359 => "00101011",2360 => "11011000",2361 => "11100011",2362 => "10110100",2363 => "11110101",2364 => "11100101",2365 => "01100100",2366 => "01000000",2367 => "00100001",2368 => "10001010",2369 => "01001110",2370 => "10001001",2371 => "10000011",2372 => "10011111",2373 => "00000010",2374 => "11011100",2375 => "00100100",2376 => "11000000",2377 => "00101101",2378 => "10100100",2379 => "01000100",2380 => "01000101",2381 => "11111101",2382 => "01100010",2383 => "11110110",2384 => "10011011",2385 => "11111011",2386 => "01101101",2387 => "01101110",2388 => "11100011",2389 => "10111101",2390 => "10000001",2391 => "10001101",2392 => "00111111",2393 => "11001110",2394 => "01011000",2395 => "11010001",2396 => "01111011",2397 => "10101011",2398 => "01001001",2399 => "10110100",2400 => "11110000",2401 => "10010101",2402 => "01100000",2403 => "11111011",2404 => "11000101",2405 => "01011111",2406 => "00100001",2407 => "01001101",2408 => "10110100",2409 => "01110101",2410 => "11010111",2411 => "00100011",2412 => "00101111",2413 => "01001100",2414 => "00001000",2415 => "10110001",2416 => "11110110",2417 => "01001111",2418 => "00001111",2419 => "10001000",2420 => "11101000",2421 => "10111001",2422 => "10010110",2423 => "10010110",2424 => "11000101",2425 => "00000111",2426 => "11000111",2427 => "11011101",2428 => "00001111",2429 => "01110010",2430 => "11000010",2431 => "01110011",2432 => "00100110",2433 => "11001110",2434 => "10001101",2435 => "00001010",2436 => "01101100",2437 => "10011011",2438 => "10111100",2439 => "00010011",2440 => "11110000",2441 => "00100011",2442 => "00011110",2443 => "01111100",2444 => "00101110",2445 => "01011011",2446 => "00010000",2447 => "10001111",2448 => "10000110",2449 => "11011001",2450 => "11011111",2451 => "01101011",2452 => "11111000",2453 => "00111110",2454 => "00100101",2455 => "11000111",2456 => "11001110",2457 => "10111110",2458 => "10001100",2459 => "01111100",2460 => "11010000",2461 => "10000110",2462 => "11010010",2463 => "01101010",2464 => "11111011",2465 => "10110001",2466 => "00000101",2467 => "11110001",2468 => "01001110",2469 => "00011111",2470 => "00001000",2471 => "10110101",2472 => "01000111",2473 => "10010011",2474 => "10010100",2475 => "11111000",2476 => "00010010",2477 => "01000111",2478 => "00010011",2479 => "00000100",2480 => "10101000",2481 => "00011001",2482 => "11100110",2483 => "01100000",2484 => "01100010",2485 => "01111001",2486 => "10111001",2487 => "01000111",2488 => "01000011",2489 => "11011011",2490 => "10100101",2491 => "10001100",2492 => "01111010",2493 => "00100001",2494 => "01110111",2495 => "10111001",2496 => "11111110",2497 => "01100100",2498 => "00011110",2499 => "11000011",2500 => "11100010",2501 => "01011110",2502 => "11101111",2503 => "01010000",2504 => "00101101",2505 => "10010001",2506 => "10010101",2507 => "11001011",2508 => "00001101",2509 => "01101110",2510 => "10011001",2511 => "11101100",2512 => "11101000",2513 => "11110111",2514 => "11000011",2515 => "10000011",2516 => "10101111",2517 => "00011110",2518 => "01100011",2519 => "10100000",2520 => "11100011",2521 => "00000001",2522 => "11111011",2523 => "00100011",2524 => "01010110",2525 => "01111010",2526 => "00011001",2527 => "01111000",2528 => "01111010",2529 => "10011010",2530 => "00011101",2531 => "10111011",2532 => "11001000",2533 => "01111101",2534 => "00001100",2535 => "10010001",2536 => "01100100",2537 => "01011010",2538 => "00101110",2539 => "10111100",2540 => "11110100",2541 => "10100100",2542 => "00010010",2543 => "01010110",2544 => "00010111",2545 => "10001100",2546 => "11011101",2547 => "11001110",2548 => "00000001",2549 => "11110010",2550 => "01000100",2551 => "11101011",2552 => "01110100",2553 => "11110101",2554 => "10011000",2555 => "10100000",2556 => "11111111",2557 => "00111010",2558 => "10100111",2559 => "01100000",2560 => "11101000",2561 => "11111100",2562 => "10110000",2563 => "10111010",2564 => "11110010",2565 => "01000011",2566 => "10001000",2567 => "10100111",2568 => "00101111",2569 => "10010001",2570 => "00010110",2571 => "00110001",2572 => "00110011",2573 => "10100000",2574 => "00100100",2575 => "10010111",2576 => "00000001",2577 => "01101100",2578 => "01001001",2579 => "11100111",2580 => "11100010",2581 => "11000011",2582 => "01011000",2583 => "01110100",2584 => "00001010",2585 => "00010101",2586 => "11000101",2587 => "11011100",2588 => "11011111",2589 => "11111000",2590 => "00100010",2591 => "11111111",2592 => "00101000",2593 => "01010001",2594 => "10000111",2595 => "01101001",2596 => "01010010",2597 => "10010010",2598 => "01111001",2599 => "11101001",2600 => "11010100",2601 => "01011110",2602 => "01101111",2603 => "11100001",2604 => "00100100",2605 => "11011101",2606 => "00001011",2607 => "10100100",2608 => "01111111",2609 => "00101000",2610 => "00111101",2611 => "10010110",2612 => "10100110",2613 => "11001110",2614 => "11110011",2615 => "00000100",2616 => "01111000",2617 => "11001010",2618 => "01100100",2619 => "10000001",2620 => "00110001",2621 => "10001111",2622 => "10100110",2623 => "01010000",2624 => "11111001",2625 => "11010000",2626 => "10000100",2627 => "10000011",2628 => "00111110",2629 => "10100001",2630 => "10011111",2631 => "01110110",2632 => "11110010",2633 => "11110111",2634 => "01010101",2635 => "00101101",2636 => "10001100",2637 => "11010001",2638 => "00110001",2639 => "01010111",2640 => "11111000",2641 => "10100001",2642 => "01011011",2643 => "10111001",2644 => "00010000",2645 => "11010001",2646 => "11100110",2647 => "10100010",2648 => "11000111",2649 => "10000100",2650 => "11111001",2651 => "11111101",2652 => "11010011",2653 => "11011000",2654 => "10011010",2655 => "00010011",2656 => "10100000",2657 => "11000001",2658 => "10100101",2659 => "00110010",2660 => "11001001",2661 => "11000100",2662 => "00111011",2663 => "01111010",2664 => "11001011",2665 => "10000011",2666 => "10111010",2667 => "00000111",2668 => "00010000",2669 => "11000110",2670 => "11111010",2671 => "11111000",2672 => "00011110",2673 => "01101000",2674 => "00000110",2675 => "01110011",2676 => "10100000",2677 => "00110010",2678 => "01010010",2679 => "10110100",2680 => "01100101",2681 => "11010011",2682 => "01101100",2683 => "10101000",2684 => "11110010",2685 => "11111111",2686 => "00100001",2687 => "11101100",2688 => "10011000",2689 => "10101010",2690 => "11101001",2691 => "11111011",2692 => "00101100",2693 => "11001110",2694 => "11000100",2695 => "10101100",2696 => "00001011",2697 => "01110010",2698 => "11100100",2699 => "00100000",2700 => "01111001",2701 => "01000110",2702 => "00010101",2703 => "01110100",2704 => "00010011",2705 => "01101101",2706 => "11101000",2707 => "10110000",2708 => "01001001",2709 => "00001110",2710 => "11000001",2711 => "00011110",2712 => "10001001",2713 => "11001011",2714 => "11101010",2715 => "01001101",2716 => "01111011",2717 => "01100110",2718 => "01111100",2719 => "10010111",2720 => "10100001",2721 => "01101110",2722 => "11110011",2723 => "10111001",2724 => "00111001",2725 => "10010100",2726 => "01110110",2727 => "11100010",2728 => "01100101",2729 => "11010101",2730 => "11001000",2731 => "01100100",2732 => "01110111",2733 => "00001111",2734 => "11011101",2735 => "11101010",2736 => "01011010",2737 => "11001111",2738 => "01101010",2739 => "00000100",2740 => "00001101",2741 => "00110100",2742 => "01110100",2743 => "10101000",2744 => "00110001",2745 => "01100110",2746 => "01111000",2747 => "10100101",2748 => "11101010",2749 => "11011110",2750 => "01101001",2751 => "00010101",2752 => "01010000",2753 => "11101101",2754 => "10101011",2755 => "10101010",2756 => "10110110",2757 => "01000010",2758 => "10101011",2759 => "00000101",2760 => "00000001",2761 => "10101001",2762 => "01110100",2763 => "00110010",2764 => "01011000",2765 => "00000101",2766 => "10000110",2767 => "10001100",2768 => "10111111",2769 => "00111000",2770 => "11101111",2771 => "10101000",2772 => "10101111",2773 => "10011001",2774 => "01111101",2775 => "10010010",2776 => "01111100",2777 => "01100100",2778 => "10101111",2779 => "01001011",2780 => "01110010",2781 => "11001110",2782 => "00100100",2783 => "11001101",2784 => "10101001",2785 => "11110010",2786 => "00110000",2787 => "01111100",2788 => "10100110",2789 => "01001111",2790 => "11000100",2791 => "11110001",2792 => "11101101",2793 => "11000000",2794 => "11110110",2795 => "11100111",2796 => "10101110",2797 => "11111010",2798 => "10101010",2799 => "11000010",2800 => "00001110",2801 => "00100001",2802 => "10111011",2803 => "00100110",2804 => "01001101",2805 => "10101101",2806 => "00001000",2807 => "11111001",2808 => "01000110",2809 => "00100001",2810 => "01111001",2811 => "01010111",2812 => "01100100",2813 => "01100101",2814 => "00011110",2815 => "00110000",2816 => "01001111",2817 => "00101110",2818 => "11001101",2819 => "11001001",2820 => "01100101",2821 => "00100001",2822 => "10101101",2823 => "11010001",2824 => "00101011",2825 => "01001011",2826 => "01111110",2827 => "11010000",2828 => "01010001",2829 => "01110110",2830 => "01001100",2831 => "01111000",2832 => "01001000",2833 => "10000010",2834 => "01100000",2835 => "11111100",2836 => "10011110",2837 => "11011100",2838 => "10101111",2839 => "10000010",2840 => "11111101",2841 => "10010000",2842 => "10110100",2843 => "00010110",2844 => "01110101",2845 => "01011110",2846 => "10100000",2847 => "11001110",2848 => "00010011",2849 => "01101000",2850 => "10100111",2851 => "11000100",2852 => "00101001",2853 => "11111001",2854 => "11010100",2855 => "01001011",2856 => "11100111",2857 => "10001101",2858 => "00011010",2859 => "00001101",2860 => "11000111",2861 => "10101100",2862 => "01010011",2863 => "00101010",2864 => "11000010",2865 => "11011100",2866 => "01000011",2867 => "11110100",2868 => "11101011",2869 => "11111111",2870 => "11001001",2871 => "11101111",2872 => "11010010",2873 => "11100111",2874 => "10111101",2875 => "10000010",2876 => "10111011",2877 => "10001111",2878 => "10001111",2879 => "00100010",2880 => "00101010",2881 => "00001001",2882 => "00010001",2883 => "10001110",2884 => "01010000",2885 => "01000110",2886 => "11011010",2887 => "00101111",2888 => "10110011",2889 => "11000000",2890 => "00110100",2891 => "01101100",2892 => "11001010",2893 => "11100110",2894 => "10001011",2895 => "01001101",2896 => "11111100",2897 => "01001011",2898 => "01111100",2899 => "11010101",2900 => "01111000",2901 => "01110010",2902 => "01100010",2903 => "11111111",2904 => "10010011",2905 => "01100100",2906 => "11111011",2907 => "11111110",2908 => "01001101",2909 => "10011101",2910 => "11001110",2911 => "00110001",2912 => "11101011",2913 => "01111001",2914 => "00111101",2915 => "00011010",2916 => "00011010",2917 => "00110000",2918 => "00001101",2919 => "01010011",2920 => "00001011",2921 => "01111111",2922 => "10100111",2923 => "01111000",2924 => "10111001",2925 => "11100001",2926 => "01011010",2927 => "01101011",2928 => "11100100",2929 => "11100101",2930 => "11111001",2931 => "00110000",2932 => "00110000",2933 => "11110011",2934 => "11100101",2935 => "00011100",2936 => "01111000",2937 => "11000100",2938 => "00110100",2939 => "01010001",2940 => "00111000",2941 => "10111110",2942 => "00000101",2943 => "11101001",2944 => "01011101",2945 => "01110001",2946 => "11110010",2947 => "00101110",2948 => "10011101",2949 => "00100011",2950 => "10001000",2951 => "10000001",2952 => "10001000",2953 => "01001111",2954 => "10100110",2955 => "01000101",2956 => "01101010",2957 => "10010101",2958 => "10011111",2959 => "01011111",2960 => "01101001",2961 => "00101110",2962 => "10100010",2963 => "10000111",2964 => "10100111",2965 => "01111100",2966 => "01101001",2967 => "01011101",2968 => "10110000",2969 => "01111010",2970 => "01011100",2971 => "10101101",2972 => "00010010",2973 => "00110111",2974 => "00101000",2975 => "11110111",2976 => "00001011",2977 => "10010101",2978 => "01010110",2979 => "01001110",2980 => "00111000",2981 => "01111111",2982 => "00000010",2983 => "01000010",2984 => "01110010",2985 => "10101011",2986 => "11010111",2987 => "01001111",2988 => "11010110",2989 => "00110110",2990 => "01000001",2991 => "00000010",2992 => "01000110",2993 => "10001010",2994 => "11001001",2995 => "10100011",2996 => "11001110",2997 => "11110110",2998 => "11100010",2999 => "00010101",3000 => "01011100",3001 => "10010110",3002 => "01100010",3003 => "11100110",3004 => "11100010",3005 => "10000010",3006 => "00001100",3007 => "10101111",3008 => "10111101",3009 => "00010100",3010 => "00011100",3011 => "01000110",3012 => "00011101",3013 => "01100101",3014 => "01011000",3015 => "01100010",3016 => "00100001",3017 => "00100001",3018 => "11110110",3019 => "11001010",3020 => "11011100",3021 => "11100010",3022 => "10011001",3023 => "01100001",3024 => "01000101",3025 => "10001101",3026 => "00001000",3027 => "00001101",3028 => "00001010",3029 => "10100100",3030 => "10010001",3031 => "01000011",3032 => "01011000",3033 => "10100111",3034 => "11101110",3035 => "00111100",3036 => "00100110",3037 => "01100000",3038 => "01000000",3039 => "00010001",3040 => "10111100",3041 => "11110011",3042 => "01100010",3043 => "00001011",3044 => "01011101",3045 => "11010000",3046 => "01100001",3047 => "00010100",3048 => "00111101",3049 => "10000011",3050 => "11110100",3051 => "11000001",3052 => "00101101",3053 => "11010010",3054 => "11101111",3055 => "10000001",3056 => "01001011",3057 => "01111101",3058 => "10001101",3059 => "11101110",3060 => "00001011",3061 => "00100001",3062 => "01010000",3063 => "10110010",3064 => "01010000",3065 => "11011111",3066 => "10010101",3067 => "10010010",3068 => "11101110",3069 => "01100000",3070 => "10100011",3071 => "10101100",3072 => "01011001",3073 => "01110011",3074 => "00100011",3075 => "10010001",3076 => "00010001",3077 => "00100111",3078 => "10000110",3079 => "00100100",3080 => "10101000",3081 => "11000000",3082 => "00011100",3083 => "11011111",3084 => "00001001",3085 => "00110000",3086 => "10010011",3087 => "11101000",3088 => "00100010",3089 => "00111110",3090 => "00100110",3091 => "10001110",3092 => "00000110",3093 => "10000110",3094 => "10100101",3095 => "00011000",3096 => "11001111",3097 => "10100000",3098 => "01110011",3099 => "00000000",3100 => "10101100",3101 => "01100010",3102 => "01010101",3103 => "00011100",3104 => "11001001",3105 => "11011101",3106 => "00101010",3107 => "11101010",3108 => "11111101",3109 => "11100010",3110 => "00100110",3111 => "00011000",3112 => "01111101",3113 => "00111010",3114 => "01010001",3115 => "01111001",3116 => "00100001",3117 => "00100011",3118 => "00101010",3119 => "00101001",3120 => "11001101",3121 => "00100000",3122 => "10010001",3123 => "11111010",3124 => "10011011",3125 => "10001000",3126 => "01110010",3127 => "00110111",3128 => "01101101",3129 => "00110111",3130 => "11001010",3131 => "11000011",3132 => "11110000",3133 => "10000100",3134 => "11001001",3135 => "01001011",3136 => "01000100",3137 => "11001111",3138 => "11101101",3139 => "00110000",3140 => "11010111",3141 => "01110000",3142 => "11001101",3143 => "11010010",3144 => "11100110",3145 => "01001011",3146 => "00110010",3147 => "01000001",3148 => "00011101",3149 => "11100100",3150 => "10011011",3151 => "10100000",3152 => "10001001",3153 => "11010010",3154 => "10000101",3155 => "11011010",3156 => "00111101",3157 => "00101001",3158 => "01111100",3159 => "01110010",3160 => "10001001",3161 => "01100001",3162 => "01000100",3163 => "11110110",3164 => "01101100",3165 => "11111111",3166 => "01011101",3167 => "11111100",3168 => "00011101",3169 => "11101011",3170 => "01100100",3171 => "01110011",3172 => "11000101",3173 => "10011001",3174 => "01110111",3175 => "10011100",3176 => "11100110",3177 => "11110011",3178 => "01011100",3179 => "00100000",3180 => "00100101",3181 => "00111111",3182 => "01110100",3183 => "11100111",3184 => "00010011",3185 => "01100011",3186 => "11100101",3187 => "01011010",3188 => "01101111",3189 => "01001001",3190 => "10001000",3191 => "11010000",3192 => "11110001",3193 => "10111000",3194 => "11000001",3195 => "11111100",3196 => "11110001",3197 => "11011011",3198 => "01011100",3199 => "01010011",3200 => "10000110",3201 => "00000010",3202 => "01101101",3203 => "11000011",3204 => "11011110",3205 => "00100111",3206 => "00011100",3207 => "10001111",3208 => "11000001",3209 => "00111100",3210 => "11101011",3211 => "11001001",3212 => "00101000",3213 => "11101110",3214 => "10000001",3215 => "10101001",3216 => "00011110",3217 => "11000011",3218 => "00110010",3219 => "10001110",3220 => "00010001",3221 => "01001101",3222 => "11111110",3223 => "11000101",3224 => "01010010",3225 => "11100000",3226 => "01110110",3227 => "00111100",3228 => "10101100",3229 => "10011101",3230 => "10111110",3231 => "11000000",3232 => "11100011",3233 => "01110110",3234 => "01010101",3235 => "00100101",3236 => "01111011",3237 => "01110100",3238 => "00010100",3239 => "11001000",3240 => "10111100",3241 => "01101101",3242 => "01011000",3243 => "11111100",3244 => "11101110",3245 => "01110101",3246 => "10110101",3247 => "01001111",3248 => "01011000",3249 => "01001001",3250 => "00101011",3251 => "11101001",3252 => "00101011",3253 => "11011110",3254 => "11110110",3255 => "00111101",3256 => "00000001",3257 => "11111111",3258 => "01011011",3259 => "01110101",3260 => "10010010",3261 => "01010010",3262 => "10110101",3263 => "11110010",3264 => "00100101",3265 => "11101011",3266 => "00001000",3267 => "00000110",3268 => "10101000",3269 => "00010010",3270 => "01011100",3271 => "01011101",3272 => "00001111",3273 => "11110001",3274 => "11010100",3275 => "00001011",3276 => "10110110",3277 => "11011111",3278 => "11001101",3279 => "11001100",3280 => "11110000",3281 => "10010110",3282 => "00001101",3283 => "10110110",3284 => "01011100",3285 => "01010110",3286 => "11000100",3287 => "10110100",3288 => "10101100",3289 => "11001110",3290 => "11101111",3291 => "11110100",3292 => "01110010",3293 => "00001100",3294 => "00110011",3295 => "10110001",3296 => "01110111",3297 => "01110110",3298 => "01001111",3299 => "11111100",3300 => "01110111",3301 => "11000111",3302 => "10000101",3303 => "11001011",3304 => "10010010",3305 => "00110001",3306 => "00100001",3307 => "01000010",3308 => "10101001",3309 => "10101101",3310 => "11010101",3311 => "10001111",3312 => "11011001",3313 => "11100111",3314 => "00110110",3315 => "00001001",3316 => "01011010",3317 => "11111110",3318 => "10011000",3319 => "01101000",3320 => "01001100",3321 => "00000110",3322 => "11111100",3323 => "01101001",3324 => "11101111",3325 => "01110110",3326 => "10111110",3327 => "01110000",3328 => "11101100",3329 => "11100011",3330 => "10110111",3331 => "00110011",3332 => "11111011",3333 => "11001010",3334 => "11101110",3335 => "00001110",3336 => "00100111",3337 => "00111110",3338 => "00000101",3339 => "10010100",3340 => "10001010",3341 => "11011000",3342 => "01000100",3343 => "11010100",3344 => "01010001",3345 => "00000000",3346 => "00101011",3347 => "11100000",3348 => "01110110",3349 => "10111100",3350 => "11111011",3351 => "11100111",3352 => "01000011",3353 => "10111101",3354 => "10001111",3355 => "11011011",3356 => "11111011",3357 => "01100101",3358 => "00111111",3359 => "00110001",3360 => "11001111",3361 => "10000011",3362 => "10110101",3363 => "10000100",3364 => "10011010",3365 => "01101011",3366 => "00010110",3367 => "01110111",3368 => "00010011",3369 => "01110101",3370 => "11000100",3371 => "11101000",3372 => "01011000",3373 => "00111011",3374 => "11100100",3375 => "11100000",3376 => "00101110",3377 => "11001010",3378 => "11101000",3379 => "11101001",3380 => "01100110",3381 => "01111001",3382 => "11010001",3383 => "01100100",3384 => "10100010",3385 => "10110110",3386 => "10101000",3387 => "11010111",3388 => "10101101",3389 => "10010011",3390 => "11011110",3391 => "11100110",3392 => "01001001",3393 => "00111101",3394 => "10110000",3395 => "11101101",3396 => "00101001",3397 => "00000110",3398 => "11100010",3399 => "10100101",3400 => "11000001",3401 => "11100101",3402 => "11101001",3403 => "11000001",3404 => "11001100",3405 => "00010111",3406 => "10101011",3407 => "01110010",3408 => "00000011",3409 => "00110011",3410 => "10101111",3411 => "11110101",3412 => "00110111",3413 => "11011101",3414 => "01111011",3415 => "01100011",3416 => "01001101",3417 => "10001111",3418 => "10010011",3419 => "01111011",3420 => "10110110",3421 => "00010110",3422 => "01010111",3423 => "01011111",3424 => "11100011",3425 => "11110001",3426 => "01000101",3427 => "00010110",3428 => "00111110",3429 => "01010011",3430 => "11001100",3431 => "11001101",3432 => "10100001",3433 => "10101101",3434 => "01010000",3435 => "11101110",3436 => "10011100",3437 => "01010011",3438 => "11100111",3439 => "11111100",3440 => "10010010",3441 => "01011110",3442 => "10110010",3443 => "00011001",3444 => "10000011",3445 => "10101011",3446 => "00110001",3447 => "11100001",3448 => "01110100",3449 => "00011010",3450 => "10000010",3451 => "00000001",3452 => "00100111",3453 => "00010010",3454 => "11010010",3455 => "10110100",3456 => "11110001",3457 => "11100001",3458 => "01010111",3459 => "01111110",3460 => "10111000",3461 => "11010011",3462 => "00010011",3463 => "10010111",3464 => "00110100",3465 => "10000000",3466 => "00000010",3467 => "11011111",3468 => "00101111",3469 => "01011110",3470 => "11110100",3471 => "11110001",3472 => "10010001",3473 => "01101100",3474 => "10100110",3475 => "10110100",3476 => "10111101",3477 => "01000001",3478 => "01100011",3479 => "10100010",3480 => "01011101",3481 => "00000001",3482 => "01000111",3483 => "00001101",3484 => "00011001",3485 => "10000001",3486 => "01001101",3487 => "01000110",3488 => "00110011",3489 => "01110011",3490 => "10000110",3491 => "11000011",3492 => "01001111",3493 => "11101001",3494 => "01010011",3495 => "01110101",3496 => "01101111",3497 => "01010011",3498 => "11001110",3499 => "00001111",3500 => "01010000",3501 => "10001110",3502 => "00111100",3503 => "11011000",3504 => "01000000",3505 => "10111110",3506 => "00110101",3507 => "11000010",3508 => "11001101",3509 => "11110000",3510 => "00111111",3511 => "11110110",3512 => "01010100",3513 => "00001110",3514 => "01010000",3515 => "10001011",3516 => "01011101",3517 => "10000101",3518 => "11111111",3519 => "10001011",3520 => "10101110",3521 => "00101100",3522 => "11011111",3523 => "00100101",3524 => "10011001",3525 => "10110111",3526 => "01110010",3527 => "11111000",3528 => "11010100",3529 => "01001000",3530 => "01100100",3531 => "01100101",3532 => "01111111",3533 => "10010000",3534 => "00111010",3535 => "01111000",3536 => "01111000",3537 => "01110001",3538 => "00011100",3539 => "00111100",3540 => "11011100",3541 => "10011111",3542 => "10010011",3543 => "10001100",3544 => "10011110",3545 => "10101101",3546 => "00000100",3547 => "10000001",3548 => "10000011",3549 => "00000001",3550 => "00011100",3551 => "11111011",3552 => "00001110",3553 => "01111010",3554 => "10000010",3555 => "11100011",3556 => "10111011",3557 => "10001100",3558 => "00000000",3559 => "00010001",3560 => "11101011",3561 => "10111110",3562 => "10010001",3563 => "01111111",3564 => "01001100",3565 => "11100010",3566 => "01110111",3567 => "10110010",3568 => "11001001",3569 => "11001110",3570 => "01010001",3571 => "01000000",3572 => "01101010",3573 => "01101101",3574 => "00001101",3575 => "11100101",3576 => "01101000",3577 => "10001011",3578 => "00011001",3579 => "00001111",3580 => "01111010",3581 => "00100111",3582 => "00101001",3583 => "01110011",3584 => "10101100",3585 => "01010011",3586 => "01111100",3587 => "01001000",3588 => "00100111",3589 => "11111000",3590 => "00000100",3591 => "01001110",3592 => "11100000",3593 => "10011101",3594 => "00010110",3595 => "00100000",3596 => "01111101",3597 => "01101010",3598 => "01011010",3599 => "11001110",3600 => "00000101",3601 => "11110111",3602 => "11110110",3603 => "01010100",3604 => "01010000",3605 => "01101000",3606 => "00100110",3607 => "11000100",3608 => "01111101",3609 => "10010111",3610 => "00010001",3611 => "11000001",3612 => "01010110",3613 => "10110000",3614 => "10011001",3615 => "11110010",3616 => "10010100",3617 => "00000110",3618 => "10101100",3619 => "00000110",3620 => "01000110",3621 => "00100110",3622 => "01100000",3623 => "11010101",3624 => "01111100",3625 => "11011010",3626 => "10001100",3627 => "11100110",3628 => "11110110",3629 => "11111101",3630 => "10110000",3631 => "00100110",3632 => "11100000",3633 => "00000110",3634 => "01110011",3635 => "11110101",3636 => "01001010",3637 => "11011011",3638 => "00000111",3639 => "11010011",3640 => "10110001",3641 => "00010010",3642 => "01011000",3643 => "10010000",3644 => "11100100",3645 => "10110010",3646 => "00100101",3647 => "01110100",3648 => "10010100",3649 => "11111001",3650 => "00111010",3651 => "01111000",3652 => "00111101",3653 => "11010001",3654 => "11111101",3655 => "00000001",3656 => "00100100",3657 => "01100110",3658 => "00010010",3659 => "00101010",3660 => "01010011",3661 => "00011110",3662 => "01000111",3663 => "11101001",3664 => "11111010",3665 => "00011001",3666 => "00000000",3667 => "00010000",3668 => "00101001",3669 => "11111000",3670 => "11100110",3671 => "01111000",3672 => "01000011",3673 => "10100000",3674 => "01100111",3675 => "01100010",3676 => "00010000",3677 => "01011101",3678 => "11000011",3679 => "01011010",3680 => "10101111",3681 => "00001100",3682 => "10011100",3683 => "10001000",3684 => "01101011",3685 => "00010101",3686 => "00111110",3687 => "00101101",3688 => "11011011",3689 => "10010110",3690 => "00101101",3691 => "10011101",3692 => "10011001",3693 => "11110101",3694 => "01000011",3695 => "11001000",3696 => "10011110",3697 => "01000010",3698 => "01010101",3699 => "01010111",3700 => "10100111",3701 => "10000100",3702 => "00010111",3703 => "00111011",3704 => "00001110",3705 => "10111100",3706 => "10101000",3707 => "10101000",3708 => "11011011",3709 => "11011011",3710 => "11010100",3711 => "00100110",3712 => "00100100",3713 => "01011101",3714 => "01000100",3715 => "00011111",3716 => "01010110",3717 => "01101100",3718 => "00000111",3719 => "00000000",3720 => "00000011",3721 => "11111010",3722 => "10100101",3723 => "10100111",3724 => "10010101",3725 => "01011111",3726 => "01111110",3727 => "10111011",3728 => "11010010",3729 => "11001010",3730 => "11010101",3731 => "00011000",3732 => "10011111",3733 => "01011110",3734 => "01110100",3735 => "01001011",3736 => "11111101",3737 => "11001000",3738 => "00110011",3739 => "01000011",3740 => "11101010",3741 => "10000000",3742 => "11011110",3743 => "00001110",3744 => "00011110",3745 => "01110100",3746 => "01000101",3747 => "11001001",3748 => "00010010",3749 => "10111101",3750 => "00010100",3751 => "00101001",3752 => "10101110",3753 => "11000001",3754 => "11001010",3755 => "10101011",3756 => "10001000",3757 => "10001100",3758 => "11101100",3759 => "11000000",3760 => "10110111",3761 => "00001101",3762 => "01010101",3763 => "01001111",3764 => "11111011",3765 => "01001111",3766 => "10100010",3767 => "01110010",3768 => "01001111",3769 => "00011100",3770 => "01101001",3771 => "00111010",3772 => "01001101",3773 => "10010011",3774 => "11011101",3775 => "00001111",3776 => "01100010",3777 => "00110110",3778 => "01011110",3779 => "10001000",3780 => "11110011",3781 => "00011101",3782 => "10100100",3783 => "11010001",3784 => "10111110",3785 => "00101100",3786 => "10011001",3787 => "11001111",3788 => "00011101",3789 => "10101101",3790 => "01111010",3791 => "11110111",3792 => "01110100",3793 => "00111110",3794 => "10011100",3795 => "00110111",3796 => "11111110",3797 => "10110101",3798 => "00011101",3799 => "10110001",3800 => "00100011",3801 => "10111010",3802 => "10111100",3803 => "00101101",3804 => "10001110",3805 => "11011100",3806 => "11110011",3807 => "11001001",3808 => "11100101",3809 => "10110110",3810 => "11101011",3811 => "00000100",3812 => "01101101",3813 => "00110010",3814 => "00000101",3815 => "01100011",3816 => "10000110",3817 => "00110001",3818 => "11001010",3819 => "00000000",3820 => "01110000",3821 => "11101110",3822 => "10001110",3823 => "00101000",3824 => "00010101",3825 => "00000011",3826 => "01010001",3827 => "10001000",3828 => "10001010",3829 => "11110001",3830 => "11100000",3831 => "01100111",3832 => "00001111",3833 => "01100001",3834 => "00011101",3835 => "11010111",3836 => "10010010",3837 => "11111010",3838 => "01101110",3839 => "01001010",3840 => "11000011",3841 => "10111111",3842 => "00101011",3843 => "00111011",3844 => "01111101",3845 => "11101011",3846 => "00001010",3847 => "10100011",3848 => "00010100",3849 => "01101000",3850 => "10110010",3851 => "11101100",3852 => "01100010",3853 => "00001100",3854 => "01110011",3855 => "01101011",3856 => "01011100",3857 => "00010011",3858 => "00010110",3859 => "10100001",3860 => "10000111",3861 => "10100101",3862 => "11101100",3863 => "11001011",3864 => "01000100",3865 => "11010110",3866 => "00111000",3867 => "11101100",3868 => "11001100",3869 => "00001100",3870 => "00010010",3871 => "11101111",3872 => "01101011",3873 => "11000001",3874 => "00000100",3875 => "01000001",3876 => "01000011",3877 => "10000001",3878 => "00001001",3879 => "10011000",3880 => "00101000",3881 => "01111101",3882 => "10000000",3883 => "01101011",3884 => "01101110",3885 => "00010100",3886 => "11111101",3887 => "10010000",3888 => "10011010",3889 => "01011001",3890 => "11011100",3891 => "00011001",3892 => "10000101",3893 => "00111010",3894 => "10001101",3895 => "10011110",3896 => "10010111",3897 => "00000000",3898 => "01010101",3899 => "11110111",3900 => "10101011",3901 => "10010110",3902 => "00010101",3903 => "10101010",3904 => "00000101",3905 => "10100000",3906 => "10100101",3907 => "10011001",3908 => "00111110",3909 => "01110100",3910 => "00011100",3911 => "11000001",3912 => "01010110",3913 => "11100110",3914 => "01110000",3915 => "01111110",3916 => "01100110",3917 => "01001000",3918 => "01100101",3919 => "00111011",3920 => "10100011",3921 => "10100101",3922 => "01011010",3923 => "01111011",3924 => "10101000",3925 => "00000110",3926 => "11111000",3927 => "00001110",3928 => "10100110",3929 => "11001011",3930 => "10101111",3931 => "11011110",3932 => "00110100",3933 => "10010010",3934 => "11101000",3935 => "00000110",3936 => "10000000",3937 => "00111001",3938 => "01100101",3939 => "10110011",3940 => "11001100",3941 => "10000001",3942 => "01101101",3943 => "00111000",3944 => "00111111",3945 => "11010010",3946 => "00101111",3947 => "11011111",3948 => "01111101",3949 => "01000110",3950 => "10111100",3951 => "11000101",3952 => "01001111",3953 => "11100011",3954 => "10111000",3955 => "00111001",3956 => "01100011",3957 => "11011000",3958 => "01010001",3959 => "11111000",3960 => "10001110",3961 => "00100000",3962 => "01010000",3963 => "10000000",3964 => "01111101",3965 => "01100111",3966 => "01111110",3967 => "00100000",3968 => "01100101",3969 => "11011011",3970 => "10011111",3971 => "10110011",3972 => "01111010",3973 => "11110111",3974 => "00111001",3975 => "01000000",3976 => "11011011",3977 => "11101110",3978 => "01101000",3979 => "01101110",3980 => "00110101",3981 => "11000001",3982 => "10100001",3983 => "01101101",3984 => "11001001",3985 => "01000010",3986 => "11101001",3987 => "01101011",3988 => "00001111",3989 => "01010110",3990 => "00101011",3991 => "00000000",3992 => "00011011",3993 => "10100101",3994 => "10111010",3995 => "11111010",3996 => "00111101",3997 => "00001001",3998 => "01101110",3999 => "00000110",4000 => "11100101",4001 => "11010001",4002 => "10011011",4003 => "00011111",4004 => "10111110",4005 => "10111000",4006 => "10010011",4007 => "01010100",4008 => "11110000",4009 => "00010100",4010 => "10111100",4011 => "00100011",4012 => "01100010",4013 => "10100110",4014 => "00100000",4015 => "11001001",4016 => "10011101",4017 => "10001101",4018 => "00101110",4019 => "11010101",4020 => "11101111",4021 => "10110001",4022 => "10010100",4023 => "00011110",4024 => "10000001",4025 => "10101010",4026 => "10101011",4027 => "10001011",4028 => "01101111",4029 => "01111001",4030 => "11001111",4031 => "01011000",4032 => "10110110",4033 => "11101011",4034 => "11001101",4035 => "11111111",4036 => "00110111",4037 => "11100011",4038 => "10110001",4039 => "00101100",4040 => "01000001",4041 => "11110100",4042 => "00111110",4043 => "11010110",4044 => "00100011",4045 => "11110110",4046 => "10100100",4047 => "11001010",4048 => "00111001",4049 => "11001011",4050 => "01110001",4051 => "10110010",4052 => "10011001",4053 => "11000010",4054 => "01111100",4055 => "01101001",4056 => "01111110",4057 => "11000111",4058 => "00000000",4059 => "00100101",4060 => "11010110",4061 => "11001101",4062 => "00000011",4063 => "00111101",4064 => "01001101",4065 => "01011111",4066 => "00111111",4067 => "01001010",4068 => "01000100",4069 => "11011001",4070 => "10001101",4071 => "10001101",4072 => "11100101",4073 => "10010000",4074 => "10010110",4075 => "00001110",4076 => "01001000",4077 => "01110010",4078 => "10100100",4079 => "10011011",4080 => "10111110",4081 => "11100000",4082 => "10101011",4083 => "00111011",4084 => "10000111",4085 => "11000001",4086 => "11000110",4087 => "01000110",4088 => "10000110",4089 => "11000100",4090 => "00000011",4091 => "01011000",4092 => "10011100",4093 => "00100101",4094 => "01100111",4095 => "01011111",4096 => "01000110",4097 => "10100100",4098 => "00010101",4099 => "11101011",4100 => "10111111",4101 => "00011001",4102 => "01101001",4103 => "10010011",4104 => "00011100",4105 => "01111011",4106 => "00000000",4107 => "00011111",4108 => "00100111",4109 => "10010011",4110 => "01101011",4111 => "00110010",4112 => "11111001",4113 => "01100100",4114 => "10111000",4115 => "01010100",4116 => "11110010",4117 => "01000000",4118 => "01111000",4119 => "10010110",4120 => "11000100",4121 => "01101011",4122 => "00011000",4123 => "01000001",4124 => "10011100",4125 => "01100110",4126 => "00101100",4127 => "10010110",4128 => "10110000",4129 => "00001110",4130 => "10100000",4131 => "00000101",4132 => "00000101",4133 => "00011011",4134 => "00110110",4135 => "00100010",4136 => "00000010",4137 => "01000111",4138 => "01000010",4139 => "00101010",4140 => "00010011",4141 => "10111100",4142 => "00011101",4143 => "10101111",4144 => "00100001",4145 => "11101011",4146 => "11110000",4147 => "00100111",4148 => "01001100",4149 => "01001111",4150 => "00001111",4151 => "01010111",4152 => "01010100",4153 => "00101110",4154 => "10101001",4155 => "10100010",4156 => "10000101",4157 => "10000000",4158 => "01100010",4159 => "01000101",4160 => "00010110",4161 => "01000100",4162 => "01111100",4163 => "00001111",4164 => "11110001",4165 => "10010110",4166 => "10101010",4167 => "11000001",4168 => "01011001",4169 => "10001100",4170 => "11111111",4171 => "00011110",4172 => "00101101",4173 => "01110001",4174 => "10011110",4175 => "01101110",4176 => "10111010",4177 => "10101101",4178 => "00111111",4179 => "11001100",4180 => "00001000",4181 => "10110001",4182 => "00100111",4183 => "11111111",4184 => "11001011",4185 => "01011111",4186 => "10010001",4187 => "10101100",4188 => "01010001",4189 => "00100011",4190 => "00000001",4191 => "11010111",4192 => "01100110",4193 => "11011111",4194 => "00011011",4195 => "00000010",4196 => "10001101",4197 => "10110001",4198 => "01111010",4199 => "01010100",4200 => "11101001",4201 => "00010110",4202 => "10100000",4203 => "00110100",4204 => "11110001",4205 => "01100111",4206 => "00000111",4207 => "00100110",4208 => "00011101",4209 => "00100111",4210 => "00110011",4211 => "01001001",4212 => "11001101",4213 => "11010110",4214 => "01101100",4215 => "01000000",4216 => "10110101",4217 => "11110011",4218 => "01110010",4219 => "11011000",4220 => "11100101",4221 => "01011111",4222 => "11000110",4223 => "10010010",4224 => "10010110",4225 => "10111101",4226 => "10111110",4227 => "01001111",4228 => "01010010",4229 => "00100011",4230 => "00100100",4231 => "10110100",4232 => "11110011",4233 => "11111010",4234 => "10000111",4235 => "10110001",4236 => "01001111",4237 => "11001110",4238 => "01001011",4239 => "01011001",4240 => "10110010",4241 => "01100101",4242 => "00100110",4243 => "10110001",4244 => "00011001",4245 => "01001011",4246 => "00111101",4247 => "11011101",4248 => "10000000",4249 => "11101110",4250 => "00100010",4251 => "00011000",4252 => "00101001",4253 => "01110001",4254 => "10101110",4255 => "01110010",4256 => "10001000",4257 => "00101000",4258 => "11111101",4259 => "00100001",4260 => "11011001",4261 => "01101110",4262 => "11100111",4263 => "10010101",4264 => "11111111",4265 => "00000010",4266 => "00011011",4267 => "01011110",4268 => "10001101",4269 => "00111101",4270 => "11111111",4271 => "10011100",4272 => "10001001",4273 => "01100101",4274 => "01000011",4275 => "10001000",4276 => "11001000",4277 => "10101001",4278 => "00110000",4279 => "10111101",4280 => "10011110",4281 => "01011111",4282 => "10011010",4283 => "01000101",4284 => "10100011",4285 => "01101101",4286 => "00110001",4287 => "01010001",4288 => "10111110",4289 => "10111111",4290 => "11010000",4291 => "11000111",4292 => "01011100",4293 => "01111000",4294 => "10100111",4295 => "11100110",4296 => "10110010",4297 => "10001110",4298 => "11100100",4299 => "10110001",4300 => "00110110",4301 => "10100011",4302 => "00001001",4303 => "01011100",4304 => "01110100",4305 => "11011001",4306 => "11101100",4307 => "01001101",4308 => "10101011",4309 => "00111001",4310 => "01000100",4311 => "11000000",4312 => "00111101",4313 => "01001010",4314 => "01101000",4315 => "00010101",4316 => "00100111",4317 => "01101001",4318 => "01001001",4319 => "11101111",4320 => "10111000",4321 => "10000110",4322 => "01111001",4323 => "11000100",4324 => "00000110",4325 => "00100000",4326 => "11001011",4327 => "11100011",4328 => "11110111",4329 => "01100010",4330 => "11101010",4331 => "11111110",4332 => "11110101",4333 => "00110001",4334 => "01000001",4335 => "10101011",4336 => "01101111",4337 => "11001101",4338 => "10010101",4339 => "00110001",4340 => "10010100",4341 => "10100110",4342 => "00000011",4343 => "01101101",4344 => "01101000",4345 => "10011011",4346 => "00100010",4347 => "00101100",4348 => "10000101",4349 => "10100111",4350 => "01100100",4351 => "11010110",4352 => "10011101",4353 => "00010011",4354 => "00000111",4355 => "11001111",4356 => "01011100",4357 => "01010001",4358 => "10011101",4359 => "11111110",4360 => "11001110",4361 => "10001101",4362 => "10001011",4363 => "01101110",4364 => "01100110",4365 => "00110010",4366 => "01010011",4367 => "00010011",4368 => "11101010",4369 => "00101011",4370 => "00010011",4371 => "10101001",4372 => "01110000",4373 => "01110111",4374 => "01000000",4375 => "01100111",4376 => "00000101",4377 => "01111101",4378 => "11100001",4379 => "00000010",4380 => "00011101",4381 => "01110001",4382 => "10010100",4383 => "01001100",4384 => "01110110",4385 => "01101101",4386 => "00001000",4387 => "00101011",4388 => "01110101",4389 => "01011111",4390 => "11101101",4391 => "10000100",4392 => "01101000",4393 => "10101010",4394 => "01110000",4395 => "11111110",4396 => "00011001",4397 => "11110001",4398 => "00100100",4399 => "01010000",4400 => "00010010",4401 => "00001011",4402 => "00001111",4403 => "01011111",4404 => "10011110",4405 => "10111011",4406 => "01001100",4407 => "01000100",4408 => "11101110",4409 => "11110111",4410 => "01111110",4411 => "11101001",4412 => "11011100",4413 => "01100101",4414 => "01111010",4415 => "10001001",4416 => "01100100",4417 => "10000111",4418 => "10101100",4419 => "01010000",4420 => "10101010",4421 => "11010010",4422 => "00010101",4423 => "00000101",4424 => "01100010",4425 => "10000001",4426 => "01000001",4427 => "10000000",4428 => "00011101",4429 => "11100000",4430 => "01110111",4431 => "00001001",4432 => "10101111",4433 => "00001010",4434 => "11010100",4435 => "00100010",4436 => "10011110",4437 => "10000010",4438 => "01011011",4439 => "00101101",4440 => "10100000",4441 => "00111000",4442 => "00100011",4443 => "00011110",4444 => "00110110",4445 => "01111001",4446 => "11101011",4447 => "01000010",4448 => "01110011",4449 => "10010011",4450 => "00111001",4451 => "00000011",4452 => "01010001",4453 => "10110101",4454 => "00101111",4455 => "10001000",4456 => "10011110",4457 => "10010101",4458 => "10000001",4459 => "01100011",4460 => "11100101",4461 => "00010110",4462 => "01010010",4463 => "11001111",4464 => "10110010",4465 => "10101111",4466 => "10011001",4467 => "10100011",4468 => "00111001",4469 => "11001011",4470 => "00010111",4471 => "01011010",4472 => "11000101",4473 => "00110000",4474 => "10101000",4475 => "00011110",4476 => "00111110",4477 => "11000111",4478 => "11011011",4479 => "10111100",4480 => "00000101",4481 => "01111011",4482 => "10001110",4483 => "00100101",4484 => "00110000",4485 => "11010000",4486 => "01110001",4487 => "00100001",4488 => "01100011",4489 => "01101101",4490 => "11100011",4491 => "00111011",4492 => "10100110",4493 => "11110100",4494 => "01001101",4495 => "11101101",4496 => "11111101",4497 => "01000101",4498 => "01110010",4499 => "00011000",4500 => "10001101",4501 => "11010111",4502 => "00000000",4503 => "10000101",4504 => "01110000",4505 => "01100100",4506 => "10100111",4507 => "10011011",4508 => "11011111",4509 => "10000111",4510 => "01101110",4511 => "00110101",4512 => "01010010",4513 => "10000101",4514 => "00000101",4515 => "10110000",4516 => "00010111",4517 => "01101111",4518 => "10101010",4519 => "00101111",4520 => "00000110",4521 => "11110111",4522 => "10100111",4523 => "10011110",4524 => "00101001",4525 => "10011011",4526 => "01100010",4527 => "00000110",4528 => "10100010",4529 => "10010010",4530 => "00100110",4531 => "11000010",4532 => "11101010",4533 => "11000001",4534 => "11100100",4535 => "01011010",4536 => "01110001",4537 => "11111001",4538 => "11100011",4539 => "10110011",4540 => "00000101",4541 => "00100011",4542 => "10100010",4543 => "00101100",4544 => "11101111",4545 => "00110111",4546 => "11001110",4547 => "01100111",4548 => "11001000",4549 => "01001001",4550 => "01100001",4551 => "10000011",4552 => "11110010",4553 => "10000110",4554 => "10110011",4555 => "01011000",4556 => "01110100",4557 => "11100001",4558 => "00100010",4559 => "00110011",4560 => "01011110",4561 => "10001010",4562 => "01001001",4563 => "01110101",4564 => "00111001",4565 => "10101011",4566 => "11001000",4567 => "10101001",4568 => "11000010",4569 => "01000100",4570 => "11110010",4571 => "11011100",4572 => "01111000",4573 => "11010110",4574 => "00001110",4575 => "11000010",4576 => "00001100",4577 => "11110010",4578 => "10001000",4579 => "10111100",4580 => "10000111",4581 => "00100100",4582 => "11011110",4583 => "01000100",4584 => "10011111",4585 => "11010101",4586 => "01011010",4587 => "10111110",4588 => "00100111",4589 => "11010111",4590 => "11110101",4591 => "11001101",4592 => "01011101",4593 => "01111011",4594 => "01000000",4595 => "11011000",4596 => "10001110",4597 => "01001100",4598 => "01111101",4599 => "00010111",4600 => "00000001",4601 => "01101010",4602 => "10100001",4603 => "01101100",4604 => "10011101",4605 => "00111111",4606 => "01111010",4607 => "10110001",4608 => "00000011",4609 => "00110001",4610 => "11100000",4611 => "00101101",4612 => "01000010",4613 => "11110101",4614 => "01101010",4615 => "00110111",4616 => "01111001",4617 => "01000011",4618 => "01111110",4619 => "10000111",4620 => "00101110",4621 => "00001110",4622 => "00010010",4623 => "00110110",4624 => "00010110",4625 => "11111111",4626 => "01010001",4627 => "00111000",4628 => "01001100",4629 => "00100011",4630 => "01101010",4631 => "10101001",4632 => "11011011",4633 => "11110011",4634 => "11110010",4635 => "10111011",4636 => "00010000",4637 => "01011010",4638 => "11001100",4639 => "01111101",4640 => "00000100",4641 => "10001000",4642 => "01101111",4643 => "11101111",4644 => "11101110",4645 => "00000110",4646 => "01010111",4647 => "11011101",4648 => "11110010",4649 => "11101110",4650 => "01000101",4651 => "10111010",4652 => "10110111",4653 => "10001010",4654 => "10110100",4655 => "00100011",4656 => "10011011",4657 => "10010010",4658 => "00000010",4659 => "10010010",4660 => "11111010",4661 => "01111010",4662 => "01011111",4663 => "11110101",4664 => "10010001",4665 => "10110010",4666 => "11011100",4667 => "01100010",4668 => "01101000",4669 => "01011101",4670 => "10011001",4671 => "01110000",4672 => "11111001",4673 => "01011000",4674 => "00101101",4675 => "11101001",4676 => "10000101",4677 => "11011011",4678 => "01000000",4679 => "00101001",4680 => "10101000",4681 => "00101100",4682 => "00010100",4683 => "11100111",4684 => "01111110",4685 => "01000010",4686 => "10001000",4687 => "11000100",4688 => "00111100",4689 => "11001010",4690 => "00001001",4691 => "11110011",4692 => "10001001",4693 => "11001010",4694 => "00111001",4695 => "11100001",4696 => "10111011",4697 => "10011110",4698 => "00010001",4699 => "00110001",4700 => "01111111",4701 => "10110100",4702 => "01011010",4703 => "11111111",4704 => "11000101",4705 => "11001100",4706 => "00001101",4707 => "00010000",4708 => "01100100",4709 => "00101101",4710 => "01011011",4711 => "10001010",4712 => "00100000",4713 => "00010001",4714 => "10110001",4715 => "10011010",4716 => "10001010",4717 => "11100101",4718 => "00101011",4719 => "10000010",4720 => "01100110",4721 => "10011100",4722 => "00101110",4723 => "01000011",4724 => "00110001",4725 => "10100110",4726 => "00111001",4727 => "10111100",4728 => "01111111",4729 => "10011001",4730 => "10010100",4731 => "10001011",4732 => "01111100",4733 => "01110101",4734 => "10110111",4735 => "01110001",4736 => "10001010",4737 => "01001000",4738 => "00000111",4739 => "00001100",4740 => "11010111",4741 => "11000000",4742 => "00101010",4743 => "01101100",4744 => "01101111",4745 => "10010110",4746 => "01100001",4747 => "10011111",4748 => "00000110",4749 => "11101101",4750 => "10111000",4751 => "11001010",4752 => "10010000",4753 => "11011100",4754 => "01101011",4755 => "10011110",4756 => "00010000",4757 => "00110011",4758 => "01110000",4759 => "10011101",4760 => "11100111",4761 => "10111010",4762 => "10101110",4763 => "11000010",4764 => "01110110",4765 => "00010100",4766 => "01110010",4767 => "10011010",4768 => "10101111",4769 => "01011101",4770 => "01110011",4771 => "11100100",4772 => "11101000",4773 => "01111000",4774 => "10001000",4775 => "10101001",4776 => "10011010",4777 => "00101011",4778 => "10000000",4779 => "10000101",4780 => "10111100",4781 => "10111111",4782 => "01010010",4783 => "01111110",4784 => "11110111",4785 => "00010110",4786 => "11011001",4787 => "00010111",4788 => "00011101",4789 => "10101001",4790 => "00111011",4791 => "00000101",4792 => "11111111",4793 => "00111001",4794 => "01101111",4795 => "01011110",4796 => "00111001",4797 => "01000011",4798 => "11010011",4799 => "11111010",4800 => "00100110",4801 => "00000011",4802 => "01001101",4803 => "01110010",4804 => "11100111",4805 => "01100110",4806 => "11101111",4807 => "00010100",4808 => "00111011",4809 => "00011010",4810 => "00111110",4811 => "11111010",4812 => "11011000",4813 => "00110010",4814 => "10110110",4815 => "01111110",4816 => "10100011",4817 => "01001000",4818 => "10111000",4819 => "01000100",4820 => "10010011",4821 => "01111000",4822 => "00110001",4823 => "11100100",4824 => "11110010",4825 => "00101110",4826 => "11000010",4827 => "01111010",4828 => "01001110",4829 => "00010110",4830 => "00010110",4831 => "11100110",4832 => "00000001",4833 => "01000101",4834 => "11111101",4835 => "10000001",4836 => "00111110",4837 => "11001110",4838 => "10001100",4839 => "01110110",4840 => "11101100",4841 => "01101110",4842 => "00000010",4843 => "01000110",4844 => "01111011",4845 => "10110110",4846 => "11111001",4847 => "01010001",4848 => "00100011",4849 => "10100101",4850 => "00101011",4851 => "00000010",4852 => "11111011",4853 => "10000111",4854 => "10101011",4855 => "10100001",4856 => "11000100",4857 => "11111001",4858 => "01010010",4859 => "00010111",4860 => "01101011",4861 => "01100010",4862 => "00111101",4863 => "00011000",4864 => "00111010",4865 => "11101101",4866 => "00100001",4867 => "00111011",4868 => "10000111",4869 => "01110000",4870 => "10010100",4871 => "00110010",4872 => "11100001",4873 => "00100010",4874 => "10110111",4875 => "11110011",4876 => "01101101",4877 => "10101100",4878 => "00000100",4879 => "11010110",4880 => "11100101",4881 => "00110000",4882 => "00011100",4883 => "11000011",4884 => "11100110",4885 => "00011000",4886 => "01000000",4887 => "01110111",4888 => "01000010",4889 => "00101110",4890 => "00111000",4891 => "00010111",4892 => "01101111",4893 => "11101101",4894 => "11101001",4895 => "10110100",4896 => "01010010",4897 => "00101011",4898 => "00000010",4899 => "11000101",4900 => "11000011",4901 => "11110000",4902 => "11011011",4903 => "10111100",4904 => "11010101",4905 => "10110010",4906 => "11110000",4907 => "11111111",4908 => "11011111",4909 => "00111111",4910 => "00010000",4911 => "00011001",4912 => "10111011",4913 => "01101100",4914 => "00001100",4915 => "01011011",4916 => "10001010",4917 => "11000010",4918 => "10000000",4919 => "10000100",4920 => "01000000",4921 => "00000000",4922 => "01111000",4923 => "10001101",4924 => "00100101",4925 => "10000011",4926 => "01110001",4927 => "01011101",4928 => "00000011",4929 => "10110000",4930 => "01100001",4931 => "01001111",4932 => "11011110",4933 => "11110010",4934 => "10100000",4935 => "10000111",4936 => "00110100",4937 => "00010011",4938 => "11001111",4939 => "01100101",4940 => "10100101",4941 => "10111101",4942 => "10001011",4943 => "00110101",4944 => "00101001",4945 => "10010011",4946 => "00111000",4947 => "11010111",4948 => "10111100",4949 => "01010010",4950 => "01010011",4951 => "10111011",4952 => "10111010",4953 => "11111110",4954 => "00001000",4955 => "10100100",4956 => "00011011",4957 => "10100011",4958 => "00100000",4959 => "00010010",4960 => "10010110",4961 => "01110101",4962 => "01101101",4963 => "00100110",4964 => "00110001",4965 => "00100111",4966 => "10101110",4967 => "00111000",4968 => "00001000",4969 => "10011110",4970 => "10011001",4971 => "01001110",4972 => "10101110",4973 => "01110111",4974 => "00010100",4975 => "01110010",4976 => "11100001",4977 => "10010000",4978 => "10110010",4979 => "01111110",4980 => "00110001",4981 => "11100111",4982 => "01010011",4983 => "00100101",4984 => "00100010",4985 => "10111010",4986 => "10110001",4987 => "01100010",4988 => "00000101",4989 => "10100000",4990 => "01000100",4991 => "11000111",4992 => "00001001",4993 => "00101011",4994 => "01110101",4995 => "10011101",4996 => "10101101",4997 => "10111001",4998 => "10101001",4999 => "01110001",5000 => "11010101",5001 => "11010100",5002 => "01001010",5003 => "10110000",5004 => "01011100",5005 => "00001010",5006 => "01001001",5007 => "00001101",5008 => "10011010",5009 => "11001000",5010 => "00111001",5011 => "11001110",5012 => "01001100",5013 => "11101101",5014 => "01001111",5015 => "01011100",5016 => "01111010",5017 => "00010011",5018 => "01111000",5019 => "11010101",5020 => "11011010",5021 => "11100001",5022 => "11000111",5023 => "00100101",5024 => "11000010",5025 => "10001010",5026 => "11001101",5027 => "11010111",5028 => "10010000",5029 => "01000101",5030 => "11000000",5031 => "10101100",5032 => "01100100",5033 => "10111001",5034 => "01000110",5035 => "00111010",5036 => "11110101",5037 => "01000000",5038 => "11010001",5039 => "01000000",5040 => "01110101",5041 => "11001101",5042 => "01110000",5043 => "00010011",5044 => "10000101",5045 => "01101001",5046 => "11101111",5047 => "01000000",5048 => "01010111",5049 => "01111011",5050 => "01000001",5051 => "11000010",5052 => "10110011",5053 => "10000011",5054 => "01000000",5055 => "01000101",5056 => "11111100",5057 => "11001000",5058 => "00100001",5059 => "10001011",5060 => "00010101",5061 => "00111000",5062 => "00001010",5063 => "10000111",5064 => "11110001",5065 => "10101011",5066 => "00001001",5067 => "00011110",5068 => "01111111",5069 => "01101010",5070 => "11111101",5071 => "10110001",5072 => "00111011",5073 => "11000010",5074 => "11101000",5075 => "01011010",5076 => "00100100",5077 => "11100111",5078 => "10010101",5079 => "11000111",5080 => "10111100",5081 => "10011000",5082 => "00000001",5083 => "00101110",5084 => "10110000",5085 => "01010000",5086 => "10011111",5087 => "10001000",5088 => "10100111",5089 => "11101110",5090 => "10101010",5091 => "10100111",5092 => "10110111",5093 => "00111011",5094 => "11111110",5095 => "11000101",5096 => "01000000",5097 => "11100001",5098 => "11001111",5099 => "00100100",5100 => "11111101",5101 => "01100000",5102 => "10111000",5103 => "00000101",5104 => "10101111",5105 => "00101111",5106 => "00000110",5107 => "10010010",5108 => "10001001",5109 => "01110101",5110 => "01000011",5111 => "10100110",5112 => "01000010",5113 => "01011010",5114 => "11011001",5115 => "10110000",5116 => "00110111",5117 => "00010100",5118 => "01111011",5119 => "10110111",5120 => "00011000",5121 => "00000100",5122 => "00101010",5123 => "01111110",5124 => "01001111",5125 => "10001101",5126 => "11111101",5127 => "11000101",5128 => "10100001",5129 => "10110011",5130 => "10101110",5131 => "00011111",5132 => "01101110",5133 => "01011000",5134 => "11110010",5135 => "01110010",5136 => "10100101",5137 => "01111100",5138 => "01011110",5139 => "00100001",5140 => "00011100",5141 => "00111111",5142 => "00010110",5143 => "10000101",5144 => "00100010",5145 => "11010011",5146 => "10011011",5147 => "10100101",5148 => "11110111",5149 => "01011001",5150 => "00001100",5151 => "01000001",5152 => "01000100",5153 => "11100010",5154 => "11010011",5155 => "10001011",5156 => "00011010",5157 => "00010011",5158 => "00001110",5159 => "10011100",5160 => "10011110",5161 => "10111010",5162 => "00101111",5163 => "10111110",5164 => "10110111",5165 => "10100001",5166 => "01010010",5167 => "01101001",5168 => "10101000",5169 => "01001110",5170 => "01100111",5171 => "01110100",5172 => "01001100",5173 => "00000001",5174 => "00100001",5175 => "01000101",5176 => "01011111",5177 => "00101111",5178 => "11001111",5179 => "00111001",5180 => "01101010",5181 => "00001000",5182 => "01011000",5183 => "10011011",5184 => "00000010",5185 => "01100111",5186 => "00011000",5187 => "10101100",5188 => "01010110",5189 => "00110000",5190 => "00000011",5191 => "11101010",5192 => "11001001",5193 => "01100010",5194 => "01000111",5195 => "11100010",5196 => "11001010",5197 => "00101101",5198 => "01101110",5199 => "01001101",5200 => "00010011",5201 => "01110010",5202 => "10111010",5203 => "10001101",5204 => "11010110",5205 => "11100101",5206 => "01110000",5207 => "01110000",5208 => "00000001",5209 => "01010100",5210 => "11100011",5211 => "10110110",5212 => "01110110",5213 => "10010010",5214 => "10101010",5215 => "11111010",5216 => "01000011",5217 => "01111100",5218 => "11011001",5219 => "00000110",5220 => "10001000",5221 => "11111100",5222 => "00000101",5223 => "11111100",5224 => "00011001",5225 => "10011011",5226 => "10010101",5227 => "10100111",5228 => "01001001",5229 => "01000010",5230 => "01000101",5231 => "00001111",5232 => "01011011",5233 => "01110100",5234 => "00111010",5235 => "10110110",5236 => "00100110",5237 => "01011001",5238 => "10001111",5239 => "11110101",5240 => "00110101",5241 => "11111111",5242 => "00000000",5243 => "00010011",5244 => "11000101",5245 => "00110000",5246 => "10111010",5247 => "01011100",5248 => "00001000",5249 => "00111001",5250 => "01100010",5251 => "10011010",5252 => "01000100",5253 => "11000000",5254 => "01111110",5255 => "11100010",5256 => "10110110",5257 => "00110100",5258 => "11001100",5259 => "11110001",5260 => "00001110",5261 => "00001011",5262 => "00101101",5263 => "00100010",5264 => "10110001",5265 => "00001111",5266 => "11010011",5267 => "11010101",5268 => "00100010",5269 => "01000101",5270 => "00111111",5271 => "01101010",5272 => "10100011",5273 => "10001100",5274 => "10111110",5275 => "00110100",5276 => "11011001",5277 => "10101011",5278 => "01111010",5279 => "10110100",5280 => "00111010",5281 => "11111010",5282 => "01111001",5283 => "01110100",5284 => "11100010",5285 => "00110000",5286 => "00000001",5287 => "11001100",5288 => "11101000",5289 => "10111001",5290 => "01011100",5291 => "10110100",5292 => "01100000",5293 => "10101100",5294 => "11000000",5295 => "01100110",5296 => "10001100",5297 => "00111101",5298 => "10100111",5299 => "11101111",5300 => "01110000",5301 => "01000001",5302 => "11101101",5303 => "10011110",5304 => "10110111",5305 => "00101111",5306 => "11111100",5307 => "11111100",5308 => "01011000",5309 => "10100011",5310 => "11000101",5311 => "00001011",5312 => "10110100",5313 => "00001011",5314 => "01001010",5315 => "01000000",5316 => "00010101",5317 => "11011001",5318 => "01110011",5319 => "11111111",5320 => "01110010",5321 => "01000011",5322 => "01101111",5323 => "11011000",5324 => "01001111",5325 => "00110101",5326 => "11111100",5327 => "01011111",5328 => "11110000",5329 => "11001111",5330 => "01010001",5331 => "10101101",5332 => "10100011",5333 => "01000100",5334 => "00111001",5335 => "10011110",5336 => "11001110",5337 => "00000011",5338 => "00010100",5339 => "00011101",5340 => "11111010",5341 => "11000011",5342 => "11010010",5343 => "00011111",5344 => "11111100",5345 => "11101010",5346 => "01000100",5347 => "00010110",5348 => "01110111",5349 => "11001011",5350 => "00100011",5351 => "01010010",5352 => "01000110",5353 => "11101000",5354 => "00000010",5355 => "11011111",5356 => "00100010",5357 => "01010000",5358 => "10011011",5359 => "01011110",5360 => "10100111",5361 => "11001111",5362 => "00100110",5363 => "10000000",5364 => "11011101",5365 => "00101110",5366 => "00000011",5367 => "01010100",5368 => "10111101",5369 => "10010010",5370 => "11001101",5371 => "00000001",5372 => "00111001",5373 => "00100111",5374 => "00100100",5375 => "10110100",5376 => "00000001",5377 => "00011101",5378 => "01101100",5379 => "00000001",5380 => "11100001",5381 => "01010010",5382 => "01101110",5383 => "11010101",5384 => "01000000",5385 => "01000100",5386 => "00010010",5387 => "01110000",5388 => "00000000",5389 => "01110110",5390 => "10101110",5391 => "11000101",5392 => "00010011",5393 => "01011110",5394 => "10010100",5395 => "11000000",5396 => "01010010",5397 => "11100110",5398 => "10001011",5399 => "01101110",5400 => "11100000",5401 => "00011010",5402 => "01111101",5403 => "01001100",5404 => "11100010",5405 => "11010011",5406 => "10100011",5407 => "00000000",5408 => "00110100",5409 => "00000100",5410 => "01100001",5411 => "01000111",5412 => "00100000",5413 => "11111110",5414 => "11000010",5415 => "10011111",5416 => "11000011",5417 => "00001100",5418 => "11010000",5419 => "00011011",5420 => "00111011",5421 => "00000000",5422 => "10011101",5423 => "00110010",5424 => "11011001",5425 => "01100111",5426 => "00010111",5427 => "10011001",5428 => "01000000",5429 => "00011111",5430 => "00111001",5431 => "11101010",5432 => "11101100",5433 => "00000000",5434 => "11110110",5435 => "01110100",5436 => "01000010",5437 => "00011111",5438 => "11000101",5439 => "00011111",5440 => "01001110",5441 => "00011001",5442 => "01110100",5443 => "01101011",5444 => "11101000",5445 => "00001011",5446 => "00100110",5447 => "10111111",5448 => "00101010",5449 => "01001010",5450 => "00100101",5451 => "00110111",5452 => "10110111",5453 => "01101100",5454 => "01110010",5455 => "01111011",5456 => "11010101",5457 => "01100101",5458 => "00100100",5459 => "00111101",5460 => "11011010",5461 => "10011101",5462 => "10111010",5463 => "00110010",5464 => "01000010",5465 => "10001111",5466 => "01111001",5467 => "01000110",5468 => "11101011",5469 => "01101101",5470 => "01000010",5471 => "10010110",5472 => "10101100",5473 => "10110000",5474 => "01001000",5475 => "00000011",5476 => "10110010",5477 => "10101101",5478 => "10100010",5479 => "01110011",5480 => "01001000",5481 => "10101000",5482 => "11011110",5483 => "11101111",5484 => "11001011",5485 => "10110011",5486 => "10000101",5487 => "11011001",5488 => "10000111",5489 => "11010011",5490 => "01001100",5491 => "10101100",5492 => "00000000",5493 => "00100011",5494 => "11000100",5495 => "00011000",5496 => "00011000",5497 => "01010110",5498 => "01000010",5499 => "10001101",5500 => "00110111",5501 => "00010111",5502 => "11011111",5503 => "10011001",5504 => "11001110",5505 => "11010101",5506 => "00111001",5507 => "01101011",5508 => "01100000",5509 => "11111001",5510 => "01010110",5511 => "00111000",5512 => "01101110",5513 => "10100011",5514 => "11111110",5515 => "00010100",5516 => "11110110",5517 => "00111011",5518 => "00110101",5519 => "10101000",5520 => "10100111",5521 => "01011011",5522 => "00110111",5523 => "01110111",5524 => "11000100",5525 => "10111010",5526 => "10010101",5527 => "00100010",5528 => "10001000",5529 => "10110110",5530 => "11111001",5531 => "01010111",5532 => "01011011",5533 => "01100100",5534 => "11000111",5535 => "11111000",5536 => "00000101",5537 => "11111111",5538 => "00101110",5539 => "11110001",5540 => "11001100",5541 => "01101111",5542 => "10101111",5543 => "11100010",5544 => "11100101",5545 => "01100011",5546 => "11101100",5547 => "01001001",5548 => "11110000",5549 => "10010111",5550 => "10101100",5551 => "00000011",5552 => "10001100",5553 => "10000100",5554 => "11111111",5555 => "10010010",5556 => "11110000",5557 => "00001000",5558 => "11011011",5559 => "10001100",5560 => "10101010",5561 => "11100111",5562 => "10111001",5563 => "01011000",5564 => "11010001",5565 => "00101001",5566 => "10110100",5567 => "00011101",5568 => "11011101",5569 => "01100000",5570 => "01110110",5571 => "11100000",5572 => "00011010",5573 => "11111100",5574 => "11001000",5575 => "10001110",5576 => "01001010",5577 => "11011010",5578 => "11101000",5579 => "01010111",5580 => "11111001",5581 => "11100110",5582 => "01111101",5583 => "11110001",5584 => "01001011",5585 => "11010010",5586 => "10101110",5587 => "00001100",5588 => "00011001",5589 => "01000111",5590 => "00100001",5591 => "01001011",5592 => "11010001",5593 => "11001100",5594 => "00001111",5595 => "01001011",5596 => "01010110",5597 => "00110001",5598 => "00100110",5599 => "11000101",5600 => "00011011",5601 => "11000011",5602 => "01101101",5603 => "10100111",5604 => "00111101",5605 => "11011000",5606 => "01110010",5607 => "11111001",5608 => "01011111",5609 => "01111010",5610 => "10010100",5611 => "00110101",5612 => "01101100",5613 => "10100100",5614 => "11011000",5615 => "01001011",5616 => "01011110",5617 => "00011111",5618 => "11110100",5619 => "00011011",5620 => "01010001",5621 => "01010000",5622 => "00010011",5623 => "11011100",5624 => "00011011",5625 => "00111111",5626 => "10000000",5627 => "10010111",5628 => "11100010",5629 => "01010101",5630 => "01011011",5631 => "10010000",5632 => "11100100",5633 => "11001110",5634 => "01000011",5635 => "01110101",5636 => "10001100",5637 => "01101101",5638 => "10101100",5639 => "00100010",5640 => "11001011",5641 => "11000000",5642 => "00110100",5643 => "11010110",5644 => "11001000",5645 => "01001000",5646 => "00110000",5647 => "01000001",5648 => "10000001",5649 => "00110010",5650 => "01100000",5651 => "11101100",5652 => "00100101",5653 => "10000000",5654 => "10111000",5655 => "00101010",5656 => "10000001",5657 => "10111111",5658 => "00000010",5659 => "11101000",5660 => "10011001",5661 => "01110011",5662 => "11001010",5663 => "10100111",5664 => "11111111",5665 => "10000000",5666 => "00111110",5667 => "11110101",5668 => "10110100",5669 => "00111010",5670 => "11111000",5671 => "10001001",5672 => "10110011",5673 => "10101010",5674 => "01010111",5675 => "10111101",5676 => "00101001",5677 => "11111011",5678 => "01010100",5679 => "11011010",5680 => "10011001",5681 => "10011011",5682 => "00010100",5683 => "00000101",5684 => "10100001",5685 => "01010011",5686 => "11100011",5687 => "01000100",5688 => "01111011",5689 => "01010110",5690 => "01010001",5691 => "11100011",5692 => "00100111",5693 => "01011110",5694 => "01100111",5695 => "11000111",5696 => "00101101",5697 => "01000000",5698 => "10100001",5699 => "00111110",5700 => "01001101",5701 => "01011110",5702 => "00111100",5703 => "10100100",5704 => "01011111",5705 => "00000101",5706 => "10110110",5707 => "00111000",5708 => "00011110",5709 => "10011011",5710 => "10000001",5711 => "00000010",5712 => "10011100",5713 => "00110110",5714 => "11100000",5715 => "11110101",5716 => "00011101",5717 => "11010110",5718 => "00101001",5719 => "10110111",5720 => "11110111",5721 => "10111110",5722 => "00001010",5723 => "00001110",5724 => "01011110",5725 => "10111100",5726 => "01101100",5727 => "00001001",5728 => "00000011",5729 => "11000111",5730 => "11001111",5731 => "00011000",5732 => "01110100",5733 => "11100000",5734 => "10001100",5735 => "11100000",5736 => "00010111",5737 => "10010001",5738 => "01011011",5739 => "01001010",5740 => "01000001",5741 => "11111010",5742 => "01001101",5743 => "01111000",5744 => "11100100",5745 => "11110100",5746 => "10001100",5747 => "01000011",5748 => "01110111",5749 => "10100100",5750 => "10001011",5751 => "01010110",5752 => "10110110",5753 => "01111010",5754 => "11110111",5755 => "10000001",5756 => "10100101",5757 => "10011001",5758 => "11110101",5759 => "10101000",5760 => "00001110",5761 => "11111110",5762 => "11011101",5763 => "11100110",5764 => "01100101",5765 => "10110110",5766 => "00000101",5767 => "10011110",5768 => "00011111",5769 => "10111100",5770 => "00101010",5771 => "01111001",5772 => "01001001",5773 => "00101000",5774 => "00010100",5775 => "10111010",5776 => "01100000",5777 => "01100000",5778 => "10111000",5779 => "00010100",5780 => "11101111",5781 => "11011101",5782 => "00111101",5783 => "01000001",5784 => "11010110",5785 => "00101001",5786 => "11000011",5787 => "01110111",5788 => "00101001",5789 => "10010101",5790 => "01000110",5791 => "00000101",5792 => "00110000",5793 => "11001101",5794 => "11000111",5795 => "01101111",5796 => "10100011",5797 => "00111110",5798 => "11010101",5799 => "10101010",5800 => "01111111",5801 => "11100101",5802 => "00110011",5803 => "11100011",5804 => "00000011",5805 => "00000000",5806 => "01110111",5807 => "01001110",5808 => "01010101",5809 => "01100000",5810 => "01011100",5811 => "00111011",5812 => "11110010",5813 => "10111010",5814 => "01100111",5815 => "10101100",5816 => "01011011",5817 => "01101011",5818 => "11111001",5819 => "00110110",5820 => "00110110",5821 => "11001101",5822 => "01101111",5823 => "00000011",5824 => "11000010",5825 => "11000110",5826 => "11010011",5827 => "11010101",5828 => "10010001",5829 => "01111010",5830 => "01100000",5831 => "01111011",5832 => "01110101",5833 => "10001100",5834 => "10001100",5835 => "10111010",5836 => "10001110",5837 => "01101010",5838 => "00010001",5839 => "00101111",5840 => "00001110",5841 => "01100101",5842 => "11111011",5843 => "10011001",5844 => "11110110",5845 => "11101011",5846 => "11011110",5847 => "00010010",5848 => "11100010",5849 => "00110110",5850 => "01010111",5851 => "01011100",5852 => "11100101",5853 => "10101110",5854 => "00110110",5855 => "00111000",5856 => "00011001",5857 => "01001010",5858 => "11011000",5859 => "10001011",5860 => "10100101",5861 => "11101110",5862 => "11110110",5863 => "01010101",5864 => "11001010",5865 => "00010001",5866 => "11100111",5867 => "01000001",5868 => "11100110",5869 => "01101000",5870 => "00000011",5871 => "00101111",5872 => "00011010",5873 => "10100101",5874 => "11101010",5875 => "10101011",5876 => "10011011",5877 => "10000001",5878 => "11110000",5879 => "01011100",5880 => "10001000",5881 => "10100101",5882 => "00000011",5883 => "11101000",5884 => "11101000",5885 => "11010000",5886 => "01011011",5887 => "01000011",5888 => "10011110",5889 => "00110010",5890 => "11010111",5891 => "11000101",5892 => "00001110",5893 => "10011100",5894 => "11011000",5895 => "10010010",5896 => "00111111",5897 => "00100001",5898 => "01000110",5899 => "11000111",5900 => "01111000",5901 => "11111110",5902 => "10101001",5903 => "10110110",5904 => "00110000",5905 => "11111000",5906 => "00001110",5907 => "00000000",5908 => "11110110",5909 => "10000001",5910 => "00011010",5911 => "01101110",5912 => "11010011",5913 => "11001111",5914 => "00011011",5915 => "10101101",5916 => "01111010",5917 => "01001101",5918 => "01100001",5919 => "00111000",5920 => "00111011",5921 => "01000110",5922 => "10101000",5923 => "01101110",5924 => "01111101",5925 => "10110111",5926 => "10011000",5927 => "11100111",5928 => "00110100",5929 => "10111100",5930 => "00111000",5931 => "01100111",5932 => "00110101",5933 => "11101100",5934 => "00111101",5935 => "10101011",5936 => "10011010",5937 => "10111010",5938 => "01010010",5939 => "01111011",5940 => "01100101",5941 => "11000110",5942 => "00110101",5943 => "01000111",5944 => "01110000",5945 => "00000011",5946 => "00101100",5947 => "10100100",5948 => "10000001",5949 => "00100100",5950 => "00111111",5951 => "00100010",5952 => "11011001",5953 => "01100001",5954 => "10000001",5955 => "01101010",5956 => "10110100",5957 => "11000101",5958 => "01110111",5959 => "11100100",5960 => "00111111",5961 => "10101101",5962 => "10010010",5963 => "01110110",5964 => "11010010",5965 => "01111000",5966 => "00010010",5967 => "10010010",5968 => "10000101",5969 => "11011000",5970 => "10101101",5971 => "00111111",5972 => "11100010",5973 => "10110010",5974 => "10011000",5975 => "10000001",5976 => "00101111",5977 => "01000111",5978 => "11111011",5979 => "11111111",5980 => "01101110",5981 => "00011011",5982 => "00010000",5983 => "01000100",5984 => "00110110",5985 => "10101100",5986 => "11111010",5987 => "10111101",5988 => "11001101",5989 => "10100110",5990 => "11100000",5991 => "01101101",5992 => "01100011",5993 => "10010101",5994 => "01100110",5995 => "00111011",5996 => "00001111",5997 => "01000001",5998 => "11001001",5999 => "01110111",6000 => "11011100",6001 => "00100111",6002 => "00000110",6003 => "11001001",6004 => "11101000",6005 => "01001100",6006 => "10011111",6007 => "10011110",6008 => "11000101",6009 => "11000010",6010 => "00100010",6011 => "10100011",6012 => "00011011",6013 => "10001011",6014 => "10011111",6015 => "00011110",6016 => "10000110",6017 => "00011011",6018 => "11011111",6019 => "10011010",6020 => "11001010",6021 => "01101100",6022 => "01001011",6023 => "11011001",6024 => "01011000",6025 => "00110000",6026 => "10100110",6027 => "00010001",6028 => "10010110",6029 => "10101000",6030 => "11001000",6031 => "11111001",6032 => "11011110",6033 => "10101000",6034 => "11000000",6035 => "10010010",6036 => "11101000",6037 => "11101111",6038 => "10111010",6039 => "11100100",6040 => "00111110",6041 => "10001010",6042 => "11001000",6043 => "10101000",6044 => "11011001",6045 => "11101100",6046 => "00011010",6047 => "00110100",6048 => "11010110",6049 => "00100111",6050 => "01110100",6051 => "01101011",6052 => "01111111",6053 => "10001111",6054 => "11001100",6055 => "01011000",6056 => "11011110",6057 => "10111011",6058 => "01101101",6059 => "11111101",6060 => "00100001",6061 => "00001101",6062 => "11010001",6063 => "10001010",6064 => "01001010",6065 => "01001101",6066 => "11111000",6067 => "10111011",6068 => "11011010",6069 => "10011101",6070 => "00011110",6071 => "01111011",6072 => "11111010",6073 => "01101110",6074 => "01000011",6075 => "11010011",6076 => "00001101",6077 => "00101000",6078 => "10010001",6079 => "11100010",6080 => "00110000",6081 => "11101001",6082 => "00010010",6083 => "01110101",6084 => "00111011",6085 => "10011010",6086 => "01110010",6087 => "01010111",6088 => "10110011",6089 => "10000011",6090 => "00010100",6091 => "10000001",6092 => "01000010",6093 => "01111010",6094 => "11000110",6095 => "11101001",6096 => "11110100",6097 => "11100001",6098 => "00011100",6099 => "11100111",6100 => "00011011",6101 => "01001011",6102 => "11110100",6103 => "00110100",6104 => "00111011",6105 => "11010011",6106 => "00100111",6107 => "00111011",6108 => "11001110",6109 => "10011000",6110 => "00101010",6111 => "00010000",6112 => "00111000",6113 => "11111011",6114 => "10101010",6115 => "11000110",6116 => "11000111",6117 => "11110011",6118 => "01000010",6119 => "10110010",6120 => "10001010",6121 => "00110000",6122 => "11010001",6123 => "01011110",6124 => "10101110",6125 => "11000100",6126 => "11101010",6127 => "11000100",6128 => "01011100",6129 => "00110011",6130 => "01111100",6131 => "10110000",6132 => "01111011",6133 => "10111101",6134 => "00001010",6135 => "00100001",6136 => "10001101",6137 => "00100101",6138 => "11010110",6139 => "01010101",6140 => "01111100",6141 => "11100010",6142 => "10100001",6143 => "00101011",6144 => "11110000",6145 => "10110001",6146 => "01010010",6147 => "11110000",6148 => "10000000",6149 => "11111100",6150 => "01101010",6151 => "11010010",6152 => "01010000",6153 => "00010101",6154 => "10110100",6155 => "00011110",6156 => "01011001",6157 => "11100101",6158 => "01000101",6159 => "01011010",6160 => "10010100",6161 => "00101101",6162 => "00101011",6163 => "11011001",6164 => "10111001",6165 => "10101111",6166 => "10011100",6167 => "01011110",6168 => "10001011",6169 => "01001111",6170 => "10010111",6171 => "01110000",6172 => "00000000",6173 => "00101011",6174 => "10000000",6175 => "00011001",6176 => "01011101",6177 => "00100101",6178 => "11101001",6179 => "00001110",6180 => "11111100",6181 => "11000111",6182 => "00011011",6183 => "10101111",6184 => "00001110",6185 => "00101101",6186 => "11010010",6187 => "00101100",6188 => "10100001",6189 => "10011010",6190 => "00111000",6191 => "01100110",6192 => "00100000",6193 => "11011100",6194 => "01010110",6195 => "01110110",6196 => "01100111",6197 => "10111111",6198 => "10110100",6199 => "11010110",6200 => "10010000",6201 => "01111001",6202 => "11111111",6203 => "10010010",6204 => "00100100",6205 => "01000100",6206 => "11111000",6207 => "01111100",6208 => "00100000",6209 => "10101010",6210 => "11110110",6211 => "00010000",6212 => "10111111",6213 => "10101010",6214 => "10011111",6215 => "00010110",6216 => "00111010",6217 => "01011011",6218 => "11011100",6219 => "10101010",6220 => "11001011",6221 => "11000010",6222 => "00110010",6223 => "11111110",6224 => "10011010",6225 => "00100100",6226 => "00000011",6227 => "01011011",6228 => "10000110",6229 => "01011001",6230 => "01000101",6231 => "00000011",6232 => "10011001",6233 => "00111110",6234 => "01001010",6235 => "01010000",6236 => "01000000",6237 => "00010010",6238 => "10101001",6239 => "11010010",6240 => "00110010",6241 => "11111000",6242 => "01001111",6243 => "11100001",6244 => "11100100",6245 => "10100101",6246 => "00010101",6247 => "00010000",6248 => "10100011",6249 => "10110010",6250 => "10001000",6251 => "11111001",6252 => "10000001",6253 => "00101001",6254 => "01111000",6255 => "01100100",6256 => "10000011",6257 => "11000111",6258 => "00010000",6259 => "10100000",6260 => "01010101",6261 => "00100011",6262 => "00100000",6263 => "01011000",6264 => "10010001",6265 => "11001000",6266 => "10001110",6267 => "00101011",6268 => "11101011",6269 => "10010001",6270 => "00100110",6271 => "10111100",6272 => "00010111",6273 => "10101001",6274 => "01100011",6275 => "10111001",6276 => "11100010",6277 => "00011100",6278 => "01001100",6279 => "00000111",6280 => "00010100",6281 => "00101100",6282 => "10101011",6283 => "01100110",6284 => "10001001",6285 => "11011111",6286 => "00100100",6287 => "01111101",6288 => "11010110",6289 => "11011111",6290 => "10000001",6291 => "10000010",6292 => "01001111",6293 => "00110000",6294 => "11101010",6295 => "10100000",6296 => "01111101",6297 => "00110010",6298 => "10100010",6299 => "01110001",6300 => "00110100",6301 => "11110101",6302 => "01110000",6303 => "01100100",6304 => "11100111",6305 => "00011100",6306 => "11011011",6307 => "11011011",6308 => "11001110",6309 => "11011011",6310 => "10110101",6311 => "00000000",6312 => "11011010",6313 => "10110111",6314 => "10000110",6315 => "11101010",6316 => "11000000",6317 => "11101001",6318 => "00110010",6319 => "11111111",6320 => "11011011",6321 => "00111101",6322 => "01100010",6323 => "01011001",6324 => "01110001",6325 => "11101001",6326 => "00000011",6327 => "00010000",6328 => "00000100",6329 => "10111001",6330 => "00010000",6331 => "01101101",6332 => "01100110",6333 => "11001001",6334 => "10011101",6335 => "01110100",6336 => "00111111",6337 => "11110011",6338 => "01101000",6339 => "00100111",6340 => "00100010",6341 => "11001001",6342 => "11110111",6343 => "01001101",6344 => "01011001",6345 => "01011000",6346 => "01101100",6347 => "10110101",6348 => "00100101",6349 => "00111111",6350 => "01011110",6351 => "01110010",6352 => "11011111",6353 => "11010100",6354 => "11001001",6355 => "10011000",6356 => "00111101",6357 => "01110101",6358 => "10111100",6359 => "01000111",6360 => "10000000",6361 => "10101000",6362 => "10011110",6363 => "10101111",6364 => "01010111",6365 => "00100100",6366 => "11110011",6367 => "11000110",6368 => "01010011",6369 => "01011100",6370 => "00001010",6371 => "11110110",6372 => "01010100",6373 => "11101001",6374 => "00110101",6375 => "10010000",6376 => "10001101",6377 => "01100100",6378 => "10111101",6379 => "01010100",6380 => "01000001",6381 => "11111010",6382 => "11001011",6383 => "10010001",6384 => "11110011",6385 => "10001001",6386 => "11110010",6387 => "10001011",6388 => "10000000",6389 => "00000001",6390 => "10101010",6391 => "11101010",6392 => "00110011",6393 => "01011101",6394 => "00111100",6395 => "11001010",6396 => "11001101",6397 => "10001001",6398 => "00100000",6399 => "11001000",6400 => "10101000",6401 => "10101001",6402 => "10110101",6403 => "10011111",6404 => "00000101",6405 => "11010000",6406 => "01110000",6407 => "01110010",6408 => "10100100",6409 => "10010001",6410 => "11101111",6411 => "11000101",6412 => "01110001",6413 => "01010000",6414 => "01101101",6415 => "11000000",6416 => "11111100",6417 => "01000101",6418 => "10010011",6419 => "00001000",6420 => "00111011",6421 => "01111100",6422 => "11011101",6423 => "11100010",6424 => "01110111",6425 => "00011001",6426 => "01001011",6427 => "11000101",6428 => "01001100",6429 => "01111100",6430 => "10100010",6431 => "11011100",6432 => "11110010",6433 => "10110111",6434 => "11110101",6435 => "10001000",6436 => "10001110",6437 => "10001110",6438 => "01011110",6439 => "10100011",6440 => "10100011",6441 => "10101111",6442 => "01101100",6443 => "01011100",6444 => "11110111",6445 => "10001100",6446 => "01100011",6447 => "11010010",6448 => "11010110",6449 => "01000100",6450 => "00110111",6451 => "10001001",6452 => "00110101",6453 => "00101010",6454 => "11000100",6455 => "10101001",6456 => "10101011",6457 => "10001100",6458 => "00010000",6459 => "00100110",6460 => "01101001",6461 => "01010111",6462 => "00111001",6463 => "00111111",6464 => "10011100",6465 => "00110010",6466 => "11000001",6467 => "01111110",6468 => "10010101",6469 => "00110111",6470 => "11111000",6471 => "01011001",6472 => "00110101",6473 => "00001100",6474 => "11111100",6475 => "11001111",6476 => "00111110",6477 => "01001001",6478 => "01011101",6479 => "11111100",6480 => "11010100",6481 => "00011110",6482 => "01010111",6483 => "11011111",6484 => "01011011",6485 => "10011101",6486 => "10110011",6487 => "01010001",6488 => "10001100",6489 => "11011101",6490 => "10111001",6491 => "00000010",6492 => "11111101",6493 => "00001100",6494 => "11111000",6495 => "11111100",6496 => "01010010",6497 => "11101001",6498 => "00100010",6499 => "01010111",6500 => "11111100",6501 => "01110110",6502 => "10010000",6503 => "00000000",6504 => "11110110",6505 => "01000100",6506 => "01110100",6507 => "10101010",6508 => "00010011",6509 => "10010001",6510 => "11101010",6511 => "01111111",6512 => "10010110",6513 => "01001000",6514 => "11100000",6515 => "11111110",6516 => "10111110",6517 => "00111001",6518 => "01011001",6519 => "01101110",6520 => "11011100",6521 => "01111010",6522 => "01010111",6523 => "00101001",6524 => "01000000",6525 => "11111001",6526 => "10110010",6527 => "10111110",6528 => "00100001",6529 => "11000100",6530 => "01001000",6531 => "00001110",6532 => "10000001",6533 => "10111001",6534 => "01111111",6535 => "00111100",6536 => "00111101",6537 => "10000100",6538 => "11110001",6539 => "10011011",6540 => "01101101",6541 => "01010011",6542 => "11101100",6543 => "11101100",6544 => "11000000",6545 => "00110000",6546 => "10000101",6547 => "11011010",6548 => "01111110",6549 => "11001110",6550 => "11111010",6551 => "11110001",6552 => "00101101",6553 => "10001010",6554 => "10001111",6555 => "10100011",6556 => "11100110",6557 => "10101111",6558 => "00101001",6559 => "00110010",6560 => "00100101",6561 => "11110100",6562 => "10011011",6563 => "01000011",6564 => "00110011",6565 => "11101101",6566 => "01110011",6567 => "01011100",6568 => "00111001",6569 => "01011000",6570 => "01100101",6571 => "01111100",6572 => "11011100",6573 => "01001000",6574 => "10101100",6575 => "01000000",6576 => "00101100",6577 => "00110101",6578 => "01111110",6579 => "11001000",6580 => "00111111",6581 => "01100111",6582 => "11001010",6583 => "01110111",6584 => "11110000",6585 => "01101001",6586 => "01001100",6587 => "11111010",6588 => "11001110",6589 => "01100011",6590 => "01110000",6591 => "10101101",6592 => "10000110",6593 => "11001000",6594 => "01011101",6595 => "01111111",6596 => "10101000",6597 => "10111110",6598 => "01001110",6599 => "00000010",6600 => "11101001",6601 => "10011000",6602 => "11101011",6603 => "11110110",6604 => "11010010",6605 => "11001110",6606 => "00000111",6607 => "00001011",6608 => "10110011",6609 => "00111111",6610 => "00111000",6611 => "00011101",6612 => "00111101",6613 => "00101010",6614 => "00001101",6615 => "01000111",6616 => "01100111",6617 => "01000010",6618 => "00000011",6619 => "00000011",6620 => "00100011",6621 => "10001111",6622 => "00001110",6623 => "01010011",6624 => "11100110",6625 => "01111001",6626 => "10111000",6627 => "00000000",6628 => "10001011",6629 => "11001101",6630 => "11111111",6631 => "10000100",6632 => "10000010",6633 => "00111001",6634 => "00101111",6635 => "10111111",6636 => "01001110",6637 => "01111011",6638 => "01101010",6639 => "01010011",6640 => "10001100",6641 => "10111001",6642 => "10101001",6643 => "00001110",6644 => "00001010",6645 => "01100111",6646 => "10000011",6647 => "01110000",6648 => "11100011",6649 => "00001110",6650 => "10101100",6651 => "00101010",6652 => "10011110",6653 => "11000011",6654 => "00010011",6655 => "01110001",6656 => "10010011",6657 => "01101101",6658 => "00101100",6659 => "10001001",6660 => "11101001",6661 => "01010000",6662 => "11010111",6663 => "11100100",6664 => "10101111",6665 => "11001100",6666 => "00001110",6667 => "00111101",6668 => "01100111",6669 => "11101101",6670 => "11100110",6671 => "10110010",6672 => "10100000",6673 => "11011100",6674 => "10110101",6675 => "11100011",6676 => "10101101",6677 => "00111100",6678 => "11000001",6679 => "10101110",6680 => "01011000",6681 => "11111111",6682 => "11001001",6683 => "00110100",6684 => "11110101",6685 => "11101010",6686 => "10100101",6687 => "11000001",6688 => "00001000",6689 => "01011110",6690 => "00100111",6691 => "01111011",6692 => "01110000",6693 => "10001101",6694 => "01001110",6695 => "10110111",6696 => "01011001",6697 => "10111101",6698 => "00010001",6699 => "11101000",6700 => "00110110",6701 => "00101011",6702 => "01010000",6703 => "00101111",6704 => "11100101",6705 => "11111111",6706 => "11000011",6707 => "10100111",6708 => "10101010",6709 => "10011011",6710 => "01001111",6711 => "11010011",6712 => "00111110",6713 => "00111111",6714 => "10110101",6715 => "11010110",6716 => "10011011",6717 => "00010100",6718 => "01001100",6719 => "11111011",6720 => "01000001",6721 => "00111001",6722 => "11111110",6723 => "10010000",6724 => "10110001",6725 => "10101111",6726 => "11010111",6727 => "10011100",6728 => "00111100",6729 => "00000100",6730 => "01101110",6731 => "00100100",6732 => "10110100",6733 => "00000100",6734 => "10010010",6735 => "11000110",6736 => "01011100",6737 => "01101000",6738 => "01100101",6739 => "10100001",6740 => "10101110",6741 => "00101101",6742 => "11011111",6743 => "00011111",6744 => "10100110",6745 => "11000000",6746 => "10000101",6747 => "10100010",6748 => "01011111",6749 => "11100100",6750 => "10111101",6751 => "01001110",6752 => "11101101",6753 => "01110111",6754 => "11010001",6755 => "00100010",6756 => "11101001",6757 => "10100110",6758 => "10100010",6759 => "11111101",6760 => "00100100",6761 => "01111011",6762 => "10100001",6763 => "10001011",6764 => "10100110",6765 => "00110100",6766 => "00111001",6767 => "11111101",6768 => "10010010",6769 => "01001010",6770 => "11100011",6771 => "11100011",6772 => "11110000",6773 => "11111001",6774 => "11010000",6775 => "11111000",6776 => "00000011",6777 => "00110010",6778 => "00110000",6779 => "01110101",6780 => "11000111",6781 => "01001001",6782 => "11111111",6783 => "01100111",6784 => "10101101",6785 => "11011000",6786 => "10101111",6787 => "10001000",6788 => "11100111",6789 => "00000010",6790 => "10010100",6791 => "00100111",6792 => "01000010",6793 => "00001111",6794 => "00000011",6795 => "11011111",6796 => "11011111",6797 => "11100100",6798 => "10111101",6799 => "01111110",6800 => "10101000",6801 => "01100010",6802 => "10100000",6803 => "01101000",6804 => "10100010",6805 => "01010100",6806 => "00001111",6807 => "11010100",6808 => "11110010",6809 => "11101010",6810 => "01011100",6811 => "00001011",6812 => "01011100",6813 => "00011111",6814 => "11011100",6815 => "00100110",6816 => "01010000",6817 => "00010111",6818 => "01001110",6819 => "00000101",6820 => "01100111",6821 => "11101010",6822 => "00010111",6823 => "01011000",6824 => "01111000",6825 => "01110010",6826 => "01010010",6827 => "01111101",6828 => "10110101",6829 => "01010110",6830 => "11100011",6831 => "00010110",6832 => "00010110",6833 => "01001011",6834 => "10111001",6835 => "01100110",6836 => "00010011",6837 => "11100000",6838 => "00001100",6839 => "01110111",6840 => "11100100",6841 => "10101001",6842 => "10011110",6843 => "10110101",6844 => "00001000",6845 => "10000100",6846 => "11001100",6847 => "11000010",6848 => "01000001",6849 => "01111110",6850 => "01001101",6851 => "00100101",6852 => "00000101",6853 => "11010100",6854 => "11111111",6855 => "11000001",6856 => "00101111",6857 => "00101011",6858 => "00111111",6859 => "01100110",6860 => "11001100",6861 => "00111111",6862 => "00101010",6863 => "11000011",6864 => "01110100",6865 => "00101100",6866 => "01101001",6867 => "11010110",6868 => "01111111",6869 => "01110001",6870 => "01011110",6871 => "00100110",6872 => "00100011",6873 => "10100101",6874 => "01010010",6875 => "11101001",6876 => "10001111",6877 => "00011010",6878 => "01101111",6879 => "01110100",6880 => "11011001",6881 => "10011000",6882 => "01000000",6883 => "00001101",6884 => "00010101",6885 => "10011101",6886 => "10010011",6887 => "10100000",6888 => "10110100",6889 => "01100010",6890 => "00011001",6891 => "00011000",6892 => "00001011",6893 => "10010011",6894 => "01110001",6895 => "10001111",6896 => "10110001",6897 => "10000110",6898 => "10011011",6899 => "01010010",6900 => "01100100",6901 => "00011111",6902 => "11100100",6903 => "00111000",6904 => "01001111",6905 => "10000110",6906 => "10000001",6907 => "11010010",6908 => "11111101",6909 => "11110001",6910 => "10010111",6911 => "01111101",6912 => "10100111",6913 => "01011001",6914 => "01110111",6915 => "10100010",6916 => "11011111",6917 => "11111000",6918 => "00101010",6919 => "10100011",6920 => "10110101",6921 => "10101110",6922 => "10100001",6923 => "01100001",6924 => "00000111",6925 => "01011001",6926 => "10000101",6927 => "00010110",6928 => "00001100",6929 => "00011110",6930 => "11000010",6931 => "00111010",6932 => "01011111",6933 => "01000011",6934 => "10111011",6935 => "00110111",6936 => "11010111",6937 => "01000110",6938 => "10001110",6939 => "11001011",6940 => "10010011",6941 => "00000100",6942 => "01001111",6943 => "01010100",6944 => "00011101",6945 => "01111011",6946 => "10011010",6947 => "10110111",6948 => "11111010",6949 => "10001000",6950 => "10101010",6951 => "00111111",6952 => "10101110",6953 => "11010010",6954 => "11011100",6955 => "11101011",6956 => "11010100",6957 => "00111111",6958 => "00101111",6959 => "10010010",6960 => "01110011",6961 => "10000100",6962 => "00100010",6963 => "01111010",6964 => "10001010",6965 => "00000000",6966 => "10010001",6967 => "01010011",6968 => "10011110",6969 => "01011010",6970 => "00010110",6971 => "10100110",6972 => "11110010",6973 => "10100111",6974 => "01001100",6975 => "10100000",6976 => "00001010",6977 => "01011011",6978 => "10001111",6979 => "01110100",6980 => "11101100",6981 => "10110101",6982 => "00100001",6983 => "01011010",6984 => "10001001",6985 => "01101100",6986 => "01000011",6987 => "10111010",6988 => "11001001",6989 => "01011010",6990 => "01000000",6991 => "00110111",6992 => "00010011",6993 => "01100100",6994 => "01110100",6995 => "11000101",6996 => "11101101",6997 => "11001010",6998 => "01101000",6999 => "01011100",7000 => "01110100",7001 => "10000110",7002 => "10101101",7003 => "00110111",7004 => "10101101",7005 => "10110010",7006 => "11100010",7007 => "10000001",7008 => "11101001",7009 => "11101100",7010 => "11001101",7011 => "10000100",7012 => "10011101",7013 => "11110100",7014 => "11101011",7015 => "11001010",7016 => "00111011",7017 => "11111111",7018 => "10101100",7019 => "11011001",7020 => "00110100",7021 => "01001110",7022 => "10110111",7023 => "10001010",7024 => "10001101",7025 => "10000001",7026 => "01111101",7027 => "00101010",7028 => "00010101",7029 => "00100010",7030 => "10010000",7031 => "10010110",7032 => "00111010",7033 => "10011001",7034 => "00110000",7035 => "11010001",7036 => "00100111",7037 => "10010111",7038 => "11001011",7039 => "00000110",7040 => "10000111",7041 => "10010110",7042 => "11101001",7043 => "00101000",7044 => "01010100",7045 => "11111111",7046 => "00101000",7047 => "11000011",7048 => "01110100",7049 => "01001100",7050 => "01010101",7051 => "11010000",7052 => "11101111",7053 => "11000011",7054 => "01000011",7055 => "10100000",7056 => "01110000",7057 => "00111011",7058 => "00001101",7059 => "00001111",7060 => "01011000",7061 => "11011111",7062 => "00011000",7063 => "00001001",7064 => "01001001",7065 => "01010001",7066 => "00111111",7067 => "00110000",7068 => "11011101",7069 => "01110101",7070 => "01000111",7071 => "11001101",7072 => "10100110",7073 => "01111111",7074 => "11110010",7075 => "10010001",7076 => "00110101",7077 => "11110111",7078 => "01001011",7079 => "11010011",7080 => "00000000",7081 => "10100111",7082 => "00010010",7083 => "00101100",7084 => "10100111",7085 => "11000001",7086 => "11111100",7087 => "01000010",7088 => "00001101",7089 => "00011011",7090 => "10010101",7091 => "01001111",7092 => "00110110",7093 => "11100100",7094 => "01100101",7095 => "01110110",7096 => "01111011",7097 => "10000000",7098 => "01000101",7099 => "11001110",7100 => "00100111",7101 => "00111100",7102 => "11100010",7103 => "00000001",7104 => "10111001",7105 => "00100101",7106 => "00111001",7107 => "01011000",7108 => "11111110",7109 => "10010110",7110 => "01010011",7111 => "00110100",7112 => "01000101",7113 => "01011101",7114 => "11110101",7115 => "11111010",7116 => "01101100",7117 => "10100001",7118 => "10001001",7119 => "10111111",7120 => "11100111",7121 => "10011101",7122 => "01001010",7123 => "11101100",7124 => "10010010",7125 => "00000011",7126 => "11101001",7127 => "10001010",7128 => "11001110",7129 => "11110000",7130 => "10100000",7131 => "11010111",7132 => "00001110",7133 => "00000100",7134 => "00100101",7135 => "10101101",7136 => "11101101",7137 => "10001001",7138 => "11001111",7139 => "10101011",7140 => "00111111",7141 => "11100100",7142 => "11000001",7143 => "10100001",7144 => "11100101",7145 => "00001100",7146 => "10111110",7147 => "11010100",7148 => "11100000",7149 => "00101101",7150 => "10110011",7151 => "01100111",7152 => "01010100",7153 => "11101111",7154 => "00100001",7155 => "00001111",7156 => "00110111",7157 => "10110011",7158 => "01100001",7159 => "11010001",7160 => "00111011",7161 => "01000100",7162 => "00100101",7163 => "11111111",7164 => "00011110",7165 => "01000111",7166 => "10000100",7167 => "11000010",7168 => "11010011",7169 => "00000111",7170 => "01000000",7171 => "01001010",7172 => "10011100",7173 => "10001011",7174 => "11000100",7175 => "11001001",7176 => "00100000",7177 => "01110011",7178 => "11010001",7179 => "01001010",7180 => "11110111",7181 => "11010000",7182 => "00011100",7183 => "11110111",7184 => "00010000",7185 => "01011110",7186 => "00110001",7187 => "00001110",7188 => "11010110",7189 => "00110010",7190 => "01101101",7191 => "11011111",7192 => "01101111",7193 => "00000101",7194 => "10000010",7195 => "11010111",7196 => "10111001",7197 => "01011111",7198 => "01110101",7199 => "00010001",7200 => "11111010",7201 => "11001011",7202 => "00110001",7203 => "01110111",7204 => "00110010",7205 => "00110000",7206 => "11000110",7207 => "00110001",7208 => "11111100",7209 => "10110111",7210 => "01001001",7211 => "01010000",7212 => "01111101",7213 => "00101001",7214 => "01101001",7215 => "11100010",7216 => "10010001",7217 => "01010000",7218 => "01101110",7219 => "00010010",7220 => "00101110",7221 => "11110010",7222 => "00100100",7223 => "01101100",7224 => "11001001",7225 => "01101010",7226 => "11111100",7227 => "11000111",7228 => "10011011",7229 => "00100110",7230 => "10011001",7231 => "00000011",7232 => "10101010",7233 => "00011100",7234 => "11111001",7235 => "11010100",7236 => "01111000",7237 => "10111111",7238 => "10000010",7239 => "11001110",7240 => "01101111",7241 => "10110010",7242 => "00111010",7243 => "10010010",7244 => "01110101",7245 => "01011111",7246 => "00011111",7247 => "10000101",7248 => "10101110",7249 => "01110110",7250 => "01010111",7251 => "10100101",7252 => "00101110",7253 => "10001000",7254 => "00101010",7255 => "11010010",7256 => "10111100",7257 => "11100100",7258 => "00111110",7259 => "01000011",7260 => "01101110",7261 => "10011100",7262 => "11111110",7263 => "11000001",7264 => "01100110",7265 => "00000001",7266 => "00000001",7267 => "11010111",7268 => "00011100",7269 => "11011011",7270 => "01100001",7271 => "00101110",7272 => "11010010",7273 => "11101110",7274 => "10011000",7275 => "10110001",7276 => "00000001",7277 => "01101101",7278 => "00110000",7279 => "11001111",7280 => "11010011",7281 => "11111100",7282 => "00100101",7283 => "00001111",7284 => "00010001",7285 => "01000011",7286 => "01001001",7287 => "10011001",7288 => "01001110",7289 => "01101111",7290 => "11110111",7291 => "00110001",7292 => "10100111",7293 => "10111010",7294 => "00010101",7295 => "00001010",7296 => "01001101",7297 => "00100001",7298 => "10111010",7299 => "11110010",7300 => "01001001",7301 => "01010111",7302 => "11101101",7303 => "10101011",7304 => "00010111",7305 => "00101001",7306 => "11110100",7307 => "00001111",7308 => "01100111",7309 => "11000110",7310 => "10110100",7311 => "01000110",7312 => "10010100",7313 => "00000010",7314 => "00111000",7315 => "11100001",7316 => "01110000",7317 => "11111000",7318 => "01000100",7319 => "00101101",7320 => "11110011",7321 => "11100111",7322 => "01100111",7323 => "11101100",7324 => "01000010",7325 => "11101111",7326 => "01000110",7327 => "10000000",7328 => "10000110",7329 => "00000110",7330 => "01100010",7331 => "11000101",7332 => "00000000",7333 => "00110010",7334 => "00010101",7335 => "01011001",7336 => "11101000",7337 => "11010101",7338 => "00001000",7339 => "10010010",7340 => "01110101",7341 => "01110110",7342 => "01000000",7343 => "00011110",7344 => "11100010",7345 => "01110101",7346 => "01011001",7347 => "01101011",7348 => "11001000",7349 => "00001111",7350 => "01001111",7351 => "00101001",7352 => "11001101",7353 => "11011111",7354 => "10000000",7355 => "01010010",7356 => "01001101",7357 => "00010011",7358 => "11011100",7359 => "11110111",7360 => "01101001",7361 => "00110011",7362 => "11101110",7363 => "00101011",7364 => "10010010",7365 => "00101010",7366 => "01011000",7367 => "00110011",7368 => "10000001",7369 => "00010001",7370 => "11101011",7371 => "01111110",7372 => "10100001",7373 => "11101111",7374 => "10111100",7375 => "01111101",7376 => "01110000",7377 => "00011000",7378 => "01000101",7379 => "01111000",7380 => "10011100",7381 => "00110100",7382 => "10011101",7383 => "11001111",7384 => "10110000",7385 => "11000010",7386 => "01101000",7387 => "01010100",7388 => "00011010",7389 => "11011010",7390 => "10000111",7391 => "01001111",7392 => "00110101",7393 => "01100111",7394 => "11000101",7395 => "01001001",7396 => "00000010",7397 => "10000111",7398 => "01110011",7399 => "11110001",7400 => "10010100",7401 => "10110101",7402 => "11110100",7403 => "10010010",7404 => "01111101",7405 => "11101111",7406 => "11100101",7407 => "10100000",7408 => "01101010",7409 => "00000001",7410 => "10111100",7411 => "01111000",7412 => "01111101",7413 => "11010100",7414 => "01000000",7415 => "11000110",7416 => "10100111",7417 => "01101110",7418 => "00101001",7419 => "00000011",7420 => "10100101",7421 => "10001100",7422 => "01000001",7423 => "00110111",7424 => "11010011",7425 => "00001100",7426 => "11110101",7427 => "11110011",7428 => "10110111",7429 => "10000110",7430 => "01011011",7431 => "00010000",7432 => "11100000",7433 => "10011111",7434 => "01110100",7435 => "11011011",7436 => "11001000",7437 => "10100111",7438 => "10111101",7439 => "11101100",7440 => "10110101",7441 => "10010100",7442 => "11111010",7443 => "11010001",7444 => "01011110",7445 => "01101011",7446 => "10000000",7447 => "01010101",7448 => "00110110",7449 => "00111011",7450 => "01010111",7451 => "10011111",7452 => "10000111",7453 => "10011010",7454 => "00100001",7455 => "10011011",7456 => "00110010",7457 => "11111110",7458 => "10101110",7459 => "10011011",7460 => "00111001",7461 => "11101111",7462 => "10100110",7463 => "10001011",7464 => "01100001",7465 => "01001011",7466 => "11100110",7467 => "01001001",7468 => "11000101",7469 => "10111101",7470 => "01100010",7471 => "11001110",7472 => "10011010",7473 => "00101000",7474 => "10010000",7475 => "01010011",7476 => "11011010",7477 => "00000100",7478 => "10010000",7479 => "11001100",7480 => "00011111",7481 => "00010000",7482 => "10011100",7483 => "10000101",7484 => "01000010",7485 => "10110010",7486 => "01010011",7487 => "00010111",7488 => "10100011",7489 => "10110010",7490 => "11010001",7491 => "00100011",7492 => "11110011",7493 => "11111001",7494 => "00011110",7495 => "11000010",7496 => "10100011",7497 => "01011000",7498 => "11000110",7499 => "11101110",7500 => "00011001",7501 => "01100000",7502 => "01000011",7503 => "00110011",7504 => "11110111",7505 => "01011111",7506 => "10111110",7507 => "01010010",7508 => "11110000",7509 => "00111101",7510 => "01000100",7511 => "11111101",7512 => "11000111",7513 => "00001001",7514 => "10110011",7515 => "11000101",7516 => "01011010",7517 => "01100110",7518 => "11111100",7519 => "01011000",7520 => "01100010",7521 => "01011000",7522 => "00101101",7523 => "00000101",7524 => "11101010",7525 => "10010001",7526 => "00001111",7527 => "00101100",7528 => "00010101",7529 => "00111101",7530 => "00011000",7531 => "11101011",7532 => "01001011",7533 => "01011111",7534 => "00000010",7535 => "11100011",7536 => "10111111",7537 => "01110001",7538 => "10110010",7539 => "11010001",7540 => "00000011",7541 => "11011111",7542 => "10111111",7543 => "10000111",7544 => "10011100",7545 => "10100000",7546 => "11011100",7547 => "01010100",7548 => "11111100",7549 => "00001100",7550 => "11001011",7551 => "11000111",7552 => "01110111",7553 => "10101101",7554 => "01111011",7555 => "00110101",7556 => "10010001",7557 => "00101011",7558 => "10110011",7559 => "00000101",7560 => "11111101",7561 => "01000101",7562 => "10001000",7563 => "01000111",7564 => "01100001",7565 => "01010000",7566 => "10000010",7567 => "00110001",7568 => "11011111",7569 => "11011100",7570 => "10001000",7571 => "00100010",7572 => "01111101",7573 => "01110111",7574 => "10111011",7575 => "00100101",7576 => "00101101",7577 => "11100000",7578 => "11010110",7579 => "11000010",7580 => "00110101",7581 => "00011001",7582 => "10101000",7583 => "00011101",7584 => "00111001",7585 => "00110010",7586 => "01101001",7587 => "10010101",7588 => "00011001",7589 => "11011011",7590 => "00001000",7591 => "11000011",7592 => "10101101",7593 => "11011111",7594 => "01101101",7595 => "00010110",7596 => "10000001",7597 => "01100011",7598 => "00010011",7599 => "01111100",7600 => "00111011",7601 => "10100110",7602 => "11001111",7603 => "11110001",7604 => "01111010",7605 => "00011111",7606 => "00110100",7607 => "10101100",7608 => "00010100",7609 => "11011111",7610 => "10100101",7611 => "01101111",7612 => "11101100",7613 => "01001111",7614 => "00110000",7615 => "01110011",7616 => "10011000",7617 => "00101111",7618 => "00100101",7619 => "11010110",7620 => "11011000",7621 => "11010011",7622 => "01100101",7623 => "01010000",7624 => "10110101",7625 => "10111110",7626 => "01111100",7627 => "00001001",7628 => "00100101",7629 => "01110110",7630 => "01101000",7631 => "11100111",7632 => "01001001",7633 => "11100111",7634 => "10100100",7635 => "01000111",7636 => "11111010",7637 => "01101101",7638 => "11110001",7639 => "11011100",7640 => "10010101",7641 => "10101111",7642 => "11011010",7643 => "01011001",7644 => "10111000",7645 => "10000100",7646 => "10001000",7647 => "11000101",7648 => "11000101",7649 => "01111010",7650 => "10110011",7651 => "01001111",7652 => "10010001",7653 => "10010000",7654 => "01001010",7655 => "00000101",7656 => "00010111",7657 => "11100001",7658 => "01000111",7659 => "01001010",7660 => "00111001",7661 => "11001101",7662 => "11110111",7663 => "01110111",7664 => "01000001",7665 => "11111000",7666 => "11010001",7667 => "01000100",7668 => "10100110",7669 => "01101100",7670 => "11000001",7671 => "11010100",7672 => "01001001",7673 => "11011011",7674 => "00110111",7675 => "11011101",7676 => "10100000",7677 => "10010011",7678 => "00010101",7679 => "11010110",7680 => "01111010",7681 => "00011110",7682 => "01011000",7683 => "00000010",7684 => "11100111",7685 => "11111010",7686 => "10111000",7687 => "10110010",7688 => "10110011",7689 => "01001101",7690 => "00001110",7691 => "00000001",7692 => "00000111",7693 => "00101010",7694 => "10110010",7695 => "11010000",7696 => "01100111",7697 => "11110101",7698 => "11011100",7699 => "00000001",7700 => "01110010",7701 => "10110010",7702 => "10100100",7703 => "11110101",7704 => "10101010",7705 => "01101000",7706 => "00010111",7707 => "10110101",7708 => "10000011",7709 => "00000000",7710 => "01011101",7711 => "00011011",7712 => "00110001",7713 => "00000001",7714 => "01001000",7715 => "01111111",7716 => "11111010",7717 => "10111001",7718 => "00111110",7719 => "01111100",7720 => "11000110",7721 => "10011011",7722 => "01010101",7723 => "00100111",7724 => "01011000",7725 => "00111001",7726 => "10101111",7727 => "11110000",7728 => "00000111",7729 => "10110011",7730 => "00110010",7731 => "10010110",7732 => "10101100",7733 => "11110011",7734 => "01101110",7735 => "11001110",7736 => "11100000",7737 => "01001000",7738 => "00010010",7739 => "10011100",7740 => "11111111",7741 => "11101111",7742 => "00001111",7743 => "00001000",7744 => "00000001",7745 => "00110001",7746 => "11010011",7747 => "00011010",7748 => "00110110",7749 => "11000101",7750 => "11110101",7751 => "11001111",7752 => "11000000",7753 => "01010110",7754 => "01000110",7755 => "00000011",7756 => "01011110",7757 => "00001101",7758 => "10011001",7759 => "01010110",7760 => "00101101",7761 => "10100011",7762 => "10011000",7763 => "01111010",7764 => "10100111",7765 => "00100011",7766 => "01100100",7767 => "01111000",7768 => "10011110",7769 => "01011010",7770 => "00100100",7771 => "01001101",7772 => "11110001",7773 => "10011011",7774 => "00000111",7775 => "01101110",7776 => "10110101",7777 => "00001100",7778 => "10010101",7779 => "01010010",7780 => "00110000",7781 => "11111111",7782 => "10101100",7783 => "01110000",7784 => "01101011",7785 => "01010101",7786 => "01111001",7787 => "00111111",7788 => "01110111",7789 => "00011101",7790 => "01011010",7791 => "00110001",7792 => "10000101",7793 => "11111010",7794 => "10010000",7795 => "01011010",7796 => "00100000",7797 => "00110100",7798 => "00001101",7799 => "11100001",7800 => "01101010",7801 => "00011101",7802 => "00101011",7803 => "10101100",7804 => "10101000",7805 => "10101100",7806 => "00010111",7807 => "10001100",7808 => "11010000",7809 => "00101011",7810 => "01100010",7811 => "01111100",7812 => "10010011",7813 => "11100001",7814 => "01101111",7815 => "00011110",7816 => "00100101",7817 => "11100001",7818 => "00000101",7819 => "10001011",7820 => "10010011",7821 => "10001111",7822 => "11001001",7823 => "01101010",7824 => "00001001",7825 => "00011001",7826 => "11100101",7827 => "01101010",7828 => "11111110",7829 => "11111001",7830 => "10110000",7831 => "11010011",7832 => "01011110",7833 => "01000110",7834 => "11000010",7835 => "10001000",7836 => "00011010",7837 => "00100011",7838 => "00110110",7839 => "01000001",7840 => "11111011",7841 => "11111001",7842 => "11110110",7843 => "10000001",7844 => "00010001",7845 => "10101011",7846 => "01001100",7847 => "11111000",7848 => "10011110",7849 => "00010101",7850 => "01001010",7851 => "00110011",7852 => "01101010",7853 => "00110101",7854 => "10100111",7855 => "01001100",7856 => "01110100",7857 => "01011110",7858 => "10001101",7859 => "00111010",7860 => "01011001",7861 => "11100001",7862 => "00101111",7863 => "01001111",7864 => "01000100",7865 => "10101100",7866 => "01110011",7867 => "01000100",7868 => "10101110",7869 => "00001001",7870 => "10010001",7871 => "11100001",7872 => "10001101",7873 => "10010100",7874 => "11011000",7875 => "11110010",7876 => "01001000",7877 => "10011000",7878 => "01101011",7879 => "11010000",7880 => "00101001",7881 => "00101111",7882 => "01101110",7883 => "10011110",7884 => "11110111",7885 => "01101010",7886 => "00010110",7887 => "11110101",7888 => "11110101",7889 => "01111111",7890 => "10111111",7891 => "10011010",7892 => "00111111",7893 => "01100111",7894 => "10000110",7895 => "01010010",7896 => "11111101",7897 => "01101011",7898 => "11000011",7899 => "00111100",7900 => "01000101",7901 => "00111100",7902 => "00111110",7903 => "01000110",7904 => "01101010",7905 => "01100000",7906 => "00010000",7907 => "00001110",7908 => "11100100",7909 => "10001110",7910 => "01000011",7911 => "11001011",7912 => "11011101",7913 => "11110101",7914 => "11100010",7915 => "11010101",7916 => "11111000",7917 => "00110011",7918 => "01110110",7919 => "00100101",7920 => "01101011",7921 => "01000101",7922 => "01101101",7923 => "10000011",7924 => "01110111",7925 => "10110001",7926 => "00111001",7927 => "11000101",7928 => "00011110",7929 => "10100101",7930 => "00110110",7931 => "10110010",7932 => "01100111",7933 => "10101011",7934 => "11010101",7935 => "11010100",7936 => "01001000",7937 => "11110110",7938 => "01011010",7939 => "10100000",7940 => "11001011",7941 => "00011001",7942 => "01000110",7943 => "11110111",7944 => "01010101",7945 => "00101100",7946 => "01010101",7947 => "01100011",7948 => "00010000",7949 => "11110101",7950 => "11000010",7951 => "10101101",7952 => "11000110",7953 => "01110111",7954 => "11000111",7955 => "00011000",7956 => "00110110",7957 => "00000011",7958 => "01111010",7959 => "10101111",7960 => "11110011",7961 => "00011001",7962 => "10110001",7963 => "01001000",7964 => "00101000",7965 => "11110010",7966 => "11010111",7967 => "10110011",7968 => "00010011",7969 => "01010001",7970 => "00011000",7971 => "11101000",7972 => "01111100",7973 => "10101110",7974 => "10111111",7975 => "01111101",7976 => "11110110",7977 => "01100101",7978 => "10111000",7979 => "11000110",7980 => "01110110",7981 => "00010111",7982 => "10100111",7983 => "01010110",7984 => "00001101",7985 => "01110100",7986 => "11111100",7987 => "10010001",7988 => "10000110",7989 => "10001010",7990 => "11010111",7991 => "11101011",7992 => "11011111",7993 => "01000101",7994 => "01101100",7995 => "01011011",7996 => "01110001",7997 => "11001101",7998 => "10011001",7999 => "11100001",8000 => "10001101",8001 => "10011110",8002 => "10001100",8003 => "10011100",8004 => "11000000",8005 => "00000000",8006 => "00011000",8007 => "00101110",8008 => "11100111",8009 => "01100010",8010 => "01100100",8011 => "00010001",8012 => "00101000",8013 => "00110100",8014 => "00111110",8015 => "01100101",8016 => "01101110",8017 => "01001111",8018 => "10000100",8019 => "10001110",8020 => "10110011",8021 => "10110101",8022 => "00001011",8023 => "00001001",8024 => "00100111",8025 => "10000110",8026 => "01101110",8027 => "10101011",8028 => "10100011",8029 => "11110010",8030 => "10001100",8031 => "00000001",8032 => "01101001",8033 => "01100011",8034 => "10111000",8035 => "01101110",8036 => "10011111",8037 => "11011001",8038 => "00110101",8039 => "10010001",8040 => "10100000",8041 => "00100100",8042 => "11100110",8043 => "10111110",8044 => "01010000",8045 => "11100011",8046 => "00110011",8047 => "11001001",8048 => "11111101",8049 => "11100110",8050 => "10100111",8051 => "01100011",8052 => "01110111",8053 => "01111101",8054 => "10100001",8055 => "00110001",8056 => "00101111",8057 => "00100110",8058 => "10000010",8059 => "10010001",8060 => "10010001",8061 => "01010010",8062 => "11010011",8063 => "11000011",8064 => "00110011",8065 => "01011011",8066 => "11111111",8067 => "00001111",8068 => "01001110",8069 => "00101010",8070 => "00110010",8071 => "01111111",8072 => "00000011",8073 => "11010100",8074 => "01001110",8075 => "01101111",8076 => "01101011",8077 => "10101010",8078 => "00001101",8079 => "00111110",8080 => "00110101",8081 => "00000000",8082 => "01100011",8083 => "01110010",8084 => "00101011",8085 => "11000000",8086 => "01101001",8087 => "10001011",8088 => "11110111",8089 => "00001100",8090 => "11101101",8091 => "10100101",8092 => "01000010",8093 => "10100100",8094 => "11111010",8095 => "11000000",8096 => "10000011",8097 => "00010000",8098 => "10100110",8099 => "11101101",8100 => "11000011",8101 => "01010111",8102 => "00001110",8103 => "01010000",8104 => "11110000",8105 => "10010000",8106 => "10101010",8107 => "00111101",8108 => "01111110",8109 => "10110011",8110 => "01101010",8111 => "00011011",8112 => "00001100",8113 => "00110010",8114 => "11010101",8115 => "01000101",8116 => "00011101",8117 => "00001100",8118 => "00000011",8119 => "00000100",8120 => "00111101",8121 => "11011110",8122 => "10100011",8123 => "10111110",8124 => "01001010",8125 => "11000001",8126 => "10111101",8127 => "10001001",8128 => "10101000",8129 => "10001010",8130 => "00001101",8131 => "00111011",8132 => "11100100",8133 => "00001111",8134 => "01001010",8135 => "11000101",8136 => "11011011",8137 => "01000010",8138 => "01010010",8139 => "11000111",8140 => "10110011",8141 => "01111100",8142 => "11111010",8143 => "10011010",8144 => "01110100",8145 => "01001111",8146 => "10000010",8147 => "00111010",8148 => "01101110",8149 => "10000001",8150 => "00111000",8151 => "10101010",8152 => "11011000",8153 => "11001111",8154 => "01100110",8155 => "11111100",8156 => "00100000",8157 => "11101010",8158 => "01100110",8159 => "00001000",8160 => "11100100",8161 => "01110101",8162 => "11001010",8163 => "10000010",8164 => "11110101",8165 => "01100010",8166 => "10110100",8167 => "11000001",8168 => "00011010",8169 => "01100110",8170 => "10111101",8171 => "10001110",8172 => "01001110",8173 => "00000010",8174 => "11100010",8175 => "11010111",8176 => "10001011",8177 => "10011101",8178 => "00010001",8179 => "00011100",8180 => "01100001",8181 => "01101111",8182 => "10111100",8183 => "01101010",8184 => "01111010",8185 => "10100111",8186 => "01110010",8187 => "00101100",8188 => "11001101",8189 => "01101010",8190 => "11010101",8191 => "10000011",8192 => "01011111",8193 => "01000011",8194 => "00110000",8195 => "11011110",8196 => "00101001",8197 => "00101101",8198 => "11110000",8199 => "00011101",8200 => "00000010",8201 => "10001011",8202 => "11011100",8203 => "10000000",8204 => "00010101",8205 => "10011011",8206 => "11100111",8207 => "00001111",8208 => "11100001",8209 => "00110001",8210 => "11010010",8211 => "11101110",8212 => "01101010",8213 => "11010100",8214 => "01010100",8215 => "10010011",8216 => "01000101",8217 => "01000000",8218 => "10100101",8219 => "11111011",8220 => "01100100",8221 => "10110100",8222 => "10001101",8223 => "00111000",8224 => "11011010",8225 => "11010000",8226 => "01110001",8227 => "00100001",8228 => "00010101",8229 => "11111001",8230 => "01101011",8231 => "01101000",8232 => "00100111",8233 => "11111001",8234 => "10000011",8235 => "11111110",8236 => "10101100",8237 => "10101111",8238 => "11000111",8239 => "00100101",8240 => "00111111",8241 => "10100011",8242 => "10111000",8243 => "11101110",8244 => "11101111",8245 => "10110011",8246 => "11101010",8247 => "01101110",8248 => "00100011",8249 => "10101010",8250 => "11101100",8251 => "00011000",8252 => "11011011",8253 => "00010010",8254 => "01111101",8255 => "11101010",8256 => "01001011",8257 => "10100101",8258 => "10101001",8259 => "01000101",8260 => "01110111",8261 => "01000111",8262 => "00111011",8263 => "01111100",8264 => "11111010",8265 => "11111101",8266 => "01000111",8267 => "11010100",8268 => "11011100",8269 => "00000111",8270 => "11100011",8271 => "00110011",8272 => "10101100",8273 => "10111001",8274 => "10010000",8275 => "10100001",8276 => "00001101",8277 => "11100010",8278 => "01000100",8279 => "10111000",8280 => "01111011",8281 => "00100100",8282 => "00111110",8283 => "00100101",8284 => "00110100",8285 => "01010101",8286 => "00001010",8287 => "11001010",8288 => "01101110",8289 => "11011101",8290 => "00100011",8291 => "00110110",8292 => "00111110",8293 => "10111001",8294 => "10111110",8295 => "11101011",8296 => "01100101",8297 => "10010100",8298 => "00011100",8299 => "10010101",8300 => "01001110",8301 => "01010000",8302 => "11011110",8303 => "00101011",8304 => "11111001",8305 => "11011100",8306 => "11110100",8307 => "01101011",8308 => "00101011",8309 => "00011010",8310 => "11000001",8311 => "00100101",8312 => "00010000",8313 => "00000101",8314 => "11100110",8315 => "10000111",8316 => "01100111",8317 => "01100101",8318 => "01011011",8319 => "11101000",8320 => "00000010",8321 => "10111101",8322 => "11000011",8323 => "00110001",8324 => "00110011",8325 => "00111000",8326 => "10001100",8327 => "01011101",8328 => "00100110",8329 => "00011101",8330 => "10001101",8331 => "00100101",8332 => "00110111",8333 => "01010011",8334 => "10010100",8335 => "11000010",8336 => "11101110",8337 => "11000001",8338 => "11101011",8339 => "11101011",8340 => "10000100",8341 => "10000111",8342 => "11110110",8343 => "00100000",8344 => "11101001",8345 => "10011000",8346 => "00111111",8347 => "11100000",8348 => "01001101",8349 => "11110101",8350 => "11111000",8351 => "11001011",8352 => "01111110",8353 => "01000100",8354 => "10101100",8355 => "00010000",8356 => "01011101",8357 => "10011110",8358 => "10111100",8359 => "10000000",8360 => "00011111",8361 => "01010001",8362 => "00100110",8363 => "11010111",8364 => "00011101",8365 => "00110001",8366 => "11100011",8367 => "00111000",8368 => "10100010",8369 => "10001110",8370 => "00111011",8371 => "01111000",8372 => "00100001",8373 => "10100111",8374 => "00011110",8375 => "11000111",8376 => "10001000",8377 => "01001011",8378 => "10111111",8379 => "00011000",8380 => "00111010",8381 => "01010000",8382 => "00111110",8383 => "10100011",8384 => "10010010",8385 => "00011111",8386 => "10101100",8387 => "00010110",8388 => "11001011",8389 => "00000011",8390 => "00100100",8391 => "11000110",8392 => "10010110",8393 => "01010100",8394 => "00100000",8395 => "00101101",8396 => "11110000",8397 => "01001000",8398 => "01010101",8399 => "11111101",8400 => "01111000",8401 => "01101111",8402 => "11010100",8403 => "01100110",8404 => "00001100",8405 => "11011101",8406 => "10100000",8407 => "10110100",8408 => "11000011",8409 => "10100101",8410 => "00101101",8411 => "10111010",8412 => "00001000",8413 => "10110111",8414 => "00001101",8415 => "01110100",8416 => "11000010",8417 => "00111010",8418 => "01010100",8419 => "11110101",8420 => "01011101",8421 => "00000101",8422 => "11011100",8423 => "11000110",8424 => "01010110",8425 => "11101001",8426 => "01011011",8427 => "01010001",8428 => "10101011",8429 => "11000100",8430 => "00001111",8431 => "11000010",8432 => "00101100",8433 => "01110111",8434 => "00110100",8435 => "00000111",8436 => "11011111",8437 => "10011111",8438 => "11011010",8439 => "10001010",8440 => "00101000",8441 => "10000110",8442 => "11110001",8443 => "01001010",8444 => "01010000",8445 => "00010100",8446 => "00101101",8447 => "01001101",8448 => "10000000",8449 => "00100101",8450 => "11010100",8451 => "01101010",8452 => "01000001",8453 => "10011100",8454 => "11110001",8455 => "01101000",8456 => "10011101",8457 => "00011100",8458 => "10000110",8459 => "10101011",8460 => "01100110",8461 => "01110101",8462 => "01100001",8463 => "11110101",8464 => "10110100",8465 => "10110001",8466 => "11010111",8467 => "00100001",8468 => "00011110",8469 => "11000110",8470 => "01110001",8471 => "10010110",8472 => "11111010",8473 => "01000110",8474 => "11110010",8475 => "00111110",8476 => "10011010",8477 => "00001001",8478 => "11001100",8479 => "01100000",8480 => "10100000",8481 => "00000000",8482 => "00010010",8483 => "11011100",8484 => "00111000",8485 => "11110010",8486 => "10110001",8487 => "00011011",8488 => "10100110",8489 => "00110101",8490 => "10111011",8491 => "11010000",8492 => "01011100",8493 => "10110100",8494 => "01110101",8495 => "10011111",8496 => "00101010",8497 => "01011011",8498 => "11100101",8499 => "11100011",8500 => "01000011",8501 => "00100010",8502 => "00001011",8503 => "01010101",8504 => "10010011",8505 => "10111110",8506 => "00101101",8507 => "00001101",8508 => "00011001",8509 => "11100001",8510 => "00001010",8511 => "01011111",8512 => "11111001",8513 => "10111011",8514 => "00011011",8515 => "11010111",8516 => "00100111",8517 => "11110000",8518 => "10011000",8519 => "10000011",8520 => "11110001",8521 => "00111111",8522 => "01000011",8523 => "00101110",8524 => "11100011",8525 => "10110100",8526 => "10110011",8527 => "11111100",8528 => "01001110",8529 => "01111000",8530 => "01100001",8531 => "10101010",8532 => "11111111",8533 => "00111011",8534 => "01100111",8535 => "01101111",8536 => "01011010",8537 => "01001001",8538 => "01001100",8539 => "10111101",8540 => "10001110",8541 => "01101100",8542 => "01101100",8543 => "11110100",8544 => "00011100",8545 => "10111011",8546 => "01100100",8547 => "11100000",8548 => "00110111",8549 => "00010101",8550 => "00100000",8551 => "11011111",8552 => "11100110",8553 => "11010000",8554 => "01010001",8555 => "11000001",8556 => "01111010",8557 => "11110010",8558 => "10110101",8559 => "01100000",8560 => "00010000",8561 => "10101110",8562 => "10101000",8563 => "11111111",8564 => "01000100",8565 => "01100111",8566 => "00101111",8567 => "11010000",8568 => "10001100",8569 => "10011100",8570 => "01001010",8571 => "00010100",8572 => "00110111",8573 => "01110110",8574 => "11000100",8575 => "10101111",8576 => "00100011",8577 => "11011011",8578 => "10000010",8579 => "11111001",8580 => "11101100",8581 => "10110011",8582 => "11011110",8583 => "00000001",8584 => "01100100",8585 => "11010011",8586 => "10111000",8587 => "10010010",8588 => "00111100",8589 => "00000011",8590 => "00011010",8591 => "11110111",8592 => "11011111",8593 => "00000100",8594 => "00010011",8595 => "01000011",8596 => "00010010",8597 => "10001111",8598 => "00101101",8599 => "01111111",8600 => "00111110",8601 => "10000000",8602 => "00010110",8603 => "00110101",8604 => "10100001",8605 => "01101111",8606 => "00110010",8607 => "10111100",8608 => "00000110",8609 => "11001100",8610 => "01010001",8611 => "00011000",8612 => "00111011",8613 => "00010011",8614 => "01000010",8615 => "01000011",8616 => "00101010",8617 => "01101011",8618 => "00111110",8619 => "01000001",8620 => "00100000",8621 => "00001101",8622 => "00011101",8623 => "11001111",8624 => "01001111",8625 => "10111111",8626 => "01011010",8627 => "11010110",8628 => "11100010",8629 => "10100110",8630 => "00001110",8631 => "11110001",8632 => "01010011",8633 => "11010001",8634 => "10100000",8635 => "00100011",8636 => "01000001",8637 => "11010010",8638 => "10101101",8639 => "11000000",8640 => "11001001",8641 => "11001100",8642 => "10000000",8643 => "01011101",8644 => "11101001",8645 => "11110001",8646 => "11110100",8647 => "10101011",8648 => "00011001",8649 => "10101001",8650 => "01111101",8651 => "00110110",8652 => "01001100",8653 => "11011100",8654 => "00000111",8655 => "11001011",8656 => "00001001",8657 => "10110110",8658 => "00010101",8659 => "01110011",8660 => "01001011",8661 => "01100110",8662 => "11010010",8663 => "10001011",8664 => "10010000",8665 => "10100011",8666 => "00111001",8667 => "01010000",8668 => "00101101",8669 => "10010001",8670 => "00010101",8671 => "10101010",8672 => "01111100",8673 => "10110010",8674 => "11100001",8675 => "11011101",8676 => "00011000",8677 => "00111101",8678 => "01110100",8679 => "01100110",8680 => "11001001",8681 => "10110010",8682 => "10000001",8683 => "10100001",8684 => "10111111",8685 => "11101111",8686 => "01001001",8687 => "11110010",8688 => "00001111",8689 => "01011110",8690 => "00010110",8691 => "00001010",8692 => "10000101",8693 => "01110000",8694 => "01101111",8695 => "10010100",8696 => "11010111",8697 => "01100110",8698 => "10111101",8699 => "10110101",8700 => "10110000",8701 => "01111010",8702 => "01100110",8703 => "01100011",8704 => "01100011",8705 => "11110011",8706 => "01000100",8707 => "01100110",8708 => "10101011",8709 => "11110110",8710 => "00111001",8711 => "11010011",8712 => "00010001",8713 => "11111100",8714 => "10110111",8715 => "10011001",8716 => "00111001",8717 => "00110011",8718 => "01111101",8719 => "11110000",8720 => "10110001",8721 => "10010100",8722 => "11001010",8723 => "11010011",8724 => "10001010",8725 => "10111111",8726 => "11000111",8727 => "00011011",8728 => "01000101",8729 => "00100000",8730 => "01010111",8731 => "00010001",8732 => "11110100",8733 => "00111000",8734 => "01000010",8735 => "11111011",8736 => "01001000",8737 => "11001000",8738 => "01010110",8739 => "11010111",8740 => "01101001",8741 => "01001010",8742 => "11100111",8743 => "00111101",8744 => "01100011",8745 => "10001100",8746 => "10010110",8747 => "01000110",8748 => "11010001",8749 => "01000000",8750 => "10111001",8751 => "00011000",8752 => "01001110",8753 => "11000011",8754 => "00001110",8755 => "01001000",8756 => "00000011",8757 => "00001110",8758 => "01010000",8759 => "11110010",8760 => "01000111",8761 => "00001010",8762 => "01101000",8763 => "00110101",8764 => "11110110",8765 => "10100111",8766 => "10110001",8767 => "11000111",8768 => "10101011",8769 => "00100100",8770 => "00010101",8771 => "01000011",8772 => "11100001",8773 => "01010011",8774 => "00001110",8775 => "10011010",8776 => "11100001",8777 => "11000010",8778 => "11001001",8779 => "10001100",8780 => "01111110",8781 => "11111110",8782 => "11001100",8783 => "01100101",8784 => "10011100",8785 => "10000000",8786 => "01000100",8787 => "00110011",8788 => "01101101",8789 => "10111110",8790 => "11100111",8791 => "01101010",8792 => "01010101",8793 => "11010000",8794 => "00011001",8795 => "10111010",8796 => "11010100",8797 => "00111110",8798 => "10100011",8799 => "10011001",8800 => "00000110",8801 => "11100110",8802 => "01111011",8803 => "11110101",8804 => "01010101",8805 => "11011010",8806 => "11100110",8807 => "11111110",8808 => "10111001",8809 => "01100110",8810 => "01110101",8811 => "00100010",8812 => "11110010",8813 => "01110010",8814 => "01101111",8815 => "10101111",8816 => "10111111",8817 => "01010000",8818 => "11111010",8819 => "00100100",8820 => "01011111",8821 => "11101001",8822 => "01001001",8823 => "00001101",8824 => "11100010",8825 => "10100100",8826 => "11011000",8827 => "00000011",8828 => "10000101",8829 => "10110010",8830 => "11111000",8831 => "10011001",8832 => "11100100",8833 => "11111011",8834 => "01111100",8835 => "01011001",8836 => "11001101",8837 => "01110011",8838 => "10101000",8839 => "10101111",8840 => "10010011",8841 => "00111001",8842 => "11011010",8843 => "00000100",8844 => "01101100",8845 => "00010101",8846 => "11000110",8847 => "01000101",8848 => "10001000",8849 => "10100000",8850 => "10111101",8851 => "00111101",8852 => "01011100",8853 => "11010001",8854 => "10111010",8855 => "11001101",8856 => "01111101",8857 => "11100001",8858 => "11100110",8859 => "01100011",8860 => "01100001",8861 => "01111011",8862 => "00010011",8863 => "11011000",8864 => "11000000",8865 => "10010001",8866 => "00000110",8867 => "00111111",8868 => "00101100",8869 => "00000011",8870 => "10110011",8871 => "10011100",8872 => "10011000",8873 => "10110001",8874 => "10100111",8875 => "00000000",8876 => "11110101",8877 => "11010111",8878 => "11010100",8879 => "00001111",8880 => "01011000",8881 => "10011011",8882 => "11100111",8883 => "00010010",8884 => "00010000",8885 => "10111110",8886 => "00100101",8887 => "00011100",8888 => "01010111",8889 => "11010101",8890 => "11111011",8891 => "00010010",8892 => "01101111",8893 => "10000111",8894 => "01000011",8895 => "01011111",8896 => "10111011",8897 => "01101101",8898 => "11100001",8899 => "11011011",8900 => "01101001",8901 => "00001111",8902 => "11110110",8903 => "01000101",8904 => "10101100",8905 => "00110111",8906 => "11001101",8907 => "01000110",8908 => "11010111",8909 => "11110001",8910 => "01100011",8911 => "10010011",8912 => "10100101",8913 => "10011100",8914 => "10011111",8915 => "01101011",8916 => "00101100",8917 => "01110001",8918 => "01010100",8919 => "01100101",8920 => "10000100",8921 => "11011110",8922 => "11000100",8923 => "11100001",8924 => "00100111",8925 => "10111000",8926 => "10100011",8927 => "00001010",8928 => "00111000",8929 => "10000100",8930 => "11100110",8931 => "11100100",8932 => "00011101",8933 => "00011011",8934 => "11010100",8935 => "01110000",8936 => "01011101",8937 => "00111010",8938 => "11110100",8939 => "10000100",8940 => "10110110",8941 => "01110011",8942 => "00101001",8943 => "11100010",8944 => "11100100",8945 => "01010100",8946 => "10101000",8947 => "01001011",8948 => "11011010",8949 => "11110100",8950 => "01000111",8951 => "00000101",8952 => "11011000",8953 => "10111111",8954 => "01101011",8955 => "00001001",8956 => "00111010",8957 => "00110101",8958 => "10000001",8959 => "01101111",8960 => "10010011",8961 => "00000101",8962 => "00110000",8963 => "10010110",8964 => "01101111",8965 => "00001011",8966 => "11100101",8967 => "10001000",8968 => "10000011",8969 => "10110101",8970 => "00110000",8971 => "01100011",8972 => "00100010",8973 => "00110011",8974 => "11111001",8975 => "00010111",8976 => "01011101",8977 => "01011011",8978 => "11001101",8979 => "10101111",8980 => "00011010",8981 => "11011110",8982 => "00111001",8983 => "11111000",8984 => "11000111",8985 => "00110110",8986 => "11111011",8987 => "10001101",8988 => "11101001",8989 => "10011101",8990 => "11000010",8991 => "11111110",8992 => "11000110",8993 => "01101110",8994 => "01001000",8995 => "00011000",8996 => "10000011",8997 => "11111000",8998 => "11110111",8999 => "11101111",9000 => "00000101",9001 => "10100110",9002 => "11101111",9003 => "00000010",9004 => "00111011",9005 => "01011101",9006 => "01011101",9007 => "10111101",9008 => "01010000",9009 => "00010010",9010 => "10000000",9011 => "00111100",9012 => "10100101",9013 => "00011011",9014 => "01010101",9015 => "01011101",9016 => "10100001",9017 => "00111111",9018 => "00101000",9019 => "11101101",9020 => "01111010",9021 => "11100101",9022 => "11011010",9023 => "11110100",9024 => "11001011",9025 => "00000111",9026 => "10000001",9027 => "10001001",9028 => "01110101",9029 => "01100101",9030 => "01111011",9031 => "10000110",9032 => "01101111",9033 => "10000110",9034 => "00000001",9035 => "01101010",9036 => "00011010",9037 => "11110100",9038 => "11011101",9039 => "10101010",9040 => "01000101",9041 => "10011111",9042 => "00101101",9043 => "11010111",9044 => "10010110",9045 => "11111011",9046 => "10011101",9047 => "10111101",9048 => "10111010",9049 => "01111011",9050 => "10011111",9051 => "10100001",9052 => "01110101",9053 => "01010100",9054 => "10111001",9055 => "10011000",9056 => "00100100",9057 => "10110110",9058 => "01101110",9059 => "00110111",9060 => "11010101",9061 => "00011000",9062 => "01001110",9063 => "01110110",9064 => "01000011",9065 => "01110111",9066 => "00101000",9067 => "10100111",9068 => "11011010",9069 => "01011111",9070 => "10111101",9071 => "10011000",9072 => "00001101",9073 => "10010011",9074 => "00011010",9075 => "01100000",9076 => "10100011",9077 => "11111101",9078 => "00000000",9079 => "10011110",9080 => "11001011",9081 => "10010000",9082 => "10001101",9083 => "11001000",9084 => "11011101",9085 => "10010011",9086 => "11010010",9087 => "01001100",9088 => "00110000",9089 => "11101100",9090 => "01110101",9091 => "00110100",9092 => "00101001",9093 => "10100000",9094 => "11100011",9095 => "00111100",9096 => "01010010",9097 => "01101000",9098 => "10100101",9099 => "01110111",9100 => "10110010",9101 => "11011011",9102 => "01011100",9103 => "11010110",9104 => "01010011",9105 => "00110101",9106 => "11101011",9107 => "10010011",9108 => "00100001",9109 => "00110110",9110 => "01100110",9111 => "00101000",9112 => "10000011",9113 => "11011000",9114 => "11001000",9115 => "00110101",9116 => "10110110",9117 => "11001000",9118 => "00010001",9119 => "11010111",9120 => "00100100",9121 => "01111000",9122 => "11100010",9123 => "00110000",9124 => "11001011",9125 => "01101100",9126 => "00110000",9127 => "00001011",9128 => "00010101",9129 => "11011111",9130 => "00010101",9131 => "00000110",9132 => "00001101",9133 => "11111111",9134 => "10111100",9135 => "00110110",9136 => "01111001",9137 => "01110000",9138 => "11001100",9139 => "11100100",9140 => "11101111",9141 => "00110001",9142 => "11010101",9143 => "10111110",9144 => "00000101",9145 => "11110101",9146 => "10000111",9147 => "01111110",9148 => "11001100",9149 => "00100011",9150 => "11000000",9151 => "00011111",9152 => "10000010",9153 => "00000111",9154 => "11000110",9155 => "01000010",9156 => "11001111",9157 => "10000100",9158 => "00011010",9159 => "10001010",9160 => "11000101",9161 => "10110001",9162 => "10111010",9163 => "00100111",9164 => "01100111",9165 => "11111110",9166 => "00011010",9167 => "10001001",9168 => "10000011",9169 => "01101111",9170 => "01011101",9171 => "01110001",9172 => "11010100",9173 => "10001011",9174 => "10010000",9175 => "11011001",9176 => "01111111",9177 => "11011001",9178 => "01010111",9179 => "01111100",9180 => "11000001",9181 => "01101010",9182 => "11110000",9183 => "10001100",9184 => "11000101",9185 => "10111001",9186 => "01001110",9187 => "10011000",9188 => "01111111",9189 => "11100010",9190 => "01101001",9191 => "01101101",9192 => "11100011",9193 => "11000111",9194 => "10010010",9195 => "10010000",9196 => "01101011",9197 => "00011111",9198 => "10001111",9199 => "11110110",9200 => "00000010",9201 => "10110001",9202 => "00010100",9203 => "11001011",9204 => "10101101",9205 => "00000001",9206 => "10100000",9207 => "01000001",9208 => "11101011",9209 => "01000011",9210 => "00000111",9211 => "10101101",9212 => "00010100",9213 => "10001001",9214 => "00000001",9215 => "01010101",9216 => "10110011",9217 => "10000000",9218 => "10101010",9219 => "00111111",9220 => "10011110",9221 => "10100110",9222 => "10000110",9223 => "00111101",9224 => "00100000",9225 => "01100100",9226 => "10111010",9227 => "10111110",9228 => "10011111",9229 => "10110111",9230 => "01011011",9231 => "00111100",9232 => "00000101",9233 => "11000110",9234 => "01001101",9235 => "01011101",9236 => "01110011",9237 => "10101010",9238 => "11011010",9239 => "11011011",9240 => "00110101",9241 => "00011001",9242 => "01101110",9243 => "01111011",9244 => "00011000",9245 => "11111110",9246 => "00111000",9247 => "00110010",9248 => "00111111",9249 => "10100100",9250 => "10111010",9251 => "00011110",9252 => "10100111",9253 => "00000000",9254 => "01011101",9255 => "11100101",9256 => "01010010",9257 => "10101000",9258 => "01111101",9259 => "11111000",9260 => "01101011",9261 => "00000010",9262 => "10010100",9263 => "01000100",9264 => "01100110",9265 => "01011100",9266 => "10110111",9267 => "10110011",9268 => "01011011",9269 => "00010100",9270 => "01100100",9271 => "01111100",9272 => "11101000",9273 => "11110110",9274 => "00010110",9275 => "00000010",9276 => "11001111",9277 => "00000110",9278 => "01010100",9279 => "10101101",9280 => "10100011",9281 => "10011001",9282 => "01101011",9283 => "01000111",9284 => "01000000",9285 => "10111001",9286 => "11000011",9287 => "01001011",9288 => "01011010",9289 => "01110000",9290 => "00101011",9291 => "10101001",9292 => "00010000",9293 => "10000111",9294 => "00010001",9295 => "11000111",9296 => "10000010",9297 => "01010011",9298 => "10110100",9299 => "00111000",9300 => "00000010",9301 => "00111000",9302 => "00100100",9303 => "11101110",9304 => "01000001",9305 => "01110101",9306 => "00101001",9307 => "11010101",9308 => "10111111",9309 => "00001011",9310 => "00111101",9311 => "01101001",9312 => "10110111",9313 => "11100100",9314 => "11110010",9315 => "10011010",9316 => "01110011",9317 => "10111100",9318 => "10000111",9319 => "00010000",9320 => "11110010",9321 => "00010100",9322 => "00011011",9323 => "10011010",9324 => "10110111",9325 => "11011001",9326 => "11100101",9327 => "00011011",9328 => "01100011",9329 => "00101000",9330 => "11011011",9331 => "01110101",9332 => "11111001",9333 => "10011000",9334 => "10110000",9335 => "10001000",9336 => "11010110",9337 => "00000011",9338 => "01010000",9339 => "01001001",9340 => "00111000",9341 => "00011000",9342 => "11000111",9343 => "01100011",9344 => "10000110",9345 => "11111101",9346 => "01011010",9347 => "10110001",9348 => "00000011",9349 => "01000001",9350 => "01000000",9351 => "01010100",9352 => "00110010",9353 => "10110010",9354 => "10111111",9355 => "11000011",9356 => "01011101",9357 => "00111000",9358 => "00000011",9359 => "10000010",9360 => "01100100",9361 => "11100100",9362 => "01010011",9363 => "10101100",9364 => "11101001",9365 => "01100100",9366 => "11011001",9367 => "00001001",9368 => "01100001",9369 => "11101001",9370 => "10111001",9371 => "00100110",9372 => "00110100",9373 => "00001000",9374 => "10101001",9375 => "10000110",9376 => "00000101",9377 => "00000100",9378 => "01101100",9379 => "00001101",9380 => "11011000",9381 => "01000100",9382 => "11000100",9383 => "01101000",9384 => "10011010",9385 => "01111000",9386 => "10000001",9387 => "01101011",9388 => "11101000",9389 => "00101011",9390 => "10010101",9391 => "10110111",9392 => "11010001",9393 => "01100001",9394 => "01001101",9395 => "00110110",9396 => "00111101",9397 => "11110101",9398 => "00000010",9399 => "10100001",9400 => "01110111",9401 => "00101110",9402 => "11001110",9403 => "01110110",9404 => "11010110",9405 => "11010000",9406 => "10111000",9407 => "11001111",9408 => "11001001",9409 => "11101001",9410 => "11111011",9411 => "01110011",9412 => "01010011",9413 => "01101111",9414 => "01010011",9415 => "00101000",9416 => "11010111",9417 => "11001010",9418 => "10100110",9419 => "10001000",9420 => "10000101",9421 => "01010001",9422 => "11011000",9423 => "00101000",9424 => "11110011",9425 => "10101110",9426 => "10100110",9427 => "10111000",9428 => "00110111",9429 => "01001111",9430 => "00111000",9431 => "01100100",9432 => "10110001",9433 => "01010010",9434 => "01010001",9435 => "01111101",9436 => "00010000",9437 => "01111000",9438 => "01111011",9439 => "01010000",9440 => "10101110",9441 => "10001101",9442 => "00100111",9443 => "11100000",9444 => "11000010",9445 => "11110110",9446 => "11110000",9447 => "11000110",9448 => "11000111",9449 => "01000010",9450 => "10100100",9451 => "00001111",9452 => "10110100",9453 => "10011101",9454 => "11010110",9455 => "11011000",9456 => "00000100",9457 => "01100100",9458 => "10100011",9459 => "11100000",9460 => "10001011",9461 => "01011110",9462 => "11101111",9463 => "01011011",9464 => "11011111",9465 => "01001100",9466 => "01100100",9467 => "01111001",9468 => "01000010",9469 => "00011111",9470 => "10011111",9471 => "01110111",9472 => "11111011",9473 => "00110111",9474 => "00011110",9475 => "11001111",9476 => "11000110",9477 => "00011000",9478 => "11000111",9479 => "00100001",9480 => "11000111",9481 => "00010101",9482 => "00000111",9483 => "01010001",9484 => "01110111",9485 => "00000000",9486 => "01100101",9487 => "10111001",9488 => "01000010",9489 => "01111101",9490 => "00011000",9491 => "11010110",9492 => "01000001",9493 => "11001100",9494 => "00000001",9495 => "11111111",9496 => "10001010",9497 => "00000010",9498 => "11101101",9499 => "01011000",9500 => "00001011",9501 => "00110101",9502 => "10010001",9503 => "01001100",9504 => "10101011",9505 => "00111101",9506 => "11010110",9507 => "01010101",9508 => "00100101",9509 => "00000001",9510 => "10001100",9511 => "10000011",9512 => "01110010",9513 => "01010100",9514 => "11110000",9515 => "01110110",9516 => "10101100",9517 => "10110101",9518 => "11011010",9519 => "11001101",9520 => "01011011",9521 => "01010101",9522 => "11100001",9523 => "10000011",9524 => "10110111",9525 => "00011010",9526 => "00011111",9527 => "10010000",9528 => "00111111",9529 => "10110100",9530 => "01011101",9531 => "01010110",9532 => "10101101",9533 => "10010111",9534 => "01111001",9535 => "01111011",9536 => "00100101",9537 => "01100010",9538 => "01000010",9539 => "01001110",9540 => "01011001",9541 => "11010100",9542 => "01111010",9543 => "00011000",9544 => "01111010",9545 => "10001011",9546 => "11111001",9547 => "01111101",9548 => "11111010",9549 => "01010110",9550 => "00010111",9551 => "00001100",9552 => "11000000",9553 => "11000100",9554 => "01111100",9555 => "11000001",9556 => "10100110",9557 => "10100111",9558 => "00110001",9559 => "00001110",9560 => "11001001",9561 => "10101101",9562 => "00110111",9563 => "10000010",9564 => "10111111",9565 => "10100110",9566 => "00010100",9567 => "01001100",9568 => "00001010",9569 => "10000000",9570 => "10110010",9571 => "10001000",9572 => "01010000",9573 => "00111110",9574 => "11011101",9575 => "10110010",9576 => "11001001",9577 => "10100110",9578 => "01001001",9579 => "11001100",9580 => "10100100",9581 => "11100111",9582 => "10111111",9583 => "01001010",9584 => "01001100",9585 => "01011111",9586 => "10100101",9587 => "00011100",9588 => "11001011",9589 => "01111110",9590 => "01111001",9591 => "00110111",9592 => "01100111",9593 => "01001001",9594 => "10000110",9595 => "10000100",9596 => "00011001",9597 => "11110000",9598 => "01111010",9599 => "00000110",9600 => "00000111",9601 => "10000000",9602 => "10101011",9603 => "11110110",9604 => "00100011",9605 => "01110110",9606 => "10000010",9607 => "00000010",9608 => "11101011",9609 => "11110000",9610 => "11010111",9611 => "01001001",9612 => "10000100",9613 => "11011010",9614 => "00001010",9615 => "01110101",9616 => "00000101",9617 => "10000000",9618 => "10111000",9619 => "11011110",9620 => "10100110",9621 => "10010110",9622 => "00011010",9623 => "10010100",9624 => "10000001",9625 => "01001010",9626 => "00011111",9627 => "01010011",9628 => "10011000",9629 => "10000101",9630 => "01001000",9631 => "00001100",9632 => "00111011",9633 => "10000010",9634 => "01000001",9635 => "00111111",9636 => "10101100",9637 => "10000100",9638 => "00010011",9639 => "00110001",9640 => "11110101",9641 => "01011001",9642 => "01000011",9643 => "11010011",9644 => "00100000",9645 => "10111100",9646 => "11011100",9647 => "01000101",9648 => "11010000",9649 => "10001011",9650 => "11001000",9651 => "01001011",9652 => "10010010",9653 => "11110000",9654 => "01000000",9655 => "01010100",9656 => "10111110",9657 => "11011101",9658 => "01001000",9659 => "11100111",9660 => "00010110",9661 => "11000110",9662 => "10110000",9663 => "00011011",9664 => "10111101",9665 => "11100000",9666 => "11011000",9667 => "00111010",9668 => "10010111",9669 => "10001000",9670 => "10100100",9671 => "00111101",9672 => "10101010",9673 => "10011010",9674 => "01111101",9675 => "01110100",9676 => "11001000",9677 => "11110101",9678 => "01010100",9679 => "10111111",9680 => "11110110",9681 => "11110001",9682 => "11110100",9683 => "10010011",9684 => "00001111",9685 => "10010010",9686 => "10000001",9687 => "00101011",9688 => "01001100",9689 => "01110101",9690 => "11110100",9691 => "11000000",9692 => "11001110",9693 => "00001100",9694 => "00001011",9695 => "00110011",9696 => "10001001",9697 => "10000001",9698 => "00110100",9699 => "00010110",9700 => "00100010",9701 => "01101010",9702 => "01110000",9703 => "11011110",9704 => "01001011",9705 => "11100111",9706 => "10010001",9707 => "01100001",9708 => "01111011",9709 => "00100001",9710 => "11000110",9711 => "11110100",9712 => "01001111",9713 => "11010110",9714 => "11001000",9715 => "10010010",9716 => "11101000",9717 => "01111011",9718 => "00011100",9719 => "11111000",9720 => "11001110",9721 => "11011111",9722 => "10000100",9723 => "01011000",9724 => "00001101",9725 => "11001111",9726 => "10100111",9727 => "11001011",9728 => "11110000",9729 => "01100110",9730 => "10100001",9731 => "01111001",9732 => "01000111",9733 => "00111010",9734 => "01101101",9735 => "00110101",9736 => "00110110",9737 => "01011010",9738 => "01101110",9739 => "01100100",9740 => "10010011",9741 => "00111000",9742 => "11010110",9743 => "01000000",9744 => "11111000",9745 => "11100010",9746 => "01101110",9747 => "01110110",9748 => "00010100",9749 => "11011111",9750 => "00100001",9751 => "11010001",9752 => "10111011",9753 => "11101111",9754 => "00100101",9755 => "11010100",9756 => "10000011",9757 => "01011111",9758 => "01011110",9759 => "11001100",9760 => "00011100",9761 => "01100010",9762 => "10000011",9763 => "01100000",9764 => "10000111",9765 => "01010100",9766 => "00110110",9767 => "00011010",9768 => "00010011",9769 => "11011101",9770 => "00000001",9771 => "11100010",9772 => "10101001",9773 => "00111000",9774 => "01000001",9775 => "01100110",9776 => "00110111",9777 => "01101101",9778 => "01001011",9779 => "11010010",9780 => "10010111",9781 => "01000010",9782 => "01100001",9783 => "11011011",9784 => "01001000",9785 => "11111000",9786 => "10001110",9787 => "01011111",9788 => "01001010",9789 => "11001001",9790 => "01100110",9791 => "00111110",9792 => "01110010",9793 => "10111001",9794 => "10000001",9795 => "11011011",9796 => "01100000",9797 => "10000010",9798 => "11000110",9799 => "01011000",9800 => "00110000",9801 => "00100001",9802 => "00111010",9803 => "11001010",9804 => "11111000",9805 => "01000011",9806 => "00100001",9807 => "10010010",9808 => "11011010",9809 => "11100111",9810 => "01011111",9811 => "00111011",9812 => "11010101",9813 => "01010011",9814 => "00000101",9815 => "01001001",9816 => "10011010",9817 => "01110110",9818 => "10100110",9819 => "11011010",9820 => "11011011",9821 => "10000011",9822 => "00111001",9823 => "01100011",9824 => "11101101",9825 => "11001000",9826 => "11111100",9827 => "00100101",9828 => "01110000",9829 => "00100101",9830 => "00111000",9831 => "01100110",9832 => "10100000",9833 => "01101111",9834 => "10111100",9835 => "10001000",9836 => "10111111",9837 => "00111011",9838 => "10100011",9839 => "01100100",9840 => "00000110",9841 => "10110010",9842 => "01000010",9843 => "10000100",9844 => "01100100",9845 => "00100000",9846 => "11000000",9847 => "10101010",9848 => "11010001",9849 => "01100001",9850 => "01000111",9851 => "01010010",9852 => "10011000",9853 => "00100001",9854 => "00000011",9855 => "00000011",9856 => "01100000",9857 => "01110100",9858 => "10100101",9859 => "00110000",9860 => "01011000",9861 => "00010111",9862 => "01111010",9863 => "01011001",9864 => "00010010",9865 => "00101011",9866 => "01000110",9867 => "01111000",9868 => "11000111",9869 => "11101111",9870 => "01011001",9871 => "10001001",9872 => "10111011",9873 => "11100010",9874 => "11011100",9875 => "11110010",9876 => "11110010",9877 => "00001100",9878 => "01001110",9879 => "01000100",9880 => "00100001",9881 => "11101111",9882 => "11000101",9883 => "01100111",9884 => "00001100",9885 => "10000111",9886 => "01011001",9887 => "11001101",9888 => "01110110",9889 => "01011111",9890 => "00100000",9891 => "01100110",9892 => "11001111",9893 => "01001011",9894 => "10000010",9895 => "10110011",9896 => "11110100",9897 => "11001111",9898 => "11010010",9899 => "10111001",9900 => "11010110",9901 => "00000100",9902 => "11011010",9903 => "00001000",9904 => "01010000",9905 => "10101100",9906 => "11110001",9907 => "10001001",9908 => "00110010",9909 => "01100011",9910 => "10101111",9911 => "10001000",9912 => "00000010",9913 => "10111110",9914 => "10111101",9915 => "10011100",9916 => "11011111",9917 => "00101011",9918 => "11001101",9919 => "01101001",9920 => "01010000",9921 => "01000100",9922 => "10000100",9923 => "10100010",9924 => "00100100",9925 => "00111101",9926 => "00011011",9927 => "11111001",9928 => "00010111",9929 => "11000111",9930 => "00110110",9931 => "11101110",9932 => "11110001",9933 => "11111100",9934 => "11001100",9935 => "10000110",9936 => "11000100",9937 => "00011100",9938 => "00100111",9939 => "01101001",9940 => "00100100",9941 => "11111100",9942 => "01110011",9943 => "11010100",9944 => "10111100",9945 => "10111100",9946 => "10110000",9947 => "10000001",9948 => "10111101",9949 => "01010111",9950 => "11111111",9951 => "01100000",9952 => "00011111",9953 => "01111010",9954 => "00011111",9955 => "01001001",9956 => "10011011",9957 => "11100000",9958 => "11111011",9959 => "00011001",9960 => "11101111",9961 => "01101101",9962 => "10101011",9963 => "11101011",9964 => "10000011",9965 => "01110111",9966 => "00101100",9967 => "11000101",9968 => "11000011",9969 => "11000110",9970 => "10000000",9971 => "11110110",9972 => "01010111",9973 => "10100011",9974 => "00100011",9975 => "10010000",9976 => "00000011",9977 => "10011000",9978 => "11000001",9979 => "10001100",9980 => "11000100",9981 => "01100101",9982 => "10100111",9983 => "01010101",9984 => "01111010",9985 => "00011111",9986 => "01111101",9987 => "01010101",9988 => "00011000",9989 => "00000110",9990 => "00010100",9991 => "10010000",9992 => "10101000",9993 => "01001110",9994 => "11001001",9995 => "01010011",9996 => "01010110",9997 => "10110100",9998 => "11111110",9999 => "10111100",10000 => "00100101",10001 => "10111100",10002 => "00011001",10003 => "01100011",10004 => "10000101",10005 => "00101001",10006 => "00010100",10007 => "00110001",10008 => "01000101",10009 => "10110000",10010 => "01011100",10011 => "01011010",10012 => "01010010",10013 => "11110111",10014 => "10110110",10015 => "11111001",10016 => "10000110",10017 => "11101111",10018 => "11011001",10019 => "01011101",10020 => "10101110",10021 => "01011100",10022 => "10010010",10023 => "00011111",10024 => "01101000",10025 => "11101001",10026 => "00110011",10027 => "00001001",10028 => "00101100",10029 => "00010100",10030 => "00111110",10031 => "11010101",10032 => "11000111",10033 => "10011111",10034 => "11011101",10035 => "01111010",10036 => "00001000",10037 => "01101110",10038 => "01110100",10039 => "11010110",10040 => "11010100",10041 => "01101001",10042 => "01101001",10043 => "00011101",10044 => "01101000",10045 => "01000000",10046 => "11110101",10047 => "11100100",10048 => "01000110",10049 => "10111001",10050 => "11011010",10051 => "11011011",10052 => "10111101",10053 => "01011000",10054 => "10011011",10055 => "00001010",10056 => "01101100",10057 => "01000110",10058 => "00100011",10059 => "10100110",10060 => "11000100",10061 => "11101100",10062 => "00111110",10063 => "01001010",10064 => "01100111",10065 => "11100101",10066 => "00100101",10067 => "01101011",10068 => "11001000",10069 => "01011111",10070 => "10011110",10071 => "10001000",10072 => "01101000",10073 => "10000011",10074 => "00101001",10075 => "10110111",10076 => "10011101",10077 => "01100110",10078 => "00110001",10079 => "11111011",10080 => "01110110",10081 => "01000111",10082 => "01100101",10083 => "00010011",10084 => "01000110",10085 => "01011001",10086 => "01000001",10087 => "01110100",10088 => "00100101",10089 => "10000010",10090 => "11110110",10091 => "01010111",10092 => "01100001",10093 => "00000101",10094 => "01011100",10095 => "11101011",10096 => "10100010",10097 => "11101101",10098 => "11101010",10099 => "01111000",10100 => "00101110",10101 => "00000110",10102 => "11010101",10103 => "11110110",10104 => "10001001",10105 => "11100100",10106 => "11111111",10107 => "11110000",10108 => "10100101",10109 => "10100101",10110 => "00111101",10111 => "11001000",10112 => "01001101",10113 => "00001110",10114 => "01011110",10115 => "01001001",10116 => "00100100",10117 => "10100001",10118 => "11010011",10119 => "01111101",10120 => "00001000",10121 => "00010110",10122 => "11001110",10123 => "11010100",10124 => "00110101",10125 => "00010010",10126 => "11110111",10127 => "00100010",10128 => "00101110",10129 => "00101011",10130 => "11110111",10131 => "00011111",10132 => "00011101",10133 => "00010001",10134 => "10100000",10135 => "10101101",10136 => "11100100",10137 => "00110010",10138 => "10100001",10139 => "11011011",10140 => "01100110",10141 => "11001001",10142 => "01000110",10143 => "11111100",10144 => "10010101",10145 => "11100111",10146 => "00100000",10147 => "00110000",10148 => "00001011",10149 => "01011000",10150 => "01110000",10151 => "11010100",10152 => "00101000",10153 => "10000000",10154 => "10010101",10155 => "01111101",10156 => "01100011",10157 => "01111011",10158 => "11100010",10159 => "01100011",10160 => "11001000",10161 => "00100000",10162 => "01010100",10163 => "00000000",10164 => "11000110",10165 => "11110100",10166 => "10000000",10167 => "00101010",10168 => "10000000",10169 => "10100001",10170 => "01001111",10171 => "10111011",10172 => "01001000",10173 => "00010001",10174 => "00000110",10175 => "10111001",10176 => "11000011",10177 => "01101101",10178 => "00110110",10179 => "11111100",10180 => "11100100",10181 => "01110000",10182 => "10101100",10183 => "00111100",10184 => "00111101",10185 => "10111000",10186 => "00100001",10187 => "11010111",10188 => "10110010",10189 => "11100101",10190 => "11100001",10191 => "10110110",10192 => "00001110",10193 => "11011001",10194 => "11000110",10195 => "00110101",10196 => "01001100",10197 => "01110100",10198 => "00001101",10199 => "01000010",10200 => "11111000",10201 => "11110001",10202 => "10001100",10203 => "10111101",10204 => "01101100",10205 => "00111100",10206 => "11110110",10207 => "10001111",10208 => "01011110",10209 => "10000111",10210 => "00100000",10211 => "10110011",10212 => "10110000",10213 => "10001111",10214 => "00000000",10215 => "01000101",10216 => "11100111",10217 => "10101001",10218 => "10001000",10219 => "11001001",10220 => "01001100",10221 => "11101110",10222 => "01110110",10223 => "10001111",10224 => "00000001",10225 => "10111001",10226 => "11000101",10227 => "01101110",10228 => "01010110",10229 => "11111110",10230 => "11000100",10231 => "00110101",10232 => "01010000",10233 => "00000001",10234 => "00111101",10235 => "11000001",10236 => "10100011",10237 => "01010101",10238 => "00101111",10239 => "10110000",10240 => "10001111",10241 => "01000101",10242 => "11011010",10243 => "11011111",10244 => "10111010",10245 => "11111110",10246 => "01000000",10247 => "01100010",10248 => "10111011",10249 => "11011101",10250 => "00011110",10251 => "11101110",10252 => "10111010",10253 => "00110110",10254 => "01100001",10255 => "00101111",10256 => "11111101",10257 => "10110111",10258 => "00000000",10259 => "10110010",10260 => "11110010",10261 => "00010100",10262 => "01011010",10263 => "11110010",10264 => "10001001",10265 => "00010111",10266 => "00010101",10267 => "00011101",10268 => "01100001",10269 => "10011010",10270 => "11010111",10271 => "10001100",10272 => "11111011",10273 => "00101001",10274 => "10010000",10275 => "10110101",10276 => "01010111",10277 => "10101010",10278 => "01111111",10279 => "00101100",10280 => "10101011",10281 => "01110110",10282 => "01100000",10283 => "11011010",10284 => "10101000",10285 => "11100011",10286 => "00001101",10287 => "11100000",10288 => "11100100",10289 => "11000000",10290 => "00110001",10291 => "11000100",10292 => "00011000",10293 => "10001011",10294 => "10010110",10295 => "10100000",10296 => "00110110",10297 => "01111011",10298 => "11110011",10299 => "00100100",10300 => "00101111",10301 => "11101000",10302 => "11010010",10303 => "10001101",10304 => "00001010",10305 => "10000010",10306 => "01101111",10307 => "01001111",10308 => "11111101",10309 => "01000010",10310 => "01010101",10311 => "00010000",10312 => "01001001",10313 => "11101101",10314 => "10001111",10315 => "01010100",10316 => "01001110",10317 => "11001000",10318 => "11100001",10319 => "00100101",10320 => "11011100",10321 => "10110010",10322 => "11100011",10323 => "00000010",10324 => "10001100",10325 => "00101110",10326 => "01001001",10327 => "00110011",10328 => "11001101",10329 => "00111000",10330 => "01110010",10331 => "11000000",10332 => "00100111",10333 => "01011110",10334 => "10100111",10335 => "01110000",10336 => "10000101",10337 => "01010010",10338 => "01111010",10339 => "01101111",10340 => "11110111",10341 => "11001000",10342 => "11010110",10343 => "10010110",10344 => "10110111",10345 => "01100111",10346 => "01110000",10347 => "10000001",10348 => "00001000",10349 => "01001111",10350 => "10011011",10351 => "00010001",10352 => "11000111",10353 => "01110011",10354 => "01001000",10355 => "10011000",10356 => "11111101",10357 => "10100100",10358 => "00101001",10359 => "10010111",10360 => "00101000",10361 => "00101110",10362 => "10010001",10363 => "11011101",10364 => "10000101",10365 => "00010010",10366 => "01010111",10367 => "00100011",10368 => "00101001",10369 => "01000101",10370 => "01100000",10371 => "11111010",10372 => "01001011",10373 => "01001100",10374 => "01001110",10375 => "00011111",10376 => "11100010",10377 => "00101000",10378 => "11010110",10379 => "11101010",10380 => "10100111",10381 => "00101001",10382 => "00001001",10383 => "10000111",10384 => "11001000",10385 => "11000000",10386 => "11110010",10387 => "11111001",10388 => "11110101",10389 => "00000111",10390 => "01100111",10391 => "10000110",10392 => "10100100",10393 => "00001111",10394 => "00100111",10395 => "11101010",10396 => "10110110",10397 => "10010010",10398 => "11010100",10399 => "01100111",10400 => "01000011",10401 => "01111100",10402 => "00011100",10403 => "01011101",10404 => "00011101",10405 => "00011011",10406 => "01100100",10407 => "11101101",10408 => "01100010",10409 => "01011101",10410 => "01110110",10411 => "10011101",10412 => "11101110",10413 => "11111100",10414 => "00011010",10415 => "10100010",10416 => "01110101",10417 => "10100011",10418 => "01010110",10419 => "01000100",10420 => "00011001",10421 => "01010111",10422 => "10001010",10423 => "10011101",10424 => "11111101",10425 => "01001100",10426 => "10000110",10427 => "00000001",10428 => "01100110",10429 => "11111110",10430 => "10111010",10431 => "01011111",10432 => "11111110",10433 => "10101000",10434 => "01111011",10435 => "11110100",10436 => "11011001",10437 => "01110001",10438 => "10111100",10439 => "01110011",10440 => "10110101",10441 => "01101100",10442 => "00111111",10443 => "11000110",10444 => "01001110",10445 => "11111100",10446 => "10011011",10447 => "10100000",10448 => "00010000",10449 => "10000000",10450 => "00010100",10451 => "00011011",10452 => "00100100",10453 => "00111100",10454 => "00100011",10455 => "00110000",10456 => "00111101",10457 => "01000001",10458 => "00110100",10459 => "11111101",10460 => "11111000",10461 => "10001111",10462 => "10010110",10463 => "00110111",10464 => "10011110",10465 => "10001001",10466 => "00101001",10467 => "00010001",10468 => "10111100",10469 => "10010110",10470 => "10100110",10471 => "10000010",10472 => "10111001",10473 => "11110001",10474 => "01101101",10475 => "00010011",10476 => "01110111",10477 => "00100101",10478 => "11010111",10479 => "10111010",10480 => "00111011",10481 => "00000100",10482 => "11001101",10483 => "11001010",10484 => "10010010",10485 => "10100011",10486 => "11011110",10487 => "01110110",10488 => "00100101",10489 => "10011110",10490 => "10101100",10491 => "11111100",10492 => "01110101",10493 => "10000011",10494 => "11101000",10495 => "11011011",10496 => "00000110",10497 => "10101010",10498 => "10100010",10499 => "01001100",10500 => "10001110",10501 => "10000000",10502 => "00001101",10503 => "01101100",10504 => "01101111",10505 => "01011001",10506 => "10000100",10507 => "00101011",10508 => "10110101",10509 => "01101001",10510 => "11100011",10511 => "01111100",10512 => "10001000",10513 => "11111100",10514 => "11000001",10515 => "01011011",10516 => "10010100",10517 => "10100100",10518 => "10011000",10519 => "11100100",10520 => "11101101",10521 => "00100010",10522 => "00001011",10523 => "10100010",10524 => "11111111",10525 => "00010111",10526 => "00010010",10527 => "11001001",10528 => "10011001",10529 => "10101111",10530 => "01100100",10531 => "11100001",10532 => "00010000",10533 => "11110101",10534 => "00101111",10535 => "00011011",10536 => "00011111",10537 => "01010011",10538 => "10101010",10539 => "01011111",10540 => "11011001",10541 => "01101010",10542 => "00000101",10543 => "01101011",10544 => "00110100",10545 => "11110010",10546 => "00011101",10547 => "01011010",10548 => "11110010",10549 => "11111001",10550 => "01000001",10551 => "01101110",10552 => "11001110",10553 => "11101110",10554 => "00110011",10555 => "11100111",10556 => "01001011",10557 => "11111100",10558 => "11101010",10559 => "01011101",10560 => "00111000",10561 => "01011011",10562 => "01100011",10563 => "01011001",10564 => "10000111",10565 => "00111000",10566 => "00011001",10567 => "10011001",10568 => "00111110",10569 => "10110100",10570 => "00101111",10571 => "10001010",10572 => "10101100",10573 => "11101100",10574 => "01100111",10575 => "10110110",10576 => "10111100",10577 => "01011101",10578 => "10100111",10579 => "00111110",10580 => "01010001",10581 => "11111011",10582 => "00111001",10583 => "01100010",10584 => "01110011",10585 => "10011101",10586 => "00011111",10587 => "11111010",10588 => "01011100",10589 => "00111000",10590 => "10110001",10591 => "11001100",10592 => "01000100",10593 => "00100001",10594 => "10101111",10595 => "01110000",10596 => "11011100",10597 => "10010011",10598 => "00101000",10599 => "11011011",10600 => "11110110",10601 => "01000101",10602 => "01011101",10603 => "10011101",10604 => "11110110",10605 => "10111000",10606 => "11001001",10607 => "00111110",10608 => "00000011",10609 => "00110011",10610 => "01000110",10611 => "11100011",10612 => "00110000",10613 => "10110001",10614 => "11110011",10615 => "00011010",10616 => "01010100",10617 => "01110110",10618 => "01111101",10619 => "01001011",10620 => "00010110",10621 => "11111110",10622 => "00001011",10623 => "00101001",10624 => "01011101",10625 => "11100011",10626 => "00011101",10627 => "01000001",10628 => "01100111",10629 => "01110101",10630 => "11110111",10631 => "00011001",10632 => "00111100",10633 => "00110100",10634 => "01000011",10635 => "01110001",10636 => "11010101",10637 => "11010110",10638 => "01010000",10639 => "11110111",10640 => "10100111",10641 => "10100100",10642 => "00000101",10643 => "01110011",10644 => "11010011",10645 => "11111011",10646 => "01011110",10647 => "01000110",10648 => "01001000",10649 => "01100100",10650 => "11000111",10651 => "10001110",10652 => "11010010",10653 => "00111011",10654 => "10000110",10655 => "11011000",10656 => "00110011",10657 => "11011010",10658 => "01011011",10659 => "00101010",10660 => "00111000",10661 => "01001111",10662 => "00111011",10663 => "11111111",10664 => "00111101",10665 => "01101100",10666 => "01011111",10667 => "11101010",10668 => "11101010",10669 => "10000011",10670 => "00010110",10671 => "00100001",10672 => "11001000",10673 => "00100100",10674 => "11111101",10675 => "01011011",10676 => "01100010",10677 => "01101011",10678 => "10110111",10679 => "01001111",10680 => "00111111",10681 => "00110100",10682 => "01101000",10683 => "11101001",10684 => "10000101",10685 => "01100001",10686 => "00100100",10687 => "11100101",10688 => "01110001",10689 => "00000110",10690 => "01110000",10691 => "11001000",10692 => "01100000",10693 => "01101100",10694 => "01011101",10695 => "10100001",10696 => "00010110",10697 => "00011111",10698 => "01110000",10699 => "11101001",10700 => "10111000",10701 => "00000100",10702 => "11101111",10703 => "11000101",10704 => "10111111",10705 => "10001011",10706 => "00010011",10707 => "00001100",10708 => "01100111",10709 => "00101000",10710 => "00010100",10711 => "11101101",10712 => "10000110",10713 => "00101100",10714 => "11100001",10715 => "00010010",10716 => "11101110",10717 => "01001100",10718 => "11110111",10719 => "10101001",10720 => "11000011",10721 => "11000111",10722 => "11101111",10723 => "01001011",10724 => "11110010",10725 => "10100111",10726 => "00100011",10727 => "01001011",10728 => "10011001",10729 => "11100110",10730 => "11111111",10731 => "10001101",10732 => "10100010",10733 => "00010101",10734 => "00000011",10735 => "00000001",10736 => "10101010",10737 => "10001010",10738 => "11111101",10739 => "10101000",10740 => "00111110",10741 => "10101010",10742 => "10110000",10743 => "11101100",10744 => "01100110",10745 => "00010011",10746 => "11000011",10747 => "01111111",10748 => "01001001",10749 => "11010011",10750 => "01101011",10751 => "10111110",10752 => "11000100",10753 => "10011110",10754 => "10111111",10755 => "10100011",10756 => "11010111",10757 => "11010010",10758 => "01100111",10759 => "11001100",10760 => "01000101",10761 => "10001011",10762 => "10100010",10763 => "10100001",10764 => "11001010",10765 => "11111010",10766 => "01111100",10767 => "10001000",10768 => "01110010",10769 => "01111001",10770 => "00000101",10771 => "00010110",10772 => "10101010",10773 => "01000010",10774 => "01101000",10775 => "01101010",10776 => "10100001",10777 => "00000101",10778 => "11000100",10779 => "01000000",10780 => "00001101",10781 => "10111100",10782 => "10110110",10783 => "11111111",10784 => "11100010",10785 => "11001010",10786 => "01111011",10787 => "01100100",10788 => "10100011",10789 => "10011001",10790 => "11010000",10791 => "10111110",10792 => "10110101",10793 => "01010010",10794 => "01010000",10795 => "00001101",10796 => "10011110",10797 => "00011011",10798 => "10101000",10799 => "11000001",10800 => "00010111",10801 => "10101100",10802 => "10110010",10803 => "11000010",10804 => "00000001",10805 => "11011011",10806 => "10101100",10807 => "00111011",10808 => "00101111",10809 => "10000110",10810 => "01110100",10811 => "10011110",10812 => "11010010",10813 => "00011101",10814 => "11100000",10815 => "01011001",10816 => "00100011",10817 => "00000111",10818 => "00100010",10819 => "01110101",10820 => "10111011",10821 => "01010000",10822 => "01000111",10823 => "00100001",10824 => "00110111",10825 => "00100000",10826 => "01110001",10827 => "10010000",10828 => "11100111",10829 => "00011100",10830 => "01111110",10831 => "10010100",10832 => "01001011",10833 => "01001011",10834 => "11011110",10835 => "01001101",10836 => "11110000",10837 => "00010101",10838 => "10000011",10839 => "01101000",10840 => "01111111",10841 => "10100101",10842 => "01111101",10843 => "00011001",10844 => "01011111",10845 => "11110011",10846 => "00011010",10847 => "00111100",10848 => "10111110",10849 => "10010001",10850 => "00100101",10851 => "10000110",10852 => "00101110",10853 => "10001101",10854 => "01000011",10855 => "11010011",10856 => "00110011",10857 => "11110011",10858 => "00001011",10859 => "10010101",10860 => "11111010",10861 => "10011010",10862 => "11101001",10863 => "00000010",10864 => "01111110",10865 => "00111010",10866 => "00101111",10867 => "01001010",10868 => "11110100",10869 => "11000010",10870 => "11110001",10871 => "11010000",10872 => "01001010",10873 => "01101010",10874 => "11010011",10875 => "10010110",10876 => "01011000",10877 => "01001100",10878 => "11000110",10879 => "11111011",10880 => "00011011",10881 => "00000010",10882 => "10010110",10883 => "01111010",10884 => "00101000",10885 => "01001110",10886 => "10101101",10887 => "11111000",10888 => "01001100",10889 => "01000101",10890 => "00101010",10891 => "11111001",10892 => "11100000",10893 => "01011100",10894 => "01010011",10895 => "00111110",10896 => "00001010",10897 => "11110110",10898 => "01100001",10899 => "00001110",10900 => "01000100",10901 => "10100101",10902 => "00001010",10903 => "01001011",10904 => "00001100",10905 => "00110110",10906 => "10101010",10907 => "00010100",10908 => "11010101",10909 => "10011101",10910 => "00000100",10911 => "01111111",10912 => "11110101",10913 => "01111000",10914 => "01000101",10915 => "11101000",10916 => "00000100",10917 => "01100000",10918 => "00100111",10919 => "11100010",10920 => "01111111",10921 => "11001111",10922 => "01001111",10923 => "00101111",10924 => "11011001",10925 => "10111010",10926 => "01010110",10927 => "10110100",10928 => "10010111",10929 => "00101111",10930 => "10010011",10931 => "10111110",10932 => "01101000",10933 => "00101111",10934 => "11110100",10935 => "01111001",10936 => "00101100",10937 => "01001110",10938 => "01101101",10939 => "10001011",10940 => "11101000",10941 => "01111101",10942 => "00001110",10943 => "00000101",10944 => "00100010",10945 => "10010110",10946 => "00000110",10947 => "10000011",10948 => "10000001",10949 => "00110001",10950 => "11111010",10951 => "11101001",10952 => "01010010",10953 => "01110101",10954 => "00101010",10955 => "00101000",10956 => "00111110",10957 => "11011100",10958 => "00100101",10959 => "00101000",10960 => "00011000",10961 => "00111010",10962 => "01001001",10963 => "00100010",10964 => "01010111",10965 => "11010101",10966 => "00100001",10967 => "10010110",10968 => "00111010",10969 => "00001010",10970 => "01001101",10971 => "11011010",10972 => "00101011",10973 => "11110101",10974 => "11110100",10975 => "11010110",10976 => "01011000",10977 => "11001010",10978 => "10100010",10979 => "01111101",10980 => "10000110",10981 => "11100101",10982 => "10110100",10983 => "01100001",10984 => "11011100",10985 => "11111000",10986 => "10001110",10987 => "10111001",10988 => "00011110",10989 => "11100001",10990 => "00101001",10991 => "11111000",10992 => "11000111",10993 => "11010100",10994 => "11111111",10995 => "10001111",10996 => "10001010",10997 => "01001110",10998 => "11101010",10999 => "10110001",11000 => "00011101",11001 => "01100011",11002 => "01110111",11003 => "10001010",11004 => "01101101",11005 => "00010000",11006 => "01111110",11007 => "11101001",11008 => "01100010",11009 => "10110101",11010 => "01000110",11011 => "00001110",11012 => "10011110",11013 => "01101110",11014 => "00101100",11015 => "01000100",11016 => "00111000",11017 => "11110101",11018 => "10001110",11019 => "00001000",11020 => "11000111",11021 => "00000011",11022 => "01110000",11023 => "01111100",11024 => "01111101",11025 => "11000010",11026 => "00011101",11027 => "10111011",11028 => "00000001",11029 => "11101100",11030 => "00000001",11031 => "10110000",11032 => "10101110",11033 => "00011100",11034 => "11000010",11035 => "10101110",11036 => "10001000",11037 => "10010000",11038 => "11100001",11039 => "01110101",11040 => "01000010",11041 => "01110000",11042 => "11001010",11043 => "11100111",11044 => "01000110",11045 => "11111110",11046 => "01100110",11047 => "01111001",11048 => "00011011",11049 => "00111110",11050 => "01000101",11051 => "11000000",11052 => "00100010",11053 => "11001100",11054 => "00111100",11055 => "11100110",11056 => "01011001",11057 => "00100111",11058 => "00000100",11059 => "11100001",11060 => "00101100",11061 => "10111010",11062 => "00001101",11063 => "00011001",11064 => "01110000",11065 => "11001101",11066 => "00110100",11067 => "01010100",11068 => "01110101",11069 => "11011111",11070 => "10010010",11071 => "00100100",11072 => "10111110",11073 => "01001010",11074 => "00100100",11075 => "00011010",11076 => "00011011",11077 => "11101110",11078 => "01100101",11079 => "01011001",11080 => "01110100",11081 => "11101000",11082 => "10011000",11083 => "11011111",11084 => "11110011",11085 => "00001110",11086 => "01000101",11087 => "11101111",11088 => "01010010",11089 => "11111110",11090 => "01100100",11091 => "00101110",11092 => "11001000",11093 => "11101011",11094 => "00110100",11095 => "01010001",11096 => "01010010",11097 => "00010001",11098 => "10101111",11099 => "00110010",11100 => "01000111",11101 => "00001101",11102 => "10010111",11103 => "00011001",11104 => "01011101",11105 => "11001111",11106 => "11000011",11107 => "10010100",11108 => "10001011",11109 => "00001101",11110 => "11010010",11111 => "00001000",11112 => "10001011",11113 => "10011101",11114 => "00000110",11115 => "10100000",11116 => "00101101",11117 => "11111100",11118 => "10100010",11119 => "01001011",11120 => "00100111",11121 => "10111000",11122 => "01100010",11123 => "00001001",11124 => "10010100",11125 => "00000101",11126 => "00000110",11127 => "01101101",11128 => "00010001",11129 => "11001000",11130 => "10100011",11131 => "00011100",11132 => "01100011",11133 => "00000110",11134 => "11000100",11135 => "10000001",11136 => "01111111",11137 => "11111100",11138 => "11100011",11139 => "10011100",11140 => "00010001",11141 => "10110110",11142 => "01010100",11143 => "00111001",11144 => "10100011",11145 => "00011110",11146 => "00101000",11147 => "00010100",11148 => "01101011",11149 => "00010011",11150 => "10000111",11151 => "11000011",11152 => "11010010",11153 => "01111101",11154 => "00001001",11155 => "00100100",11156 => "10111010",11157 => "01111100",11158 => "11101101",11159 => "00010011",11160 => "01100100",11161 => "11000000",11162 => "00000111",11163 => "11101000",11164 => "00010000",11165 => "10111110",11166 => "01001000",11167 => "11110110",11168 => "01100011",11169 => "00100010",11170 => "01010101",11171 => "00110111",11172 => "11110011",11173 => "10110101",11174 => "01111001",11175 => "11000001",11176 => "00010010",11177 => "11000100",11178 => "10111111",11179 => "11101111",11180 => "10000011",11181 => "11011110",11182 => "01001011",11183 => "11001101",11184 => "00000101",11185 => "10000001",11186 => "01100101",11187 => "10111011",11188 => "00010110",11189 => "00110101",11190 => "00101000",11191 => "00110000",11192 => "10110111",11193 => "11100100",11194 => "11011000",11195 => "01001101",11196 => "11001001",11197 => "11001100",11198 => "00000001",11199 => "11011001",11200 => "11101011",11201 => "01011111",11202 => "00100011",11203 => "00000000",11204 => "01011011",11205 => "10011010",11206 => "00010101",11207 => "11011101",11208 => "11011100",11209 => "10011001",11210 => "10110100",11211 => "01100000",11212 => "10110000",11213 => "00100100",11214 => "01100010",11215 => "00011000",11216 => "11100001",11217 => "11001011",11218 => "00101111",11219 => "10101001",11220 => "00100001",11221 => "01101000",11222 => "00101101",11223 => "11010110",11224 => "10000101",11225 => "10011010",11226 => "10001011",11227 => "00111011",11228 => "11111100",11229 => "11001111",11230 => "11110011",11231 => "01100000",11232 => "01101001",11233 => "10101001",11234 => "11101101",11235 => "11001001",11236 => "00111110",11237 => "01011110",11238 => "11010101",11239 => "01001010",11240 => "10010010",11241 => "11011010",11242 => "11010001",11243 => "00010010",11244 => "11011001",11245 => "11011100",11246 => "00110110",11247 => "01000011",11248 => "10110011",11249 => "10010010",11250 => "01011011",11251 => "00111101",11252 => "01010110",11253 => "10101010",11254 => "11101001",11255 => "10111101",11256 => "10000011",11257 => "00010011",11258 => "00000111",11259 => "01010001",11260 => "10111001",11261 => "01011110",11262 => "01110111",11263 => "00011001",11264 => "11110000",11265 => "00110101",11266 => "11110011",11267 => "00100010",11268 => "01000000",11269 => "10101000",11270 => "01110110",11271 => "01100010",11272 => "01010010",11273 => "01011011",11274 => "00010111",11275 => "01100011",11276 => "01001001",11277 => "00000110",11278 => "01010000",11279 => "00001110",11280 => "00101100",11281 => "00110101",11282 => "11001001",11283 => "01100100",11284 => "00101100",11285 => "10011010",11286 => "01010111",11287 => "00100010",11288 => "00110101",11289 => "11110101",11290 => "10111001",11291 => "01101011",11292 => "01110010",11293 => "00000000",11294 => "10111101",11295 => "11101100",11296 => "00111011",11297 => "00100110",11298 => "01100010",11299 => "11110010",11300 => "01001001",11301 => "11011111",11302 => "11000111",11303 => "11100001",11304 => "11001110",11305 => "11001111",11306 => "00111101",11307 => "11110001",11308 => "00101110",11309 => "01101000",11310 => "01001000",11311 => "01101011",11312 => "01011010",11313 => "00101010",11314 => "01011001",11315 => "01101100",11316 => "00011001",11317 => "01000101",11318 => "01101101",11319 => "01111000",11320 => "01110010",11321 => "10000101",11322 => "10000100",11323 => "01110101",11324 => "01001001",11325 => "00100110",11326 => "11101110",11327 => "00001010",11328 => "01111110",11329 => "00001010",11330 => "01000111",11331 => "11010111",11332 => "00010111",11333 => "00100101",11334 => "10101110",11335 => "11110001",11336 => "11011101",11337 => "01101000",11338 => "11101110",11339 => "00010010",11340 => "10100111",11341 => "10001010",11342 => "10010001",11343 => "00010001",11344 => "11110000",11345 => "11110110",11346 => "11101010",11347 => "10001011",11348 => "00111011",11349 => "00101101",11350 => "10111101",11351 => "11110100",11352 => "00110001",11353 => "11010101",11354 => "01110000",11355 => "11100000",11356 => "11110111",11357 => "01011111",11358 => "10100010",11359 => "11000011",11360 => "00011000",11361 => "01111110",11362 => "11010010",11363 => "11101001",11364 => "01000100",11365 => "01101010",11366 => "01110110",11367 => "10000110",11368 => "00000111",11369 => "10100001",11370 => "01011101",11371 => "10111100",11372 => "11100110",11373 => "11000110",11374 => "10101100",11375 => "01010100",11376 => "01110011",11377 => "00001100",11378 => "11010001",11379 => "00010000",11380 => "01000111",11381 => "10111001",11382 => "01101010",11383 => "10110001",11384 => "01100010",11385 => "10001011",11386 => "00110100",11387 => "01001000",11388 => "01111010",11389 => "00010111",11390 => "10001001",11391 => "11000101",11392 => "11110101",11393 => "11100110",11394 => "01010001",11395 => "10000111",11396 => "00001110",11397 => "00111111",11398 => "10000011",11399 => "01011111",11400 => "01110101",11401 => "11110110",11402 => "00000001",11403 => "01100110",11404 => "01100101",11405 => "00101110",11406 => "10000111",11407 => "11001011",11408 => "10001110",11409 => "01001001",11410 => "01010101",11411 => "00101101",11412 => "10001110",11413 => "01101000",11414 => "10100000",11415 => "10001001",11416 => "11100011",11417 => "10100010",11418 => "11010011",11419 => "01011110",11420 => "11101011",11421 => "10000110",11422 => "10111101",11423 => "00011111",11424 => "00010011",11425 => "11110011",11426 => "01111101",11427 => "01000011",11428 => "10001101",11429 => "11111000",11430 => "11010101",11431 => "10111010",11432 => "01010000",11433 => "01011111",11434 => "01110010",11435 => "11111001",11436 => "10011001",11437 => "00000111",11438 => "10011011",11439 => "11100000",11440 => "00111100",11441 => "01111000",11442 => "11100110",11443 => "01110100",11444 => "00001000",11445 => "00001110",11446 => "00001001",11447 => "11101001",11448 => "01100110",11449 => "00001010",11450 => "10100100",11451 => "11101111",11452 => "00000100",11453 => "10010111",11454 => "11011001",11455 => "10000001",11456 => "11001011",11457 => "00001010",11458 => "00011010",11459 => "01111100",11460 => "00010101",11461 => "11111111",11462 => "11111111",11463 => "10100111",11464 => "10100000",11465 => "11111100",11466 => "10011111",11467 => "11010010",11468 => "00001100",11469 => "00010001",11470 => "00101110",11471 => "00111000",11472 => "11101011",11473 => "11101101",11474 => "11110011",11475 => "01100101",11476 => "00001011",11477 => "01000010",11478 => "11010110",11479 => "01011101",11480 => "00100110",11481 => "10100010",11482 => "00001000",11483 => "10111000",11484 => "11000101",11485 => "10010001",11486 => "00100100",11487 => "00101000",11488 => "10000010",11489 => "10100111",11490 => "11011000",11491 => "11111011",11492 => "01000011",11493 => "00010100",11494 => "00011000",11495 => "00001100",11496 => "00000110",11497 => "01100110",11498 => "00010010",11499 => "01011101",11500 => "11011111",11501 => "01110000",11502 => "01110111",11503 => "01010010",11504 => "01100100",11505 => "11100000",11506 => "00010000",11507 => "01111111",11508 => "11100000",11509 => "11101000",11510 => "10010000",11511 => "01100110",11512 => "00001101",11513 => "11010111",11514 => "01101101",11515 => "00000101",11516 => "00000100",11517 => "00001111",11518 => "11001101",11519 => "01111101",11520 => "01010011",11521 => "00011100",11522 => "00010010",11523 => "11110110",11524 => "00000010",11525 => "00000010",11526 => "10101010",11527 => "10110001",11528 => "10000000",11529 => "00011001",11530 => "01101010",11531 => "10111010",11532 => "11110011",11533 => "01110001",11534 => "10100111",11535 => "11011001",11536 => "11000001",11537 => "11011011",11538 => "11011010",11539 => "10111000",11540 => "01111110",11541 => "11011111",11542 => "00010010",11543 => "00100111",11544 => "00110000",11545 => "01001101",11546 => "11100000",11547 => "01101001",11548 => "10110110",11549 => "10111100",11550 => "11001000",11551 => "00100010",11552 => "00110101",11553 => "11100100",11554 => "10010110",11555 => "10110111",11556 => "00001110",11557 => "10100100",11558 => "00111111",11559 => "11000101",11560 => "11110000",11561 => "10011111",11562 => "00010111",11563 => "00001111",11564 => "00101000",11565 => "00110010",11566 => "00110000",11567 => "11010011",11568 => "10011110",11569 => "11001010",11570 => "11001000",11571 => "11101011",11572 => "00001001",11573 => "01011110",11574 => "11001001",11575 => "00110000",11576 => "10011001",11577 => "01100100",11578 => "11101101",11579 => "01101011",11580 => "11111001",11581 => "00010010",11582 => "00010001",11583 => "00000111",11584 => "10110011",11585 => "01101011",11586 => "00011101",11587 => "10001011",11588 => "11011011",11589 => "00010000",11590 => "01111111",11591 => "11101010",11592 => "00111011",11593 => "01010111",11594 => "10000101",11595 => "00000011",11596 => "10000010",11597 => "00010110",11598 => "11011001",11599 => "11011001",11600 => "00011111",11601 => "10000010",11602 => "10000101",11603 => "01011111",11604 => "11010100",11605 => "01110001",11606 => "00010000",11607 => "01001110",11608 => "10101100",11609 => "01010000",11610 => "10101101",11611 => "10101101",11612 => "11000110",11613 => "01111111",11614 => "01100011",11615 => "10101111",11616 => "01101000",11617 => "01101111",11618 => "10111101",11619 => "01010101",11620 => "10000100",11621 => "00101110",11622 => "00100100",11623 => "11000010",11624 => "01010011",11625 => "01011011",11626 => "00000011",11627 => "01001101",11628 => "11101000",11629 => "10111111",11630 => "10000111",11631 => "00000101",11632 => "01010011",11633 => "01101100",11634 => "11111011",11635 => "11010101",11636 => "10010111",11637 => "11010111",11638 => "11111110",11639 => "01110011",11640 => "11101110",11641 => "00110100",11642 => "10101111",11643 => "01100001",11644 => "11011100",11645 => "11010111",11646 => "01010100",11647 => "10110111",11648 => "10011011",11649 => "11101000",11650 => "10101010",11651 => "11010000",11652 => "10110110",11653 => "00010001",11654 => "11101011",11655 => "01100111",11656 => "00001111",11657 => "11111010",11658 => "00010110",11659 => "10001001",11660 => "11001101",11661 => "10001011",11662 => "01001110",11663 => "00101101",11664 => "11110011",11665 => "00010111",11666 => "10011010",11667 => "01000010",11668 => "10110101",11669 => "11001000",11670 => "11110100",11671 => "01111011",11672 => "10001010",11673 => "01001000",11674 => "00000100",11675 => "10010110",11676 => "11100100",11677 => "00010101",11678 => "11100001",11679 => "11100011",11680 => "00101000",11681 => "10100000",11682 => "10110110",11683 => "00000001",11684 => "11101101",11685 => "01011100",11686 => "10001100",11687 => "10001100",11688 => "10110110",11689 => "01011100",11690 => "10111001",11691 => "10001000",11692 => "11011111",11693 => "01011101",11694 => "00100100",11695 => "01001101",11696 => "11100000",11697 => "01000011",11698 => "11010101",11699 => "00111011",11700 => "10010001",11701 => "00010110",11702 => "01011110",11703 => "10010110",11704 => "01100100",11705 => "01000000",11706 => "11100101",11707 => "11011110",11708 => "11100000",11709 => "01100000",11710 => "01111110",11711 => "01010001",11712 => "11100001",11713 => "00111100",11714 => "00000111",11715 => "10110010",11716 => "00001011",11717 => "01010110",11718 => "10110001",11719 => "10101101",11720 => "11101000",11721 => "11011011",11722 => "10011111",11723 => "10011010",11724 => "00011110",11725 => "01110011",11726 => "11011001",11727 => "00110100",11728 => "11110000",11729 => "10101110",11730 => "01101110",11731 => "00001111",11732 => "10010011",11733 => "00010000",11734 => "10000010",11735 => "10111001",11736 => "01101000",11737 => "00110010",11738 => "00001100",11739 => "00000000",11740 => "00001110",11741 => "10101000",11742 => "00000001",11743 => "10001111",11744 => "00100110",11745 => "11110010",11746 => "11100111",11747 => "10101101",11748 => "00111010",11749 => "11110001",11750 => "10010010",11751 => "11101000",11752 => "10001001",11753 => "01000001",11754 => "11000000",11755 => "01011101",11756 => "11010101",11757 => "01101000",11758 => "01111001",11759 => "01111110",11760 => "10110000",11761 => "00101001",11762 => "11110001",11763 => "01101010",11764 => "11110111",11765 => "11100001",11766 => "10000111",11767 => "01101001",11768 => "00000000",11769 => "11010011",11770 => "10101000",11771 => "11011100",11772 => "00000100",11773 => "10100101",11774 => "00101110",11775 => "01011101",11776 => "11000101",11777 => "11000110",11778 => "11110010",11779 => "00100011",11780 => "00010100",11781 => "00010000",11782 => "00010000",11783 => "01101011",11784 => "01001000",11785 => "10011100",11786 => "10111100",11787 => "01011100",11788 => "00000101",11789 => "11000111",11790 => "11100111",11791 => "01100111",11792 => "00000101",11793 => "11101101",11794 => "00111001",11795 => "00011010",11796 => "01110110",11797 => "00100000",11798 => "00011011",11799 => "00100110",11800 => "11011101",11801 => "00110000",11802 => "00100011",11803 => "01011000",11804 => "01011101",11805 => "00110011",11806 => "10111011",11807 => "01010111",11808 => "11110011",11809 => "11100101",11810 => "11010000",11811 => "10011000",11812 => "10110011",11813 => "10001110",11814 => "10111000",11815 => "11010001",11816 => "10111011",11817 => "00111101",11818 => "01101001",11819 => "01100000",11820 => "00101110",11821 => "01110100",11822 => "11011111",11823 => "01100110",11824 => "01100011",11825 => "11000101",11826 => "11100011",11827 => "10111111",11828 => "10001110",11829 => "01110001",11830 => "11000010",11831 => "01110111",11832 => "00101010",11833 => "00011001",11834 => "11010111",11835 => "11001001",11836 => "00110000",11837 => "11011001",11838 => "00000111",11839 => "00001010",11840 => "00111001",11841 => "01100001",11842 => "00011000",11843 => "10101100",11844 => "10100000",11845 => "11000001",11846 => "11001000",11847 => "00100001",11848 => "01000000",11849 => "10011010",11850 => "00101011",11851 => "00101001",11852 => "10001101",11853 => "01010001",11854 => "10101011",11855 => "01010111",11856 => "11101101",11857 => "00001110",11858 => "11011110",11859 => "01010101",11860 => "10110101",11861 => "11000011",11862 => "10001111",11863 => "11111011",11864 => "10101101",11865 => "01110010",11866 => "11101001",11867 => "10110101",11868 => "11110100",11869 => "01100101",11870 => "01101011",11871 => "11000000",11872 => "10000010",11873 => "00000001",11874 => "01000000",11875 => "11110000",11876 => "00110101",11877 => "11100101",11878 => "11010000",11879 => "11010110",11880 => "01000001",11881 => "10100101",11882 => "10110110",11883 => "10100010",11884 => "00000010",11885 => "11011100",11886 => "11111001",11887 => "01111111",11888 => "10101011",11889 => "01101000",11890 => "11010111",11891 => "10100010",11892 => "11111010",11893 => "01001100",11894 => "00111010",11895 => "00110001",11896 => "10010011",11897 => "00000001",11898 => "11100111",11899 => "00100110",11900 => "00011000",11901 => "10101011",11902 => "01110000",11903 => "10000100",11904 => "00100100",11905 => "10011101",11906 => "11000101",11907 => "01100101",11908 => "10100101",11909 => "00001100",11910 => "00110101",11911 => "10010001",11912 => "11011110",11913 => "11010000",11914 => "01110011",11915 => "00110011",11916 => "00000011",11917 => "00110101",11918 => "10101100",11919 => "11111100",11920 => "10011011",11921 => "01110100",11922 => "11000111",11923 => "10000000",11924 => "00010110",11925 => "01100101",11926 => "10011010",11927 => "01001110",11928 => "01000011",11929 => "00011100",11930 => "11101111",11931 => "01110111",11932 => "00010011",11933 => "10010000",11934 => "00100110",11935 => "10011000",11936 => "11100110",11937 => "01011110",11938 => "11010111",11939 => "01011110",11940 => "11000101",11941 => "11100010",11942 => "11100100",11943 => "01011010",11944 => "11000111",11945 => "01000000",11946 => "00010010",11947 => "11111101",11948 => "10111011",11949 => "10000000",11950 => "10010000",11951 => "00001111",11952 => "00110011",11953 => "01111101",11954 => "00000011",11955 => "11101010",11956 => "01110101",11957 => "01011011",11958 => "00101001",11959 => "11010101",11960 => "00111000",11961 => "00001110",11962 => "01000011",11963 => "01011111",11964 => "00100001",11965 => "10001001",11966 => "00010000",11967 => "11101001",11968 => "10101011",11969 => "01110011",11970 => "11101000",11971 => "11110100",11972 => "00101101",11973 => "10110101",11974 => "10010111",11975 => "00110001",11976 => "10010100",11977 => "10111001",11978 => "11000110",11979 => "01110010",11980 => "10011111",11981 => "01001011",11982 => "00100011",11983 => "00111100",11984 => "01101100",11985 => "01101111",11986 => "11101100",11987 => "01001011",11988 => "10101110",11989 => "11001111",11990 => "01101001",11991 => "11100111",11992 => "11110111",11993 => "01011111",11994 => "00011111",11995 => "10101100",11996 => "00010101",11997 => "00111000",11998 => "00001000",11999 => "00010000",12000 => "01100000",12001 => "10000001",12002 => "00000100",12003 => "11110111",12004 => "10101111",12005 => "11100011",12006 => "01010110",12007 => "01111110",12008 => "10010110",12009 => "11001100",12010 => "00000001",12011 => "01100010",12012 => "01101000",12013 => "11001110",12014 => "10000100",12015 => "10111101",12016 => "01111100",12017 => "11000011",12018 => "01111111",12019 => "11101111",12020 => "00101100",12021 => "10000111",12022 => "00010110",12023 => "00110000",12024 => "01001101",12025 => "11110010",12026 => "10011100",12027 => "01000111",12028 => "01111001",12029 => "11000011",12030 => "01101100",12031 => "01010000",12032 => "10101000",12033 => "00100110",12034 => "00101010",12035 => "11101100",12036 => "01010001",12037 => "00010101",12038 => "11111001",12039 => "00001001",12040 => "01010010",12041 => "00010110",12042 => "00111111",12043 => "01111110",12044 => "00110110",12045 => "00010101",12046 => "10100001",12047 => "00111100",12048 => "10011001",12049 => "10011011",12050 => "10100100",12051 => "00000011",12052 => "00010001",12053 => "01101001",12054 => "01100011",12055 => "10011001",12056 => "10000100",12057 => "10001000",12058 => "11001100",12059 => "01010001",12060 => "11001011",12061 => "01010010",12062 => "11111010",12063 => "01110101",12064 => "01110101",12065 => "01111110",12066 => "01011011",12067 => "00010111",12068 => "10000100",12069 => "10110111",12070 => "01111001",12071 => "10110001",12072 => "00000100",12073 => "00010000",12074 => "01001110",12075 => "01101110",12076 => "00100100",12077 => "11100101",12078 => "10110101",12079 => "00111101",12080 => "10010111",12081 => "10001110",12082 => "11110001",12083 => "10110000",12084 => "00100100",12085 => "10101010",12086 => "00001110",12087 => "00000000",12088 => "01100011",12089 => "11011000",12090 => "01001100",12091 => "00000100",12092 => "10110000",12093 => "10001000",12094 => "11100011",12095 => "00011010",12096 => "10000101",12097 => "00100111",12098 => "11011111",12099 => "10011101",12100 => "00001010",12101 => "01111101",12102 => "10011111",12103 => "01011100",12104 => "11110011",12105 => "00101010",12106 => "01001000",12107 => "01111100",12108 => "10000100",12109 => "11100101",12110 => "10001011",12111 => "01011001",12112 => "01100101",12113 => "01011011",12114 => "01111111",12115 => "11001100",12116 => "00000001",12117 => "10011011",12118 => "11011100",12119 => "01110100",12120 => "10011010",12121 => "01000100",12122 => "00010111",12123 => "01110101",12124 => "01101011",12125 => "10000110",12126 => "01001100",12127 => "10010011",12128 => "00111110",12129 => "11100100",12130 => "01000110",12131 => "10001110",12132 => "00011011",12133 => "01010010",12134 => "01110011",12135 => "10010111",12136 => "11011000",12137 => "11111101",12138 => "00001101",12139 => "10001001",12140 => "01101010",12141 => "10111110",12142 => "10110001",12143 => "11000111",12144 => "10011001",12145 => "01100000",12146 => "01000100",12147 => "11010100",12148 => "00010010",12149 => "11001100",12150 => "10000001",12151 => "11011100",12152 => "00010100",12153 => "11100100",12154 => "01111011",12155 => "00011111",12156 => "10000000",12157 => "01111001",12158 => "10010101",12159 => "00100001",12160 => "11110000",12161 => "11101100",12162 => "00101111",12163 => "01100000",12164 => "00011011",12165 => "01000001",12166 => "01110001",12167 => "10100000",12168 => "10011110",12169 => "11001010",12170 => "11111111",12171 => "01110110",12172 => "11101101",12173 => "00100000",12174 => "11100101",12175 => "11010001",12176 => "01011101",12177 => "11101110",12178 => "00001001",12179 => "01011101",12180 => "11111110",12181 => "00011101",12182 => "01010011",12183 => "11111001",12184 => "10100101",12185 => "11011011",12186 => "11100100",12187 => "01011011",12188 => "00110100",12189 => "10100111",12190 => "10010100",12191 => "01100100",12192 => "01011111",12193 => "10111101",12194 => "10000111",12195 => "01111010",12196 => "10110000",12197 => "11110111",12198 => "00101001",12199 => "01011011",12200 => "00010100",12201 => "10010010",12202 => "01110100",12203 => "10000001",12204 => "00001011",12205 => "10000100",12206 => "10100110",12207 => "11010110",12208 => "01010110",12209 => "10001110",12210 => "10001101",12211 => "00011001",12212 => "10010101",12213 => "01001100",12214 => "11111100",12215 => "00101110",12216 => "11000000",12217 => "11111100",12218 => "10011000",12219 => "01000100",12220 => "11100101",12221 => "10100111",12222 => "11100111",12223 => "01010101",12224 => "11010011",12225 => "10010101",12226 => "11000000",12227 => "11101011",12228 => "10010101",12229 => "00011011",12230 => "00111100",12231 => "00010011",12232 => "11000000",12233 => "10001100",12234 => "11110000",12235 => "11111110",12236 => "01101010",12237 => "11110111",12238 => "00001011",12239 => "11001011",12240 => "01000011",12241 => "01110101",12242 => "11001000",12243 => "10111001",12244 => "00110111",12245 => "01011100",12246 => "11100101",12247 => "01101010",12248 => "00001110",12249 => "00011100",12250 => "10001000",12251 => "11100100",12252 => "11001101",12253 => "00100111",12254 => "10010101",12255 => "00111010",12256 => "01110011",12257 => "10001010",12258 => "01111010",12259 => "11100011",12260 => "00111011",12261 => "10111100",12262 => "01010001",12263 => "11011111",12264 => "10100101",12265 => "00001001",12266 => "11100010",12267 => "00100111",12268 => "01011100",12269 => "10010011",12270 => "00000001",12271 => "01100001",12272 => "11010100",12273 => "10011010",12274 => "00111000",12275 => "00111111",12276 => "01011100",12277 => "00110101",12278 => "01010111",12279 => "10100010",12280 => "11111001",12281 => "00000111",12282 => "11111111",12283 => "11011110",12284 => "00110000",12285 => "10100110",12286 => "11100001",12287 => "10001001",12288 => "10001011",12289 => "11011110",12290 => "10010011",12291 => "10010010",12292 => "00110000",12293 => "01100101",12294 => "10100110",12295 => "00010001",12296 => "11011000",12297 => "11111111",12298 => "00010100",12299 => "10110110",12300 => "01000001",12301 => "01101011",12302 => "10010110",12303 => "10111100",12304 => "10010100",12305 => "11011100",12306 => "01110001",12307 => "01101001",12308 => "01110000",12309 => "10010001",12310 => "01000100",12311 => "01011001",12312 => "10011111",12313 => "11101010",12314 => "01001100",12315 => "10001110",12316 => "11000011",12317 => "10101100",12318 => "11111001",12319 => "01110100",12320 => "11110110",12321 => "00111001",12322 => "10111001",12323 => "00101100",12324 => "10001110",12325 => "01010111",12326 => "01101110",12327 => "10000100",12328 => "10001101",12329 => "01000001",12330 => "11000111",12331 => "10100010",12332 => "01001110",12333 => "01100101",12334 => "11010011",12335 => "10110111",12336 => "01000000",12337 => "11111101",12338 => "00100100",12339 => "00001011",12340 => "11110111",12341 => "11001101",12342 => "00000111",12343 => "10000011",12344 => "11111001",12345 => "11101000",12346 => "10000000",12347 => "00111111",12348 => "00100101",12349 => "10111010",12350 => "00000100",12351 => "01000011",12352 => "11111000",12353 => "10001101",12354 => "10001101",12355 => "10000011",12356 => "00000011",12357 => "00111111",12358 => "11111110",12359 => "11110000",12360 => "00000111",12361 => "10111101",12362 => "01011110",12363 => "11100111",12364 => "10111011",12365 => "11011010",12366 => "00001100",12367 => "00110001",12368 => "11111100",12369 => "11111001",12370 => "00100011",12371 => "01110101",12372 => "10011100",12373 => "00111101",12374 => "00101011",12375 => "11010010",12376 => "01001010",12377 => "11001010",12378 => "10101011",12379 => "10111010",12380 => "10011010",12381 => "01110100",12382 => "00000010",12383 => "10101010",12384 => "01011000",12385 => "00000111",12386 => "01010110",12387 => "10011010",12388 => "10000100",12389 => "10010101",12390 => "00100000",12391 => "11100101",12392 => "10010101",12393 => "00011011",12394 => "11101001",12395 => "11110111",12396 => "11111111",12397 => "01110100",12398 => "01101001",12399 => "10001001",12400 => "11100001",12401 => "10100010",12402 => "10101011",12403 => "11101101",12404 => "10010111",12405 => "11110010",12406 => "00101111",12407 => "11110110",12408 => "00010110",12409 => "10001010",12410 => "00101101",12411 => "01110010",12412 => "10011100",12413 => "01100011",12414 => "10111101",12415 => "10011010",12416 => "00101100",12417 => "01010111",12418 => "11011010",12419 => "11111010",12420 => "00101011",12421 => "01011111",12422 => "01000011",12423 => "00010110",12424 => "01110110",12425 => "01110111",12426 => "01100011",12427 => "10000111",12428 => "10000011",12429 => "11001010",12430 => "01010000",12431 => "11011010",12432 => "11101101",12433 => "01010011",12434 => "10011010",12435 => "01100100",12436 => "00100011",12437 => "11011101",12438 => "01000010",12439 => "00000000",12440 => "10000101",12441 => "00110001",12442 => "01111111",12443 => "10010010",12444 => "01111100",12445 => "00101001",12446 => "01001010",12447 => "11100110",12448 => "11000101",12449 => "11110110",12450 => "10101100",12451 => "10110010",12452 => "01101100",12453 => "01110001",12454 => "01001011",12455 => "10011100",12456 => "10101001",12457 => "01000000",12458 => "10110001",12459 => "01001111",12460 => "01101110",12461 => "00101011",12462 => "10001010",12463 => "11000110",12464 => "01101011",12465 => "11101101",12466 => "01100010",12467 => "10110010",12468 => "01101000",12469 => "00010110",12470 => "11011100",12471 => "00000110",12472 => "11000011",12473 => "10000001",12474 => "11101100",12475 => "11000010",12476 => "11001110",12477 => "11001110",12478 => "01011000",12479 => "00100010",12480 => "10011001",12481 => "00100101",12482 => "01100001",12483 => "10011000",12484 => "01111101",12485 => "01000111",12486 => "00110000",12487 => "10100010",12488 => "00010011",12489 => "00010000",12490 => "00000110",12491 => "11011001",12492 => "01000101",12493 => "11100000",12494 => "00001010",12495 => "01011110",12496 => "00100010",12497 => "10011010",12498 => "00110001",12499 => "10111110",12500 => "00001000",12501 => "10000101",12502 => "10011100",12503 => "01000001",12504 => "01001000",12505 => "11001001",12506 => "11011010",12507 => "00001100",12508 => "11111111",12509 => "00100001",12510 => "11100010",12511 => "10011101",12512 => "00100111",12513 => "11110110",12514 => "10000111",12515 => "10100010",12516 => "11010100",12517 => "00000011",12518 => "01110110",12519 => "11000101",12520 => "10110000",12521 => "01111101",12522 => "01101010",12523 => "01111100",12524 => "11010010",12525 => "11010111",12526 => "11100000",12527 => "11001101",12528 => "01011011",12529 => "11111010",12530 => "11111101",12531 => "01001010",12532 => "10110100",12533 => "11010000",12534 => "10110111",12535 => "00100101",12536 => "00000001",12537 => "01100011",12538 => "11101011",12539 => "10101010",12540 => "11101011",12541 => "00001110",12542 => "10110100",12543 => "01011100",12544 => "10101001",12545 => "11110111",12546 => "11111110",12547 => "00000010",12548 => "00010000",12549 => "10010010",12550 => "01011001",12551 => "01000010",12552 => "10100000",12553 => "10111101",12554 => "00111011",12555 => "11000101",12556 => "10011111",12557 => "11000111",12558 => "11101000",12559 => "11110000",12560 => "11010111",12561 => "11010100",12562 => "11101011",12563 => "00011010",12564 => "10100110",12565 => "01101110",12566 => "00100000",12567 => "11010100",12568 => "01111101",12569 => "10011110",12570 => "01110011",12571 => "00000001",12572 => "11010100",12573 => "00010111",12574 => "01010101",12575 => "00111001",12576 => "00000001",12577 => "11000001",12578 => "01100111",12579 => "00000101",12580 => "00011110",12581 => "11011101",12582 => "10010000",12583 => "11101010",12584 => "00100010",12585 => "10110110",12586 => "10110101",12587 => "01111001",12588 => "01101011",12589 => "01001101",12590 => "01000100",12591 => "10000011",12592 => "11001111",12593 => "01111000",12594 => "01101011",12595 => "11100101",12596 => "10100111",12597 => "00011001",12598 => "00010011",12599 => "01110010",12600 => "11100110",12601 => "10010011",12602 => "10111101",12603 => "00010000",12604 => "01101010",12605 => "11110101",12606 => "10110111",12607 => "00010111",12608 => "01111000",12609 => "10011000",12610 => "11101101",12611 => "00110010",12612 => "10100011",12613 => "00010010",12614 => "00010001",12615 => "01111110",12616 => "11001001",12617 => "00110101",12618 => "00100000",12619 => "10100110",12620 => "01101000",12621 => "00010011",12622 => "10111000",12623 => "11111001",12624 => "11101010",12625 => "10111100",12626 => "00010010",12627 => "11010110",12628 => "11011001",12629 => "01010010",12630 => "00100101",12631 => "01000010",12632 => "10000100",12633 => "01101010",12634 => "00100100",12635 => "00000000",12636 => "11101011",12637 => "11001100",12638 => "00011010",12639 => "10111101",12640 => "11010101",12641 => "00110110",12642 => "11010101",12643 => "10011111",12644 => "10011010",12645 => "11110000",12646 => "00000000",12647 => "00101010",12648 => "01010110",12649 => "10110101",12650 => "10011100",12651 => "10101100",12652 => "00110111",12653 => "11111111",12654 => "11100000",12655 => "00000011",12656 => "01001100",12657 => "00010101",12658 => "10000110",12659 => "00100101",12660 => "11010000",12661 => "10011111",12662 => "00010101",12663 => "11001111",12664 => "10011110",12665 => "10100101",12666 => "10011010",12667 => "11111111",12668 => "11001110",12669 => "00011010",12670 => "01100011",12671 => "00001101",12672 => "10100100",12673 => "10100001",12674 => "10011110",12675 => "11011110",12676 => "01000100",12677 => "00011111",12678 => "11010000",12679 => "00110110",12680 => "10001010",12681 => "00000110",12682 => "10100001",12683 => "01001010",12684 => "00110100",12685 => "01000011",12686 => "11000001",12687 => "10011100",12688 => "10011011",12689 => "01010110",12690 => "00011011",12691 => "10101001",12692 => "00001010",12693 => "10101111",12694 => "11100010",12695 => "00011110",12696 => "10000100",12697 => "11110111",12698 => "10010100",12699 => "00111100",12700 => "01111111",12701 => "11111111",12702 => "10111101",12703 => "01111010",12704 => "10011011",12705 => "00000111",12706 => "00000110",12707 => "10111111",12708 => "10110001",12709 => "11011010",12710 => "11101000",12711 => "01010010",12712 => "00000000",12713 => "01000100",12714 => "11110110",12715 => "00101010",12716 => "11111110",12717 => "00110010",12718 => "11110011",12719 => "01011110",12720 => "00001010",12721 => "01000110",12722 => "11110110",12723 => "10010101",12724 => "01001100",12725 => "01011011",12726 => "00000001",12727 => "10001111",12728 => "11101110",12729 => "10101100",12730 => "11000101",12731 => "00000111",12732 => "00010001",12733 => "10111101",12734 => "11111101",12735 => "10101001",12736 => "00001110",12737 => "00011011",12738 => "00001010",12739 => "01110100",12740 => "11110010",12741 => "11000100",12742 => "11000001",12743 => "11100100",12744 => "01011001",12745 => "11110100",12746 => "00001011",12747 => "00010100",12748 => "00101010",12749 => "00110100",12750 => "01000010",12751 => "10001010",12752 => "11110110",12753 => "10011100",12754 => "11011111",12755 => "11100110",12756 => "11110011",12757 => "10001111",12758 => "11111100",12759 => "01110111",12760 => "00001010",12761 => "11110010",12762 => "11110000",12763 => "11011101",12764 => "01011110",12765 => "01111011",12766 => "11001001",12767 => "00110111",12768 => "11100111",12769 => "01010000",12770 => "01001110",12771 => "01101000",12772 => "00110100",12773 => "10110100",12774 => "01111100",12775 => "11110100",12776 => "00011010",12777 => "10100000",12778 => "11101101",12779 => "10001110",12780 => "10001011",12781 => "00001100",12782 => "10001000",12783 => "11101010",12784 => "00001000",12785 => "11101011",12786 => "10101011",12787 => "10101101",12788 => "10101101",12789 => "10111001",12790 => "00111111",12791 => "11101111",12792 => "00010101",12793 => "10111000",12794 => "01110000",12795 => "11000010",12796 => "10011011",12797 => "01101000",12798 => "11110001",12799 => "00001100",12800 => "00101111",12801 => "01010110",12802 => "10000000",12803 => "01011000",12804 => "10110111",12805 => "00000110",12806 => "00101101",12807 => "10000101",12808 => "11010101",12809 => "01010000",12810 => "00011100",12811 => "00110010",12812 => "01100000",12813 => "00000101",12814 => "00000101",12815 => "01011111",12816 => "10101000",12817 => "11010101",12818 => "10001000",12819 => "00001111",12820 => "11100001",12821 => "01010101",12822 => "11011101",12823 => "10101111",12824 => "01000010",12825 => "10111111",12826 => "10100101",12827 => "10010101",12828 => "01001000",12829 => "11001010",12830 => "01110100",12831 => "00100000",12832 => "00011001",12833 => "11111110",12834 => "10011100",12835 => "01101001",12836 => "11110101",12837 => "10011111",12838 => "11011010",12839 => "11111011",12840 => "10101000",12841 => "11100000",12842 => "01001001",12843 => "01101111",12844 => "10000011",12845 => "10110110",12846 => "00111000",12847 => "01100111",12848 => "10110111",12849 => "00000110",12850 => "10110001",12851 => "01001011",12852 => "11011111",12853 => "11010010",12854 => "10011000",12855 => "10111110",12856 => "01010001",12857 => "10010010",12858 => "10111010",12859 => "01010011",12860 => "10010101",12861 => "11000101",12862 => "11011101",12863 => "01000100",12864 => "10110010",12865 => "00110001",12866 => "11000010",12867 => "00111011",12868 => "11000001",12869 => "00001110",12870 => "00110101",12871 => "11101101",12872 => "11001001",12873 => "00110011",12874 => "11000111",12875 => "01010101",12876 => "11001011",12877 => "01111010",12878 => "00010001",12879 => "01000110",12880 => "10100000",12881 => "11110100",12882 => "01001110",12883 => "00101011",12884 => "10010001",12885 => "00111100",12886 => "11001100",12887 => "00001010",12888 => "00101011",12889 => "11110101",12890 => "00101001",12891 => "01000110",12892 => "10010101",12893 => "00111010",12894 => "00101010",12895 => "11010110",12896 => "10111111",12897 => "11001001",12898 => "10011110",12899 => "11000110",12900 => "01100001",12901 => "11001010",12902 => "01111100",12903 => "01111010",12904 => "11000010",12905 => "10101010",12906 => "11111101",12907 => "10110000",12908 => "10110111",12909 => "11000100",12910 => "01101010",12911 => "00011101",12912 => "00100100",12913 => "10001110",12914 => "11111110",12915 => "00010111",12916 => "00001011",12917 => "10111011",12918 => "11111101",12919 => "11111010",12920 => "10010010",12921 => "10110000",12922 => "11010011",12923 => "10101000",12924 => "01100101",12925 => "00111000",12926 => "00101100",12927 => "10100101",12928 => "11001010",12929 => "11111110",12930 => "10001000",12931 => "00110011",12932 => "11100110",12933 => "11101001",12934 => "00001111",12935 => "01010100",12936 => "00001110",12937 => "10110101",12938 => "11001010",12939 => "10101011",12940 => "10111011",12941 => "00110000",12942 => "11100011",12943 => "00010010",12944 => "11001011",12945 => "10000011",12946 => "01111111",12947 => "00111101",12948 => "01101110",12949 => "01111110",12950 => "01011000",12951 => "10001110",12952 => "10000110",12953 => "00101011",12954 => "00111111",12955 => "00001100",12956 => "10101011",12957 => "01111000",12958 => "11111010",12959 => "11011100",12960 => "01000101",12961 => "00010000",12962 => "10010110",12963 => "11010101",12964 => "00111001",12965 => "11100101",12966 => "01001110",12967 => "01100010",12968 => "00000111",12969 => "10001000",12970 => "10001100",12971 => "10101001",12972 => "10100010",12973 => "00001101",12974 => "11101110",12975 => "10011010",12976 => "10000001",12977 => "10010110",12978 => "11111100",12979 => "11011110",12980 => "10101101",12981 => "01011100",12982 => "11011001",12983 => "10001100",12984 => "01111100",12985 => "10101000",12986 => "01111001",12987 => "11010011",12988 => "10110011",12989 => "11001010",12990 => "01011100",12991 => "01100100",12992 => "01011000",12993 => "00110011",12994 => "11000111",12995 => "00101011",12996 => "11001000",12997 => "00110011",12998 => "11111011",12999 => "00010010",13000 => "00111111",13001 => "00000010",13002 => "11100010",13003 => "00010101",13004 => "00101101",13005 => "10111010",13006 => "01110000",13007 => "01011011",13008 => "00101000",13009 => "11110111",13010 => "01011001",13011 => "00001100",13012 => "01010000",13013 => "00001111",13014 => "11110101",13015 => "10101101",13016 => "10000001",13017 => "00010100",13018 => "01101011",13019 => "11000010",13020 => "00111010",13021 => "10110010",13022 => "10100111",13023 => "10110100",13024 => "00001100",13025 => "10100001",13026 => "11101111",13027 => "11100011",13028 => "00000101",13029 => "11111111",13030 => "01010100",13031 => "00100010",13032 => "11001111",13033 => "00010111",13034 => "10000010",13035 => "00100000",13036 => "01110110",13037 => "11000011",13038 => "01011010",13039 => "10010111",13040 => "10001010",13041 => "01110110",13042 => "01000100",13043 => "00111111",13044 => "01110001",13045 => "10111111",13046 => "10100111",13047 => "10000011",13048 => "01101110",13049 => "01001101",13050 => "01101011",13051 => "11010111",13052 => "10000010",13053 => "10001101",13054 => "00100000",13055 => "10111000",13056 => "00001110",13057 => "01110110",13058 => "01101110",13059 => "00111101",13060 => "00101111",13061 => "01101100",13062 => "00100000",13063 => "11011011",13064 => "00001110",13065 => "11110010",13066 => "10000100",13067 => "00011111",13068 => "11001011",13069 => "10111110",13070 => "10010001",13071 => "10111000",13072 => "00000110",13073 => "10000100",13074 => "11010100",13075 => "01100101",13076 => "01010000",13077 => "10010010",13078 => "00000100",13079 => "11110000",13080 => "11010011",13081 => "11111010",13082 => "10110010",13083 => "00110100",13084 => "01000001",13085 => "11010101",13086 => "11011101",13087 => "01111110",13088 => "10010111",13089 => "01010010",13090 => "10110100",13091 => "10101101",13092 => "00111111",13093 => "00110000",13094 => "10101111",13095 => "00111011",13096 => "00110111",13097 => "00010110",13098 => "01011010",13099 => "10100001",13100 => "11110111",13101 => "01011001",13102 => "01100101",13103 => "01011101",13104 => "01110000",13105 => "01110111",13106 => "00110011",13107 => "01011100",13108 => "00001101",13109 => "01011001",13110 => "00010110",13111 => "01110011",13112 => "10100110",13113 => "11011011",13114 => "01001001",13115 => "01001010",13116 => "01111101",13117 => "10011101",13118 => "00011110",13119 => "11010111",13120 => "11100010",13121 => "01111010",13122 => "11110110",13123 => "10110100",13124 => "00111000",13125 => "11011001",13126 => "10000010",13127 => "01011111",13128 => "00001001",13129 => "11000010",13130 => "10011111",13131 => "11001100",13132 => "01001101",13133 => "11010010",13134 => "00100100",13135 => "10001110",13136 => "10001101",13137 => "00011100",13138 => "01111111",13139 => "01011100",13140 => "01011001",13141 => "11111011",13142 => "01101000",13143 => "00011100",13144 => "11100101",13145 => "11101101",13146 => "11010100",13147 => "00000111",13148 => "01100110",13149 => "01101111",13150 => "10000111",13151 => "11011010",13152 => "10010101",13153 => "00101110",13154 => "11110100",13155 => "01111011",13156 => "00000010",13157 => "10000110",13158 => "00110101",13159 => "11011000",13160 => "11111011",13161 => "00100101",13162 => "01010000",13163 => "10111011",13164 => "11001111",13165 => "10011101",13166 => "01001001",13167 => "11000100",13168 => "11100101",13169 => "01010000",13170 => "01001100",13171 => "01000010",13172 => "10001010",13173 => "00000111",13174 => "01001101",13175 => "00001000",13176 => "01110100",13177 => "11111000",13178 => "00010100",13179 => "11100011",13180 => "01110010",13181 => "01100100",13182 => "01000100",13183 => "11001100",13184 => "00101101",13185 => "10011011",13186 => "11101100",13187 => "01111011",13188 => "01111101",13189 => "10010011",13190 => "10111110",13191 => "01101101",13192 => "11100011",13193 => "11001101",13194 => "00010011",13195 => "01001110",13196 => "00010101",13197 => "01010001",13198 => "01111010",13199 => "11001110",13200 => "01100000",13201 => "11100110",13202 => "11001111",13203 => "11101100",13204 => "00001101",13205 => "10000111",13206 => "00110111",13207 => "11000100",13208 => "11011110",13209 => "10100100",13210 => "00000001",13211 => "10010111",13212 => "00110100",13213 => "01000011",13214 => "01001110",13215 => "01101010",13216 => "01001010",13217 => "00000100",13218 => "10010010",13219 => "00010011",13220 => "11010000",13221 => "11010001",13222 => "00111010",13223 => "11100010",13224 => "00011001",13225 => "11000001",13226 => "11001010",13227 => "11010110",13228 => "00110010",13229 => "00010010",13230 => "11111110",13231 => "00010111",13232 => "10000111",13233 => "00110011",13234 => "01000110",13235 => "00110000",13236 => "11011101",13237 => "01001000",13238 => "10011111",13239 => "10010010",13240 => "01010011",13241 => "10110011",13242 => "11000011",13243 => "11001001",13244 => "01111111",13245 => "00000111",13246 => "10110111",13247 => "11111010",13248 => "01101111",13249 => "11011110",13250 => "00000101",13251 => "01000011",13252 => "01011001",13253 => "00000011",13254 => "00000000",13255 => "01000100",13256 => "10110101",13257 => "00001101",13258 => "10111111",13259 => "01101010",13260 => "11101000",13261 => "01001010",13262 => "11110111",13263 => "01001101",13264 => "10011100",13265 => "00101011",13266 => "00010110",13267 => "11010000",13268 => "01111011",13269 => "11101000",13270 => "11010100",13271 => "11100000",13272 => "00100111",13273 => "11001111",13274 => "01011111",13275 => "11001011",13276 => "10110001",13277 => "01110110",13278 => "01101011",13279 => "01011111",13280 => "10011010",13281 => "01011101",13282 => "10111101",13283 => "01101001",13284 => "00100011",13285 => "10001110",13286 => "00000000",13287 => "01110001",13288 => "10011000",13289 => "10010011",13290 => "10110010",13291 => "10110001",13292 => "11000110",13293 => "11100001",13294 => "00010010",13295 => "10001010",13296 => "10111001",13297 => "00111000",13298 => "01100010",13299 => "01100001",13300 => "10101001",13301 => "00100111",13302 => "00110100",13303 => "11101111",13304 => "00001011",13305 => "00100000",13306 => "11011001",13307 => "01010000",13308 => "11010000",13309 => "00100101",13310 => "11001111",13311 => "11110010",13312 => "01010111",13313 => "11101000",13314 => "10010001",13315 => "10110010",13316 => "10101001",13317 => "01110000",13318 => "00000111",13319 => "10111001",13320 => "10011011",13321 => "01100110",13322 => "11000111",13323 => "10110110",13324 => "10000111",13325 => "10011110",13326 => "00010000",13327 => "11000110",13328 => "10100110",13329 => "11000101",13330 => "01111101",13331 => "00100001",13332 => "00100101",13333 => "01010001",13334 => "00110110",13335 => "11001000",13336 => "00001001",13337 => "00010011",13338 => "11000100",13339 => "00100000",13340 => "11100111",13341 => "10111101",13342 => "00001011",13343 => "10100010",13344 => "00111101",13345 => "01010000",13346 => "01111010",13347 => "01101010",13348 => "10110001",13349 => "11000111",13350 => "00010010",13351 => "11010010",13352 => "10100011",13353 => "10100110",13354 => "11011000",13355 => "01111110",13356 => "10010110",13357 => "11100010",13358 => "11011100",13359 => "00000011",13360 => "11111011",13361 => "00001001",13362 => "00101011",13363 => "10110111",13364 => "00000010",13365 => "01101111",13366 => "10101000",13367 => "10101110",13368 => "11101100",13369 => "11011110",13370 => "10001000",13371 => "00011100",13372 => "10100101",13373 => "00110011",13374 => "01010001",13375 => "10011001",13376 => "00001001",13377 => "10111100",13378 => "00010100",13379 => "10010100",13380 => "10101101",13381 => "11000100",13382 => "00011010",13383 => "01100100",13384 => "00011000",13385 => "11010101",13386 => "00010011",13387 => "11011101",13388 => "00111101",13389 => "11010000",13390 => "11001011",13391 => "10011100",13392 => "10000101",13393 => "00100010",13394 => "10111001",13395 => "11100001",13396 => "01110100",13397 => "01111100",13398 => "00000100",13399 => "00100001",13400 => "10100110",13401 => "00000110",13402 => "11010000",13403 => "00111110",13404 => "11011110",13405 => "01001100",13406 => "00011000",13407 => "01011101",13408 => "11100111",13409 => "11111000",13410 => "10001011",13411 => "01111010",13412 => "11101001",13413 => "00011010",13414 => "00001111",13415 => "11000010",13416 => "11011000",13417 => "10111101",13418 => "10010101",13419 => "00000100",13420 => "10011010",13421 => "01010010",13422 => "01101011",13423 => "10111010",13424 => "00110110",13425 => "10101001",13426 => "01101010",13427 => "10111001",13428 => "00011001",13429 => "00111110",13430 => "01001001",13431 => "01100011",13432 => "00110010",13433 => "11101000",13434 => "00111101",13435 => "00000000",13436 => "01101010",13437 => "11101000",13438 => "00000000",13439 => "11111001",13440 => "01000000",13441 => "00110000",13442 => "00101101",13443 => "01000101",13444 => "00001100",13445 => "00010011",13446 => "00011011",13447 => "11001101",13448 => "01101111",13449 => "00100111",13450 => "11000011",13451 => "00111001",13452 => "11111100",13453 => "11110010",13454 => "01111100",13455 => "10111011",13456 => "11111000",13457 => "00010010",13458 => "11001110",13459 => "00000100",13460 => "11110110",13461 => "01010100",13462 => "10010101",13463 => "01111100",13464 => "00011011",13465 => "01010100",13466 => "11011100",13467 => "01010001",13468 => "01100010",13469 => "10011001",13470 => "10001100",13471 => "00100101",13472 => "11010101",13473 => "01101101",13474 => "10111111",13475 => "11111100",13476 => "10000000",13477 => "11000100",13478 => "00011111",13479 => "10001011",13480 => "11110100",13481 => "10100000",13482 => "00100101",13483 => "11011010",13484 => "11100001",13485 => "00101110",13486 => "11101110",13487 => "10011001",13488 => "10000010",13489 => "11100111",13490 => "00011011",13491 => "11100001",13492 => "00011101",13493 => "01010010",13494 => "01010011",13495 => "01111001",13496 => "00001101",13497 => "11001100",13498 => "01000111",13499 => "00100010",13500 => "10010110",13501 => "11001000",13502 => "01001011",13503 => "11110100",13504 => "11110110",13505 => "10100011",13506 => "11000001",13507 => "01100110",13508 => "01110010",13509 => "01011100",13510 => "11100010",13511 => "10001000",13512 => "10010001",13513 => "10100100",13514 => "10000000",13515 => "11100000",13516 => "00110000",13517 => "00110110",13518 => "00110011",13519 => "11101001",13520 => "10001101",13521 => "00011101",13522 => "10011101",13523 => "11010000",13524 => "11001000",13525 => "10001100",13526 => "01011001",13527 => "00011100",13528 => "00010110",13529 => "10001101",13530 => "01111100",13531 => "01110001",13532 => "10011000",13533 => "01010101",13534 => "10001010",13535 => "01111001",13536 => "01111100",13537 => "10111111",13538 => "01111001",13539 => "10100110",13540 => "10100110",13541 => "10000111",13542 => "00100011",13543 => "10100011",13544 => "01000011",13545 => "11111100",13546 => "01001000",13547 => "11110000",13548 => "01001001",13549 => "00111110",13550 => "11011100",13551 => "00111000",13552 => "01101000",13553 => "10100101",13554 => "01000111",13555 => "01110100",13556 => "00001110",13557 => "01100001",13558 => "00111110",13559 => "10111100",13560 => "11011100",13561 => "01110001",13562 => "10100111",13563 => "11010010",13564 => "11110010",13565 => "00010001",13566 => "10111000",13567 => "01111101",13568 => "10110101",13569 => "10100101",13570 => "11000101",13571 => "10110101",13572 => "11101011",13573 => "00100111",13574 => "01011010",13575 => "01100111",13576 => "10000100",13577 => "10000010",13578 => "11111010",13579 => "10000001",13580 => "11010001",13581 => "10111011",13582 => "10011101",13583 => "11100001",13584 => "00001010",13585 => "00001101",13586 => "10110110",13587 => "10000010",13588 => "11001110",13589 => "11011111",13590 => "11110011",13591 => "11011000",13592 => "11100110",13593 => "10011101",13594 => "11100111",13595 => "00101100",13596 => "11011010",13597 => "00110011",13598 => "01001101",13599 => "10000001",13600 => "00111110",13601 => "11101110",13602 => "11101100",13603 => "11000101",13604 => "11100100",13605 => "10111001",13606 => "00110100",13607 => "11101111",13608 => "10110000",13609 => "01101101",13610 => "00110001",13611 => "10011100",13612 => "10000001",13613 => "10101001",13614 => "10100110",13615 => "01001001",13616 => "01110111",13617 => "11010000",13618 => "10111101",13619 => "00011001",13620 => "01011000",13621 => "10010010",13622 => "10010011",13623 => "10010101",13624 => "11101110",13625 => "00010110",13626 => "00011100",13627 => "11110100",13628 => "10011101",13629 => "00010001",13630 => "00101011",13631 => "01000010",13632 => "01011101",13633 => "10010111",13634 => "11010001",13635 => "01011000",13636 => "10110000",13637 => "01011101",13638 => "00100011",13639 => "00100010",13640 => "01110110",13641 => "10100011",13642 => "01101111",13643 => "01000000",13644 => "10101101",13645 => "00010000",13646 => "01000000",13647 => "11011000",13648 => "01011010",13649 => "01111001",13650 => "10110110",13651 => "01101101",13652 => "01101101",13653 => "10010000",13654 => "01101101",13655 => "10101101",13656 => "11100100",13657 => "01001110",13658 => "01101010",13659 => "10001111",13660 => "01001011",13661 => "01001111",13662 => "00001101",13663 => "01100010",13664 => "11100111",13665 => "01001011",13666 => "11100100",13667 => "10011001",13668 => "01011100",13669 => "01000110",13670 => "01001100",13671 => "01100011",13672 => "11011011",13673 => "00100100",13674 => "00111000",13675 => "10011100",13676 => "01111000",13677 => "10111100",13678 => "00101010",13679 => "10110001",13680 => "00100011",13681 => "01010111",13682 => "10111000",13683 => "11011010",13684 => "00010110",13685 => "11010010",13686 => "01000000",13687 => "10110000",13688 => "00101100",13689 => "11110010",13690 => "00010100",13691 => "11011110",13692 => "10011110",13693 => "01011010",13694 => "01100101",13695 => "00101100",13696 => "10011000",13697 => "00010010",13698 => "00001001",13699 => "01100000",13700 => "01001111",13701 => "00110100",13702 => "00010100",13703 => "01101010",13704 => "11101101",13705 => "01110001",13706 => "01010100",13707 => "10101011",13708 => "10000010",13709 => "01011110",13710 => "01110101",13711 => "00011111",13712 => "11011101",13713 => "00011101",13714 => "11111100",13715 => "00001100",13716 => "10101011",13717 => "11101001",13718 => "11111100",13719 => "10010110",13720 => "00110011",13721 => "10110100",13722 => "10010010",13723 => "10111101",13724 => "10011100",13725 => "00000111",13726 => "11101000",13727 => "00000100",13728 => "10100100",13729 => "10110011",13730 => "01000101",13731 => "00110110",13732 => "10111101",13733 => "10010001",13734 => "10101000",13735 => "01011011",13736 => "00010101",13737 => "11110100",13738 => "11101100",13739 => "10011110",13740 => "01111001",13741 => "11000100",13742 => "00001110",13743 => "01011110",13744 => "01011010",13745 => "01111001",13746 => "11100110",13747 => "01010000",13748 => "11010111",13749 => "11001110",13750 => "11000100",13751 => "10000010",13752 => "10101001",13753 => "10100000",13754 => "10111010",13755 => "11010101",13756 => "10110111",13757 => "00111100",13758 => "11111110",13759 => "10011010",13760 => "01001010",13761 => "11111001",13762 => "00000010",13763 => "01000111",13764 => "00011010",13765 => "11011011",13766 => "01000011",13767 => "01101010",13768 => "00011101",13769 => "11100100",13770 => "01010100",13771 => "01101010",13772 => "00001010",13773 => "01100101",13774 => "01110011",13775 => "10011101",13776 => "01001101",13777 => "10011011",13778 => "01101100",13779 => "00100100",13780 => "00100011",13781 => "00110011",13782 => "00110010",13783 => "11100001",13784 => "01100010",13785 => "10010001",13786 => "10110011",13787 => "00111011",13788 => "11110010",13789 => "10010010",13790 => "11100100",13791 => "00111001",13792 => "10000010",13793 => "11001001",13794 => "01101111",13795 => "11111101",13796 => "10001011",13797 => "00000010",13798 => "11001101",13799 => "01100101",13800 => "00101010",13801 => "11000010",13802 => "00111000",13803 => "10010101",13804 => "01000010",13805 => "11000111",13806 => "01110000",13807 => "11111111",13808 => "10001111",13809 => "00111001",13810 => "11110011",13811 => "10010101",13812 => "10101010",13813 => "10100111",13814 => "00011011",13815 => "11001111",13816 => "10000010",13817 => "11111000",13818 => "10111010",13819 => "11110001",13820 => "10110110",13821 => "11111011",13822 => "00000110",13823 => "11001011",13824 => "01110100",13825 => "11111000",13826 => "11011111",13827 => "10000101",13828 => "00101110",13829 => "10000000",13830 => "00100011",13831 => "01100011",13832 => "10100110",13833 => "11001000",13834 => "11110101",13835 => "01001111",13836 => "01101011",13837 => "10010010",13838 => "11000111",13839 => "00110001",13840 => "00101011",13841 => "00000100",13842 => "11111010",13843 => "01110101",13844 => "01101100",13845 => "00101000",13846 => "11001111",13847 => "10110111",13848 => "00010101",13849 => "11111010",13850 => "00101110",13851 => "00000010",13852 => "01000110",13853 => "00100011",13854 => "11000011",13855 => "11101000",13856 => "00111000",13857 => "10010101",13858 => "01101110",13859 => "01001011",13860 => "10010100",13861 => "00001010",13862 => "00000011",13863 => "10001011",13864 => "00000111",13865 => "01110001",13866 => "11100010",13867 => "01001001",13868 => "01111100",13869 => "11011010",13870 => "01000001",13871 => "01101100",13872 => "00101110",13873 => "10110110",13874 => "11000010",13875 => "11110111",13876 => "01011000",13877 => "00011110",13878 => "10000011",13879 => "01111111",13880 => "00010011",13881 => "10010101",13882 => "00101001",13883 => "11101010",13884 => "01110101",13885 => "10100000",13886 => "01001101",13887 => "10001110",13888 => "00010100",13889 => "01111010",13890 => "01011100",13891 => "10101111",13892 => "00011111",13893 => "00000011",13894 => "00000000",13895 => "00110001",13896 => "11010111",13897 => "10011011",13898 => "01000110",13899 => "00011101",13900 => "01100101",13901 => "11011010",13902 => "00011100",13903 => "01011101",13904 => "01010011",13905 => "10110101",13906 => "00110011",13907 => "00000001",13908 => "10101110",13909 => "11101010",13910 => "01001001",13911 => "01111010",13912 => "10111010",13913 => "00111111",13914 => "01001101",13915 => "01111011",13916 => "10101101",13917 => "10011000",13918 => "10101001",13919 => "01011101",13920 => "10001100",13921 => "01100111",13922 => "11011110",13923 => "00010010",13924 => "10100110",13925 => "10101001",13926 => "00110000",13927 => "11010111",13928 => "10101100",13929 => "00010101",13930 => "00010101",13931 => "01010010",13932 => "10100001",13933 => "00010000",13934 => "00011001",13935 => "01010011",13936 => "01010100",13937 => "11001011",13938 => "10001010",13939 => "00001111",13940 => "01000000",13941 => "11110101",13942 => "01101100",13943 => "11111010",13944 => "00011001",13945 => "11110100",13946 => "01111111",13947 => "01001110",13948 => "10010110",13949 => "01100010",13950 => "00110010",13951 => "10111000",13952 => "10011001",13953 => "10010100",13954 => "00100010",13955 => "00110000",13956 => "10101101",13957 => "10001010",13958 => "00000001",13959 => "00110011",13960 => "01101110",13961 => "01011100",13962 => "00011110",13963 => "00001110",13964 => "01011001",13965 => "01101101",13966 => "11001001",13967 => "11101100",13968 => "01010101",13969 => "10101100",13970 => "01100100",13971 => "00110011",13972 => "00010000",13973 => "00001010",13974 => "01000110",13975 => "10111100",13976 => "01011101",13977 => "00010110",13978 => "11101010",13979 => "11010101",13980 => "01111000",13981 => "10000011",13982 => "10010011",13983 => "00110001",13984 => "11111010",13985 => "01001110",13986 => "01111110",13987 => "11100110",13988 => "01010110",13989 => "11001011",13990 => "00110011",13991 => "01100001",13992 => "00111010",13993 => "01110001",13994 => "00001010",13995 => "11111011",13996 => "10010010",13997 => "10000111",13998 => "00000101",13999 => "10100000",14000 => "11001010",14001 => "10000000",14002 => "00010110",14003 => "01011100",14004 => "10000111",14005 => "10000100",14006 => "00100100",14007 => "10010110",14008 => "11111000",14009 => "10010000",14010 => "00100001",14011 => "00001100",14012 => "11001000",14013 => "10101110",14014 => "00101101",14015 => "01011110",14016 => "10000001",14017 => "00011110",14018 => "00111000",14019 => "11011100",14020 => "11101111",14021 => "11110000",14022 => "11010100",14023 => "01101000",14024 => "01110110",14025 => "11100011",14026 => "00001111",14027 => "11100010",14028 => "10010001",14029 => "00100000",14030 => "10001110",14031 => "00110101",14032 => "00010010",14033 => "01101001",14034 => "00110000",14035 => "00100100",14036 => "00011001",14037 => "01101100",14038 => "10000100",14039 => "11101111",14040 => "00001010",14041 => "01111011",14042 => "00001000",14043 => "10001110",14044 => "01111101",14045 => "00010110",14046 => "11010011",14047 => "01111100",14048 => "11010001",14049 => "10110110",14050 => "10111000",14051 => "01001101",14052 => "10001101",14053 => "01111110",14054 => "01111111",14055 => "01100111",14056 => "00011100",14057 => "10000000",14058 => "00000100",14059 => "01010001",14060 => "00000010",14061 => "11011111",14062 => "01110110",14063 => "00001101",14064 => "01010011",14065 => "11110011",14066 => "10010011",14067 => "01100010",14068 => "01111000",14069 => "11000101",14070 => "10000100",14071 => "01000010",14072 => "01111001",14073 => "00111101",14074 => "01110001",14075 => "00110100",14076 => "00110110",14077 => "01010100",14078 => "00011000",14079 => "10010101",14080 => "11101011",14081 => "11111100",14082 => "10000010",14083 => "01001110",14084 => "01110000",14085 => "00100101",14086 => "01010100",14087 => "00011101",14088 => "11101011",14089 => "10110101",14090 => "11001001",14091 => "00101101",14092 => "01010000",14093 => "11001100",14094 => "10111100",14095 => "00011001",14096 => "10100001",14097 => "01101001",14098 => "01000100",14099 => "11010001",14100 => "11101101",14101 => "10110010",14102 => "10110010",14103 => "01011111",14104 => "10010011",14105 => "10010110",14106 => "00101010",14107 => "00011111",14108 => "00111010",14109 => "11011001",14110 => "10010101",14111 => "00001101",14112 => "10010001",14113 => "00000010",14114 => "11101101",14115 => "01010011",14116 => "00110110",14117 => "00100001",14118 => "01000000",14119 => "01011101",14120 => "01101110",14121 => "01000101",14122 => "10001100",14123 => "10110010",14124 => "00100101",14125 => "10101010",14126 => "10000011",14127 => "01111000",14128 => "00110101",14129 => "11011001",14130 => "01001100",14131 => "11001011",14132 => "00111000",14133 => "11101111",14134 => "10011000",14135 => "10111011",14136 => "10100010",14137 => "01011110",14138 => "00011100",14139 => "01010111",14140 => "10010111",14141 => "11111110",14142 => "01001111",14143 => "11000101",14144 => "01001110",14145 => "10011011",14146 => "11101010",14147 => "00110111",14148 => "11111110",14149 => "01111010",14150 => "00110101",14151 => "10101110",14152 => "11100010",14153 => "00000000",14154 => "00110010",14155 => "11001101",14156 => "01111000",14157 => "10000001",14158 => "11100000",14159 => "10011101",14160 => "10011001",14161 => "00011111",14162 => "00100110",14163 => "00001111",14164 => "01000100",14165 => "00010101",14166 => "01110110",14167 => "01010011",14168 => "01000011",14169 => "00111111",14170 => "10000011",14171 => "00000100",14172 => "01100111",14173 => "00001010",14174 => "10100101",14175 => "00011110",14176 => "10001001",14177 => "10000110",14178 => "00000000",14179 => "10011000",14180 => "01110011",14181 => "11110001",14182 => "10011101",14183 => "10110111",14184 => "00100010",14185 => "11010011",14186 => "11111000",14187 => "00110110",14188 => "11111110",14189 => "11111111",14190 => "11101010",14191 => "01001000",14192 => "01110000",14193 => "00101000",14194 => "00011010",14195 => "01101001",14196 => "01001111",14197 => "01011110",14198 => "00100001",14199 => "00101011",14200 => "01010101",14201 => "11001110",14202 => "11100111",14203 => "10011101",14204 => "01000000",14205 => "01100000",14206 => "10010001",14207 => "10101001",14208 => "11001110",14209 => "10000011",14210 => "10011011",14211 => "00010001",14212 => "11010110",14213 => "10100100",14214 => "10100111",14215 => "11100110",14216 => "00101001",14217 => "01110011",14218 => "11000111",14219 => "00011011",14220 => "01010010",14221 => "00101000",14222 => "11011011",14223 => "00011011",14224 => "11101111",14225 => "11110000",14226 => "11101011",14227 => "01111001",14228 => "11000101",14229 => "10001111",14230 => "11110100",14231 => "11001001",14232 => "10111111",14233 => "11100001",14234 => "11000001",14235 => "11000100",14236 => "01110100",14237 => "11010101",14238 => "01010011",14239 => "10011110",14240 => "01010111",14241 => "01101101",14242 => "00001100",14243 => "11000111",14244 => "00110011",14245 => "01111111",14246 => "10110110",14247 => "01010011",14248 => "01010111",14249 => "10010011",14250 => "00101100",14251 => "00110011",14252 => "00010001",14253 => "10010001",14254 => "01001111",14255 => "11100111",14256 => "01111111",14257 => "01100000",14258 => "00000101",14259 => "11101011",14260 => "10010111",14261 => "10101110",14262 => "11010110",14263 => "11101000",14264 => "01101111",14265 => "10101001",14266 => "11101111",14267 => "01010100",14268 => "01011011",14269 => "00000011",14270 => "11100111",14271 => "10001110",14272 => "10010000",14273 => "10001100",14274 => "01111101",14275 => "01111101",14276 => "10011100",14277 => "11101010",14278 => "01100111",14279 => "11101011",14280 => "00111001",14281 => "10001111",14282 => "11010010",14283 => "11001100",14284 => "10010000",14285 => "11111101",14286 => "01100110",14287 => "11111100",14288 => "01110101",14289 => "11100110",14290 => "00100010",14291 => "11111100",14292 => "10100011",14293 => "00100000",14294 => "00111101",14295 => "00010000",14296 => "10001011",14297 => "10011001",14298 => "11011100",14299 => "10101010",14300 => "11010000",14301 => "11011101",14302 => "00000011",14303 => "00101100",14304 => "10101000",14305 => "01100000",14306 => "01110111",14307 => "00100001",14308 => "00101110",14309 => "01000111",14310 => "01101011",14311 => "11000010",14312 => "11010001",14313 => "10101010",14314 => "00100100",14315 => "00111000",14316 => "01000110",14317 => "01111100",14318 => "10100010",14319 => "10110000",14320 => "11010001",14321 => "11011011",14322 => "00101001",14323 => "10000010",14324 => "11010010",14325 => "10101001",14326 => "11010100",14327 => "10010001",14328 => "11111110",14329 => "01101001",14330 => "11001111",14331 => "01001011",14332 => "11110101",14333 => "11110110",14334 => "10001010",14335 => "00000010",14336 => "01101110",14337 => "10000110",14338 => "01011001",14339 => "00011101",14340 => "10111100",14341 => "10100000",14342 => "01010101",14343 => "11101100",14344 => "00011110",14345 => "01101010",14346 => "01110110",14347 => "01000101",14348 => "01010001",14349 => "01001100",14350 => "01110000",14351 => "00001001",14352 => "10101000",14353 => "01001101",14354 => "01010010",14355 => "01100010",14356 => "10101101",14357 => "11101100",14358 => "11001100",14359 => "11001011",14360 => "00100000",14361 => "11101011",14362 => "00010011",14363 => "11100100",14364 => "00110101",14365 => "00110110",14366 => "10111100",14367 => "11010101",14368 => "11101011",14369 => "01011100",14370 => "01100010",14371 => "11111011",14372 => "01110100",14373 => "01110100",14374 => "01011101",14375 => "01010000",14376 => "11110100",14377 => "10101110",14378 => "01100001",14379 => "11111010",14380 => "01010100",14381 => "01100000",14382 => "10110010",14383 => "01010000",14384 => "01111010",14385 => "10100011",14386 => "10001100",14387 => "01101111",14388 => "11000011",14389 => "01011011",14390 => "10010000",14391 => "10001110",14392 => "01011110",14393 => "10110111",14394 => "01011110",14395 => "01001110",14396 => "10011100",14397 => "10011010",14398 => "10010100",14399 => "10100010",14400 => "00010100",14401 => "11110000",14402 => "01001100",14403 => "11101110",14404 => "10011100",14405 => "11000100",14406 => "10100001",14407 => "01101001",14408 => "10010100",14409 => "01000110",14410 => "00010011",14411 => "00000001",14412 => "11001011",14413 => "01111000",14414 => "01101000",14415 => "11100100",14416 => "10111011",14417 => "11000011",14418 => "10010000",14419 => "10110110",14420 => "00100100",14421 => "01100010",14422 => "01011000",14423 => "00011110",14424 => "01100100",14425 => "10101010",14426 => "10010101",14427 => "00101110",14428 => "10111010",14429 => "00000110",14430 => "10101100",14431 => "10001100",14432 => "10100001",14433 => "00100100",14434 => "11101101",14435 => "11010101",14436 => "01100101",14437 => "00010100",14438 => "00111110",14439 => "10000111",14440 => "01011111",14441 => "01001010",14442 => "11100101",14443 => "00001111",14444 => "01111011",14445 => "01100111",14446 => "11010001",14447 => "01101101",14448 => "11110010",14449 => "10101111",14450 => "10110101",14451 => "00101010",14452 => "10111010",14453 => "00001101",14454 => "10000000",14455 => "11101000",14456 => "11011101",14457 => "01000011",14458 => "01010011",14459 => "10001100",14460 => "00111010",14461 => "01010111",14462 => "00110010",14463 => "10011011",14464 => "10000010",14465 => "00111100",14466 => "10111000",14467 => "00110000",14468 => "10101100",14469 => "10010011",14470 => "11000101",14471 => "11001000",14472 => "01100100",14473 => "01101010",14474 => "00000100",14475 => "10000101",14476 => "10000101",14477 => "10001011",14478 => "00110010",14479 => "00011111",14480 => "10101001",14481 => "00010010",14482 => "00011011",14483 => "00110101",14484 => "10101001",14485 => "11111110",14486 => "01101001",14487 => "11100001",14488 => "00111110",14489 => "11010101",14490 => "10010010",14491 => "00000001",14492 => "01001110",14493 => "11101101",14494 => "01101011",14495 => "01101001",14496 => "11001001",14497 => "10110101",14498 => "01110110",14499 => "11010001",14500 => "10100001",14501 => "01101010",14502 => "00100001",14503 => "01101111",14504 => "11101011",14505 => "01111010",14506 => "10010110",14507 => "01011101",14508 => "10100010",14509 => "01111010",14510 => "11001101",14511 => "10010100",14512 => "01001001",14513 => "00001001",14514 => "01100111",14515 => "01110010",14516 => "01101100",14517 => "10001011",14518 => "00001101",14519 => "01001100",14520 => "01110100",14521 => "01101110",14522 => "01001110",14523 => "10111011",14524 => "11001010",14525 => "01111011",14526 => "10110111",14527 => "11000100",14528 => "01101111",14529 => "00101101",14530 => "01010000",14531 => "10101010",14532 => "01001010",14533 => "10100010",14534 => "10100110",14535 => "11000000",14536 => "01110110",14537 => "01111110",14538 => "00111001",14539 => "11011001",14540 => "10100001",14541 => "10111000",14542 => "11110000",14543 => "10111110",14544 => "00011111",14545 => "11001110",14546 => "01111000",14547 => "00110010",14548 => "01010110",14549 => "00010111",14550 => "10001100",14551 => "10000111",14552 => "01000110",14553 => "00000001",14554 => "11001010",14555 => "00110111",14556 => "01011010",14557 => "00101000",14558 => "01101011",14559 => "11011101",14560 => "00111000",14561 => "10110010",14562 => "00110101",14563 => "11101011",14564 => "11010110",14565 => "00101010",14566 => "01111011",14567 => "00010111",14568 => "01100010",14569 => "00100011",14570 => "11110111",14571 => "10100111",14572 => "11000111",14573 => "01101100",14574 => "01010010",14575 => "00001010",14576 => "10011010",14577 => "11110101",14578 => "00011110",14579 => "01001000",14580 => "10111101",14581 => "01000110",14582 => "11011001",14583 => "00011001",14584 => "10010101",14585 => "01110000",14586 => "11011000",14587 => "10001101",14588 => "01101011",14589 => "11101111",14590 => "01111100",14591 => "00000001",14592 => "11011100",14593 => "10101001",14594 => "10011111",14595 => "00010000",14596 => "10101111",14597 => "00101010",14598 => "00010011",14599 => "11010000",14600 => "10001010",14601 => "10011011",14602 => "10110110",14603 => "00011101",14604 => "10111100",14605 => "10111100",14606 => "00100110",14607 => "10011010",14608 => "11010111",14609 => "11101111",14610 => "00001000",14611 => "01010111",14612 => "00001110",14613 => "00010001",14614 => "00110010",14615 => "11110001",14616 => "11110011",14617 => "11110011",14618 => "00010010",14619 => "00010010",14620 => "10011111",14621 => "00111011",14622 => "01001001",14623 => "00001110",14624 => "10000000",14625 => "10101110",14626 => "11000100",14627 => "00101111",14628 => "00001110",14629 => "11100110",14630 => "10111001",14631 => "01000100",14632 => "00001011",14633 => "11011111",14634 => "00011111",14635 => "10100010",14636 => "01101011",14637 => "11000101",14638 => "00101010",14639 => "10110011",14640 => "00110000",14641 => "10001010",14642 => "11101100",14643 => "01000010",14644 => "00110000",14645 => "11001110",14646 => "10101101",14647 => "00100111",14648 => "00011010",14649 => "01110010",14650 => "00000011",14651 => "10011101",14652 => "01011101",14653 => "00110111",14654 => "11100101",14655 => "10001011",14656 => "00100010",14657 => "00111111",14658 => "10110101",14659 => "01010010",14660 => "10001110",14661 => "10110011",14662 => "01111111",14663 => "11000010",14664 => "01100011",14665 => "01001000",14666 => "11010100",14667 => "00101001",14668 => "10110000",14669 => "10100010",14670 => "01010011",14671 => "00011011",14672 => "00100101",14673 => "01000110",14674 => "01101100",14675 => "01010111",14676 => "10011110",14677 => "11001011",14678 => "10011000",14679 => "00111000",14680 => "11110011",14681 => "00101110",14682 => "11001101",14683 => "10110101",14684 => "10111111",14685 => "01011000",14686 => "00000110",14687 => "10011000",14688 => "00100110",14689 => "10110011",14690 => "11111011",14691 => "11011011",14692 => "10010111",14693 => "00101110",14694 => "01010001",14695 => "01110010",14696 => "01001111",14697 => "10000000",14698 => "00000111",14699 => "11110111",14700 => "10111111",14701 => "01110011",14702 => "00100010",14703 => "11111001",14704 => "11011000",14705 => "11010111",14706 => "01111101",14707 => "01010111",14708 => "01111110",14709 => "10001010",14710 => "00110100",14711 => "10000001",14712 => "01111011",14713 => "01010110",14714 => "10100101",14715 => "01011101",14716 => "10010101",14717 => "10110000",14718 => "00000011",14719 => "10000110",14720 => "00011100",14721 => "00010011",14722 => "01110011",14723 => "01111010",14724 => "11000001",14725 => "01000101",14726 => "01101100",14727 => "00100110",14728 => "10011111",14729 => "01001100",14730 => "10000100",14731 => "00110101",14732 => "00101111",14733 => "10100011",14734 => "10111110",14735 => "10001011",14736 => "01000100",14737 => "10111011",14738 => "10100011",14739 => "11111000",14740 => "11100000",14741 => "01000001",14742 => "10000000",14743 => "00101101",14744 => "01100010",14745 => "10100000",14746 => "11100011",14747 => "01011110",14748 => "01010011",14749 => "10100110",14750 => "11100101",14751 => "11001000",14752 => "11010000",14753 => "00111110",14754 => "11110101",14755 => "00010101",14756 => "10000110",14757 => "11101111",14758 => "10001111",14759 => "10110000",14760 => "01001011",14761 => "01110000",14762 => "01100010",14763 => "11011110",14764 => "10010011",14765 => "10110010",14766 => "11100000",14767 => "01000001",14768 => "10011000",14769 => "10010010",14770 => "10101010",14771 => "11110011",14772 => "11111001",14773 => "10110011",14774 => "00010100",14775 => "00010111",14776 => "00001100",14777 => "01000000",14778 => "10111111",14779 => "10111111",14780 => "01011010",14781 => "10000100",14782 => "11010011",14783 => "00001101",14784 => "10010001",14785 => "00010101",14786 => "11100010",14787 => "00000110",14788 => "00100100",14789 => "10101000",14790 => "00000101",14791 => "10001010",14792 => "01101111",14793 => "10100100",14794 => "00100010",14795 => "01111010",14796 => "11111011",14797 => "00111101",14798 => "10110110",14799 => "10111100",14800 => "01101100",14801 => "11010011",14802 => "11001010",14803 => "00111110",14804 => "00101100",14805 => "10111100",14806 => "11011101",14807 => "10100000",14808 => "00100001",14809 => "01001000",14810 => "00110000",14811 => "10011100",14812 => "01101010",14813 => "00111111",14814 => "10011101",14815 => "10010001",14816 => "00010000",14817 => "11000100",14818 => "11010000",14819 => "11111011",14820 => "00011010",14821 => "00111011",14822 => "10000010",14823 => "11001110",14824 => "00101001",14825 => "11000010",14826 => "00001000",14827 => "01110100",14828 => "11010110",14829 => "10000110",14830 => "00111111",14831 => "00010010",14832 => "11001110",14833 => "01001100",14834 => "00001101",14835 => "00110110",14836 => "01111100",14837 => "00001111",14838 => "11001001",14839 => "11111110",14840 => "11100001",14841 => "10110001",14842 => "00010101",14843 => "00110000",14844 => "10000110",14845 => "01011011",14846 => "10011001",14847 => "10111001",14848 => "10101110",14849 => "11000000",14850 => "01000001",14851 => "00111000",14852 => "00000100",14853 => "00101001",14854 => "01010001",14855 => "00011111",14856 => "01111011",14857 => "00010110",14858 => "00001101",14859 => "10001010",14860 => "00001000",14861 => "00001111",14862 => "01000010",14863 => "00010011",14864 => "10001001",14865 => "10001011",14866 => "00101111",14867 => "00110110",14868 => "10000111",14869 => "00000111",14870 => "01101100",14871 => "10110100",14872 => "11011111",14873 => "00010010",14874 => "01101000",14875 => "00101110",14876 => "10011001",14877 => "01010010",14878 => "00011011",14879 => "00001100",14880 => "10100100",14881 => "10000110",14882 => "00110110",14883 => "11011011",14884 => "00010100",14885 => "01100100",14886 => "10111000",14887 => "01011100",14888 => "11001101",14889 => "01000011",14890 => "00011001",14891 => "10011111",14892 => "10001100",14893 => "11110110",14894 => "01111101",14895 => "00001111",14896 => "01001111",14897 => "00110101",14898 => "10001010",14899 => "10100101",14900 => "00111100",14901 => "00000110",14902 => "01010011",14903 => "00011101",14904 => "10011110",14905 => "00010010",14906 => "00010110",14907 => "11111011",14908 => "11101000",14909 => "11010110",14910 => "10111111",14911 => "11011001",14912 => "11101000",14913 => "10001111",14914 => "10111011",14915 => "10111100",14916 => "00111110",14917 => "01100001",14918 => "10000111",14919 => "01110000",14920 => "01011100",14921 => "00100001",14922 => "10011010",14923 => "11010110",14924 => "11110111",14925 => "01110111",14926 => "00000011",14927 => "10101011",14928 => "11001101",14929 => "10011011",14930 => "00101011",14931 => "01111100",14932 => "10110001",14933 => "01010011",14934 => "10101101",14935 => "01110101",14936 => "10001000",14937 => "00101101",14938 => "00010011",14939 => "11010001",14940 => "01111010",14941 => "00111100",14942 => "11100101",14943 => "01110011",14944 => "10010101",14945 => "01100000",14946 => "00111001",14947 => "11010110",14948 => "00110110",14949 => "01011100",14950 => "10000001",14951 => "11100111",14952 => "00001011",14953 => "01111010",14954 => "11010100",14955 => "11001001",14956 => "01010111",14957 => "01010011",14958 => "00111000",14959 => "10101010",14960 => "01001111",14961 => "11001010",14962 => "01111101",14963 => "00100011",14964 => "11101010",14965 => "01011101",14966 => "01011101",14967 => "00100011",14968 => "11011111",14969 => "01001000",14970 => "00001111",14971 => "10000110",14972 => "11010110",14973 => "01001001",14974 => "11001010",14975 => "01000110",14976 => "01000000",14977 => "11100011",14978 => "10101000",14979 => "00001011",14980 => "00100010",14981 => "11110101",14982 => "10101011",14983 => "10111001",14984 => "01111000",14985 => "10111000",14986 => "01110100",14987 => "10100101",14988 => "00111010",14989 => "01111111",14990 => "11101101",14991 => "01001111",14992 => "01000011",14993 => "01000001",14994 => "01011100",14995 => "10100100",14996 => "11010011",14997 => "11000001",14998 => "00111000",14999 => "11010101",15000 => "01111000",15001 => "01101011",15002 => "01101001",15003 => "11011101",15004 => "01001111",15005 => "00010010",15006 => "00001111",15007 => "00000000",15008 => "00101111",15009 => "01100100",15010 => "10111110",15011 => "00110001",15012 => "11111111",15013 => "10000010",15014 => "01001100",15015 => "00001001",15016 => "10000000",15017 => "01001001",15018 => "10110010",15019 => "10111111",15020 => "10110111",15021 => "11010010",15022 => "01001011",15023 => "00110010",15024 => "10000101",15025 => "00100010",15026 => "10000011",15027 => "00101010",15028 => "11010111",15029 => "10111110",15030 => "10011010",15031 => "10110111",15032 => "11000001",15033 => "10111110",15034 => "11011001",15035 => "11000000",15036 => "00011100",15037 => "10001010",15038 => "10000000",15039 => "00001101",15040 => "01111100",15041 => "00101100",15042 => "11111010",15043 => "10100010",15044 => "01001010",15045 => "00010010",15046 => "11111110",15047 => "10001010",15048 => "11110010",15049 => "10001100",15050 => "11100000",15051 => "11000111",15052 => "00010011",15053 => "11111111",15054 => "11101110",15055 => "11011100",15056 => "01110101",15057 => "11111101",15058 => "10001000",15059 => "10010011",15060 => "10111010",15061 => "10010001",15062 => "10010001",15063 => "11010111",15064 => "11101100",15065 => "01011111",15066 => "01110100",15067 => "00100101",15068 => "01010101",15069 => "00100010",15070 => "10111100",15071 => "01001100",15072 => "01011110",15073 => "11010101",15074 => "10010101",15075 => "11110101",15076 => "01111100",15077 => "01100011",15078 => "10000001",15079 => "00011010",15080 => "00011000",15081 => "11011110",15082 => "00101010",15083 => "01110001",15084 => "11110111",15085 => "01100110",15086 => "11011001",15087 => "01110110",15088 => "10010001",15089 => "01001101",15090 => "11001110",15091 => "11110110",15092 => "00001000",15093 => "00111010",15094 => "00100010",15095 => "10010110",15096 => "01000011",15097 => "10011000",15098 => "01000010",15099 => "00110110",15100 => "11101101",15101 => "10010111",15102 => "01001011",15103 => "11100000",15104 => "01011001",15105 => "01001010",15106 => "10000000",15107 => "00001100",15108 => "10000111",15109 => "01101000",15110 => "11010000",15111 => "11001011",15112 => "11011011",15113 => "10101100",15114 => "00101100",15115 => "00110010",15116 => "00011100",15117 => "01000000",15118 => "11010100",15119 => "01001100",15120 => "01111101",15121 => "11101101",15122 => "00001110",15123 => "11001111",15124 => "10100100",15125 => "11111010",15126 => "10100110",15127 => "00100010",15128 => "00101000",15129 => "11101001",15130 => "10011111",15131 => "00110010",15132 => "10110111",15133 => "00110110",15134 => "10100011",15135 => "11001001",15136 => "10001101",15137 => "00000110",15138 => "10111011",15139 => "01001110",15140 => "10100110",15141 => "11011100",15142 => "01111101",15143 => "01010011",15144 => "00100011",15145 => "10011100",15146 => "00011011",15147 => "01000011",15148 => "01011111",15149 => "11001101",15150 => "11101000",15151 => "10101100",15152 => "01110110",15153 => "11000111",15154 => "10100000",15155 => "01110101",15156 => "00111110",15157 => "00010000",15158 => "11000001",15159 => "01101011",15160 => "11001101",15161 => "10000100",15162 => "10000010",15163 => "00001101",15164 => "00101011",15165 => "11100100",15166 => "00001100",15167 => "01110010",15168 => "01111100",15169 => "00001001",15170 => "11110101",15171 => "00011101",15172 => "01011111",15173 => "00101011",15174 => "10011111",15175 => "10001001",15176 => "00000000",15177 => "11000101",15178 => "01010000",15179 => "10011001",15180 => "00011011",15181 => "11100110",15182 => "00011011",15183 => "10110011",15184 => "11100101",15185 => "01110000",15186 => "11111101",15187 => "10101011",15188 => "10111000",15189 => "01010101",15190 => "10110100",15191 => "00011101",15192 => "11101110",15193 => "01010000",15194 => "01110101",15195 => "11001011",15196 => "10011010",15197 => "11011000",15198 => "10001110",15199 => "11101010",15200 => "00101010",15201 => "11110001",15202 => "10010010",15203 => "10011111",15204 => "00010000",15205 => "11010110",15206 => "11110000",15207 => "10011101",15208 => "10010111",15209 => "11101100",15210 => "10111000",15211 => "10011100",15212 => "10101111",15213 => "10000011",15214 => "11000010",15215 => "01011001",15216 => "10101110",15217 => "00110011",15218 => "11010011",15219 => "00110101",15220 => "00000001",15221 => "10010101",15222 => "00110001",15223 => "01011101",15224 => "11110010",15225 => "10111010",15226 => "01000001",15227 => "00111100",15228 => "11100101",15229 => "11010101",15230 => "10101010",15231 => "10000000",15232 => "11010000",15233 => "00011011",15234 => "11011011",15235 => "00111011",15236 => "11011001",15237 => "11010001",15238 => "01110001",15239 => "10010000",15240 => "10110000",15241 => "10010001",15242 => "11010111",15243 => "00101001",15244 => "00101001",15245 => "01011010",15246 => "00100011",15247 => "00000010",15248 => "01010001",15249 => "11011111",15250 => "11110101",15251 => "00101000",15252 => "11101001",15253 => "11010110",15254 => "01011101",15255 => "01000011",15256 => "10001001",15257 => "01011000",15258 => "11001000",15259 => "10100010",15260 => "11000101",15261 => "01011101",15262 => "10011011",15263 => "11110111",15264 => "01110110",15265 => "10001100",15266 => "11001001",15267 => "00110110",15268 => "01111000",15269 => "10011101",15270 => "01000110",15271 => "00010111",15272 => "10101111",15273 => "01101110",15274 => "01010111",15275 => "01000110",15276 => "01110110",15277 => "10111010",15278 => "11101001",15279 => "10011000",15280 => "00101010",15281 => "01100101",15282 => "11110110",15283 => "01001010",15284 => "10111010",15285 => "10000000",15286 => "00100101",15287 => "10000110",15288 => "01110010",15289 => "01001010",15290 => "01111011",15291 => "00010011",15292 => "11100100",15293 => "11000101",15294 => "11110101",15295 => "10000010",15296 => "01010111",15297 => "10100100",15298 => "10101101",15299 => "00110110",15300 => "10111000",15301 => "01111111",15302 => "00001101",15303 => "01000111",15304 => "01110011",15305 => "11000001",15306 => "11001011",15307 => "00100111",15308 => "00000010",15309 => "11101001",15310 => "10000111",15311 => "10111011",15312 => "10000001",15313 => "00110100",15314 => "00101101",15315 => "01111100",15316 => "10011110",15317 => "10001001",15318 => "11000100",15319 => "11100111",15320 => "11111111",15321 => "10111010",15322 => "01111111",15323 => "01111001",15324 => "10000000",15325 => "00010001",15326 => "10001001",15327 => "00011001",15328 => "00110010",15329 => "00100001",15330 => "10011010",15331 => "00000001",15332 => "10011110",15333 => "11100111",15334 => "00111000",15335 => "10111111",15336 => "11111110",15337 => "01110101",15338 => "10101100",15339 => "00100001",15340 => "10000000",15341 => "01010011",15342 => "00111101",15343 => "11001100",15344 => "11000100",15345 => "00010111",15346 => "11011011",15347 => "10000111",15348 => "10111100",15349 => "10010100",15350 => "01010101",15351 => "00110101",15352 => "11101001",15353 => "01000101",15354 => "01110100",15355 => "01000010",15356 => "10001001",15357 => "11010111",15358 => "01100100",15359 => "10101111",15360 => "00000101",15361 => "10100011",15362 => "01010000",15363 => "00110100",15364 => "00010111",15365 => "11011111",15366 => "10000001",15367 => "01101101",15368 => "00100011",15369 => "00000011",15370 => "11100111",15371 => "00000001",15372 => "01001001",15373 => "10101100",15374 => "00011011",15375 => "01010110",15376 => "10011110",15377 => "01111111",15378 => "00000110",15379 => "11010000",15380 => "01101000",15381 => "10010101",15382 => "11101000",15383 => "01100000",15384 => "00011011",15385 => "10111011",15386 => "00001101",15387 => "11001011",15388 => "01111110",15389 => "00011011",15390 => "10101101",15391 => "01011111",15392 => "10110100",15393 => "01010001",15394 => "10101110",15395 => "10000100",15396 => "00011001",15397 => "00001101",15398 => "00011110",15399 => "00011000",15400 => "01100110",15401 => "10000001",15402 => "01000010",15403 => "01000001",15404 => "00000010",15405 => "11110111",15406 => "10000001",15407 => "11101100",15408 => "10101100",15409 => "01100110",15410 => "10001010",15411 => "10000011",15412 => "11000010",15413 => "10001010",15414 => "11000001",15415 => "11010110",15416 => "00100100",15417 => "11011101",15418 => "01010111",15419 => "10100110",15420 => "10110001",15421 => "01010000",15422 => "11010011",15423 => "11101000",15424 => "01110100",15425 => "01001001",15426 => "01011001",15427 => "10110101",15428 => "10010111",15429 => "00011110",15430 => "10100100",15431 => "01110010",15432 => "01100011",15433 => "11001101",15434 => "01001100",15435 => "01001101",15436 => "00100000",15437 => "01110001",15438 => "10001010",15439 => "11001011",15440 => "00011011",15441 => "00011110",15442 => "00001000",15443 => "11100011",15444 => "01000010",15445 => "01010011",15446 => "11100001",15447 => "11001001",15448 => "10110100",15449 => "10101111",15450 => "11100011",15451 => "10000010",15452 => "11101001",15453 => "00001111",15454 => "10110011",15455 => "01001100",15456 => "10100100",15457 => "01001101",15458 => "10000100",15459 => "11011011",15460 => "10111000",15461 => "01101011",15462 => "00110110",15463 => "11100010",15464 => "11100111",15465 => "11110111",15466 => "11001010",15467 => "11011011",15468 => "11011001",15469 => "01111111",15470 => "10010011",15471 => "00100101",15472 => "01101010",15473 => "11100011",15474 => "01110111",15475 => "11001001",15476 => "11111110",15477 => "01000001",15478 => "01111011",15479 => "11011110",15480 => "11010100",15481 => "11001101",15482 => "11101111",15483 => "10110110",15484 => "11111001",15485 => "01100000",15486 => "11111000",15487 => "01111010",15488 => "00011011",15489 => "01010110",15490 => "11001111",15491 => "10110101",15492 => "10011100",15493 => "01111010",15494 => "01111010",15495 => "10110101",15496 => "11000111",15497 => "10000100",15498 => "00001101",15499 => "01010100",15500 => "11010010",15501 => "01011100",15502 => "10101110",15503 => "00101000",15504 => "01110000",15505 => "00011110",15506 => "00101001",15507 => "01011101",15508 => "00000011",15509 => "10010111",15510 => "00011010",15511 => "00111001",15512 => "01010100",15513 => "00111110",15514 => "01001010",15515 => "00111100",15516 => "11001001",15517 => "10110011",15518 => "01111101",15519 => "11110111",15520 => "10111001",15521 => "01000101",15522 => "01011010",15523 => "11101110",15524 => "01111100",15525 => "00001100",15526 => "10111010",15527 => "11101101",15528 => "11110101",15529 => "10011100",15530 => "00001111",15531 => "00100111",15532 => "11000111",15533 => "00100010",15534 => "10011111",15535 => "00011101",15536 => "11000110",15537 => "11111111",15538 => "01011001",15539 => "11000011",15540 => "10100100",15541 => "10100011",15542 => "00000100",15543 => "01010100",15544 => "11110001",15545 => "10110100",15546 => "00100100",15547 => "01001110",15548 => "11000110",15549 => "00100101",15550 => "01101011",15551 => "01000111",15552 => "10000110",15553 => "11010110",15554 => "10000110",15555 => "11110111",15556 => "10100000",15557 => "10000110",15558 => "10100001",15559 => "00110001",15560 => "01111101",15561 => "00000000",15562 => "11110001",15563 => "01110100",15564 => "11110000",15565 => "10100101",15566 => "00011100",15567 => "00110010",15568 => "11100110",15569 => "00111111",15570 => "11101101",15571 => "01110111",15572 => "11110001",15573 => "00100100",15574 => "00100111",15575 => "00101101",15576 => "10000110",15577 => "01100001",15578 => "00011011",15579 => "00011010",15580 => "11110110",15581 => "01000000",15582 => "00001010",15583 => "11001000",15584 => "01000100",15585 => "00000101",15586 => "00000010",15587 => "10001100",15588 => "01111100",15589 => "00011000",15590 => "10011000",15591 => "00000100",15592 => "11000100",15593 => "01110111",15594 => "00010000",15595 => "00011100",15596 => "11001110",15597 => "11000000",15598 => "00010101",15599 => "11111111",15600 => "10111110",15601 => "01100010",15602 => "10110100",15603 => "01101011",15604 => "00111001",15605 => "01011000",15606 => "11011100",15607 => "00111011",15608 => "10101101",15609 => "11111110",15610 => "01010000",15611 => "01100111",15612 => "10001100",15613 => "01101110",15614 => "01101011",15615 => "01101011",15616 => "01010100",15617 => "00000011",15618 => "11001100",15619 => "10000000",15620 => "11011011",15621 => "01010100",15622 => "10101001",15623 => "11000011",15624 => "00011001",15625 => "10111101",15626 => "10000000",15627 => "11001001",15628 => "10001010",15629 => "01100011",15630 => "01000111",15631 => "01001011",15632 => "00100100",15633 => "10101011",15634 => "10011010",15635 => "01110100",15636 => "11110010",15637 => "00101100",15638 => "00100010",15639 => "10100011",15640 => "00000111",15641 => "11010110",15642 => "01100111",15643 => "01001011",15644 => "11010000",15645 => "00100111",15646 => "10101001",15647 => "11111110",15648 => "11001001",15649 => "01000101",15650 => "11100011",15651 => "10011100",15652 => "01010011",15653 => "00000011",15654 => "00000011",15655 => "01111100",15656 => "01000000",15657 => "01010101",15658 => "01010011",15659 => "11001011",15660 => "10101010",15661 => "11100100",15662 => "11011010",15663 => "11111001",15664 => "10111111",15665 => "11011111",15666 => "11111010",15667 => "00111000",15668 => "00011000",15669 => "00100111",15670 => "01011100",15671 => "01011101",15672 => "00110100",15673 => "10011011",15674 => "00101001",15675 => "01100000",15676 => "00000000",15677 => "10100011",15678 => "00110111",15679 => "10000100",15680 => "10000001",15681 => "00000001",15682 => "10001101",15683 => "11111010",15684 => "10010100",15685 => "11001111",15686 => "11001000",15687 => "01111011",15688 => "00101010",15689 => "10000010",15690 => "10001001",15691 => "11000001",15692 => "00110100",15693 => "11111011",15694 => "00100001",15695 => "01001010",15696 => "00010110",15697 => "01100100",15698 => "00111000",15699 => "10000010",15700 => "01001001",15701 => "10101110",15702 => "01011010",15703 => "10110011",15704 => "01110100",15705 => "10110000",15706 => "11001101",15707 => "00001011",15708 => "11001000",15709 => "00001011",15710 => "10100000",15711 => "11100111",15712 => "11011100",15713 => "10010111",15714 => "11110001",15715 => "01010011",15716 => "01101101",15717 => "01110010",15718 => "10001000",15719 => "10111101",15720 => "10111000",15721 => "10010011",15722 => "00010101",15723 => "01111110",15724 => "00010011",15725 => "10111100",15726 => "11010111",15727 => "10011011",15728 => "11110100",15729 => "01111111",15730 => "10101001",15731 => "00001001",15732 => "01110110",15733 => "01011001",15734 => "10110111",15735 => "00111001",15736 => "00011011",15737 => "10111010",15738 => "00011111",15739 => "01001001",15740 => "10111110",15741 => "01110101",15742 => "10101100",15743 => "10010010",15744 => "11111101",15745 => "00111101",15746 => "10000111",15747 => "00101001",15748 => "00011101",15749 => "11010011",15750 => "01101001",15751 => "01010100",15752 => "11101000",15753 => "00000001",15754 => "01001011",15755 => "11100110",15756 => "01101000",15757 => "11010110",15758 => "10111110",15759 => "00011100",15760 => "00101100",15761 => "10110011",15762 => "10111011",15763 => "01000110",15764 => "10100001",15765 => "00000100",15766 => "10011011",15767 => "01100111",15768 => "11101111",15769 => "00010010",15770 => "01001101",15771 => "00001010",15772 => "00011100",15773 => "01010000",15774 => "01010010",15775 => "11001000",15776 => "01110010",15777 => "11001010",15778 => "00010001",15779 => "01110000",15780 => "01111101",15781 => "11001001",15782 => "10101101",15783 => "11000101",15784 => "10100100",15785 => "11101110",15786 => "00100111",15787 => "00110011",15788 => "00011000",15789 => "11111011",15790 => "00010110",15791 => "00011000",15792 => "10111111",15793 => "00011001",15794 => "11100000",15795 => "11000110",15796 => "01001100",15797 => "01001010",15798 => "11100101",15799 => "11101101",15800 => "10011011",15801 => "00110010",15802 => "00010010",15803 => "11110111",15804 => "01010100",15805 => "10110010",15806 => "00100110",15807 => "00011001",15808 => "10100011",15809 => "11000010",15810 => "01000100",15811 => "11000010",15812 => "10001011",15813 => "10111001",15814 => "01110001",15815 => "00000001",15816 => "11010000",15817 => "10110100",15818 => "10100000",15819 => "01100010",15820 => "10011101",15821 => "10010000",15822 => "01111110",15823 => "01000111",15824 => "01011001",15825 => "11100110",15826 => "00011000",15827 => "00111001",15828 => "01110011",15829 => "10010101",15830 => "00111010",15831 => "11111100",15832 => "11100100",15833 => "01101101",15834 => "10000110",15835 => "10010100",15836 => "00001101",15837 => "11001001",15838 => "01001001",15839 => "00111100",15840 => "11001010",15841 => "10010011",15842 => "00000110",15843 => "01010111",15844 => "11100000",15845 => "00110111",15846 => "01010111",15847 => "11001001",15848 => "11101110",15849 => "01111000",15850 => "10111000",15851 => "01011011",15852 => "11011000",15853 => "01111100",15854 => "10110011",15855 => "00000111",15856 => "00101111",15857 => "01110101",15858 => "10010001",15859 => "11010101",15860 => "11101111",15861 => "10010001",15862 => "10010000",15863 => "01011101",15864 => "01111101",15865 => "11010000",15866 => "00101110",15867 => "01001010",15868 => "10000111",15869 => "11010100",15870 => "00110101",15871 => "01011011",15872 => "10100011",15873 => "00010010",15874 => "11010010",15875 => "00010011",15876 => "11010111",15877 => "11011010",15878 => "11001010",15879 => "11100100",15880 => "11100111",15881 => "10001100",15882 => "10110010",15883 => "00001001",15884 => "10000000",15885 => "10001011",15886 => "11110110",15887 => "11100111",15888 => "11011010",15889 => "10010010",15890 => "11110010",15891 => "10010000",15892 => "00111111",15893 => "01000010",15894 => "10100010",15895 => "11100101",15896 => "00000100",15897 => "01110000",15898 => "10000101",15899 => "00101110",15900 => "01001000",15901 => "11001011",15902 => "00000111",15903 => "00100101",15904 => "10100011",15905 => "00011011",15906 => "01101001",15907 => "00111000",15908 => "10000011",15909 => "10110010",15910 => "10101000",15911 => "10110100",15912 => "10110011",15913 => "10000010",15914 => "01010101",15915 => "00011001",15916 => "11101001",15917 => "00101100",15918 => "01101100",15919 => "01111110",15920 => "10111101",15921 => "00011001",15922 => "11100001",15923 => "11011000",15924 => "00011111",15925 => "10110100",15926 => "10001010",15927 => "11011100",15928 => "00010110",15929 => "10111111",15930 => "11001001",15931 => "01100110",15932 => "11000100",15933 => "11000010",15934 => "00111101",15935 => "10010110",15936 => "00100011",15937 => "10011101",15938 => "10010110",15939 => "11010011",15940 => "00110101",15941 => "10011111",15942 => "01111010",15943 => "10001100",15944 => "00110010",15945 => "11111001",15946 => "00111010",15947 => "10000001",15948 => "00000001",15949 => "00111111",15950 => "01110111",15951 => "10011110",15952 => "11111010",15953 => "10000101",15954 => "01010110",15955 => "00110100",15956 => "10111111",15957 => "11011010",15958 => "01000111",15959 => "10000000",15960 => "10011011",15961 => "11101011",15962 => "01001110",15963 => "01100110",15964 => "10111100",15965 => "11111111",15966 => "11010000",15967 => "11100011",15968 => "11100010",15969 => "00100001",15970 => "10000001",15971 => "11000100",15972 => "10100001",15973 => "10001110",15974 => "11000001",15975 => "00111010",15976 => "01000011",15977 => "11001110",15978 => "11101101",15979 => "10101000",15980 => "10111110",15981 => "00001101",15982 => "00010100",15983 => "10011110",15984 => "11000111",15985 => "10011000",15986 => "11001000",15987 => "11110100",15988 => "01101000",15989 => "01010110",15990 => "11011100",15991 => "10000101",15992 => "01000111",15993 => "10111101",15994 => "11101111",15995 => "01111001",15996 => "11101010",15997 => "11101101",15998 => "01000100",15999 => "01111011",16000 => "00101001",16001 => "11011000",16002 => "00100001",16003 => "10000111",16004 => "00110101",16005 => "00001010",16006 => "01000101",16007 => "10011011",16008 => "00100011",16009 => "01111000",16010 => "11001101",16011 => "01101101",16012 => "10111000",16013 => "00001010",16014 => "10110001",16015 => "00000100",16016 => "00010011",16017 => "01100111",16018 => "00110101",16019 => "00001100",16020 => "01111010",16021 => "10011101",16022 => "10101110",16023 => "01000001",16024 => "00110101",16025 => "11001000",16026 => "10110100",16027 => "10000110",16028 => "10000010",16029 => "10000111",16030 => "00000011",16031 => "01110100",16032 => "01100110",16033 => "00101000",16034 => "00101110",16035 => "01000111",16036 => "00100010",16037 => "11101111",16038 => "11011110",16039 => "10000000",16040 => "11011011",16041 => "11000100",16042 => "01010011",16043 => "01010100",16044 => "10001100",16045 => "01110101",16046 => "01110100",16047 => "11100000",16048 => "11011111",16049 => "11011010",16050 => "11101000",16051 => "01001001",16052 => "00001010",16053 => "00001000",16054 => "10100111",16055 => "01100000",16056 => "10011110",16057 => "11010011",16058 => "10011001",16059 => "10111011",16060 => "11010001",16061 => "10111001",16062 => "10000111",16063 => "10110000",16064 => "11110011",16065 => "11100000",16066 => "11010110",16067 => "01001000",16068 => "11010110",16069 => "11010011",16070 => "00110001",16071 => "10011111",16072 => "10011000",16073 => "00011110",16074 => "01011010",16075 => "11010100",16076 => "00101000",16077 => "11000101",16078 => "01010101",16079 => "11100011",16080 => "00001011",16081 => "01000100",16082 => "01011001",16083 => "11110010",16084 => "10001001",16085 => "00001110",16086 => "00100110",16087 => "11111101",16088 => "10000111",16089 => "00100101",16090 => "10011010",16091 => "10110110",16092 => "01100000",16093 => "10110001",16094 => "00011111",16095 => "00110100",16096 => "01011111",16097 => "10110011",16098 => "11100110",16099 => "01101100",16100 => "10111001",16101 => "11111001",16102 => "01100110",16103 => "10001101",16104 => "01011101",16105 => "01000000",16106 => "11000000",16107 => "11010011",16108 => "10001111",16109 => "11011110",16110 => "11100010",16111 => "10111101",16112 => "11001100",16113 => "01111000",16114 => "11111010",16115 => "00101101",16116 => "01010101",16117 => "01000110",16118 => "11010011",16119 => "10101011",16120 => "01010110",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00111110" report "FAIL high bits" severity failure;
assert RAM(0) = "11111000" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
