 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "11101000",3 => "01111011",4 => "00001100",5 => "01001111",6 => "10100110",7 => "10110011",8 => "01000111",9 => "00000111",10 => "00111011",11 => "10001100",12 => "00000101",13 => "00111100",14 => "10001101",15 => "00111010",16 => "10100110",17 => "00011101",18 => "00110001",19 => "01010110",20 => "10011000",21 => "00000101",22 => "00111010",23 => "00100011",24 => "11000001",25 => "01010011",26 => "00110100",27 => "11001111",28 => "00001111",29 => "11010000",30 => "11110011",31 => "01000000",32 => "01000011",33 => "01011000",34 => "10011101",35 => "01001100",36 => "01010010",37 => "11111111",38 => "11101010",39 => "01111010",40 => "01010111",41 => "01011001",42 => "01000010",43 => "00110011",44 => "01010101",45 => "11100101",46 => "00001011",47 => "11111111",48 => "00111001",49 => "00111111",50 => "01100111",51 => "00011101",52 => "11000001",53 => "01110001",54 => "01001101",55 => "11011100",56 => "00111100",57 => "00010000",58 => "00101101",59 => "01100010",60 => "01001111",61 => "10010110",62 => "10000011",63 => "10010001",64 => "11111001",65 => "01100101",66 => "01101001",67 => "11010100",68 => "00111100",69 => "10011111",70 => "01010011",71 => "11101000",72 => "10111000",73 => "11111000",74 => "00101010",75 => "11100100",76 => "11011001",77 => "01001100",78 => "01111001",79 => "01010010",80 => "00111110",81 => "00100101",82 => "00001110",83 => "00000011",84 => "00000010",85 => "00001011",86 => "10001001",87 => "00010111",88 => "00010111",89 => "11100010",90 => "10010100",91 => "01101111",92 => "10101111",93 => "01100010",94 => "00101010",95 => "10101100",96 => "01010000",97 => "00010110",98 => "00110010",99 => "11011101",100 => "00111110",101 => "11100000",102 => "10100011",103 => "11110011",104 => "00101100",105 => "11101111",106 => "01000000",107 => "10011100",108 => "01010001",109 => "01000010",110 => "10000001",111 => "10000101",112 => "10111010",113 => "00001101",114 => "00100101",115 => "10011011",116 => "10010001",117 => "10011011",118 => "11010011",119 => "00010000",120 => "11110101",121 => "01110001",122 => "00111110",123 => "10111100",124 => "00001111",125 => "11100011",126 => "11111101",127 => "01111101",128 => "00011010",129 => "00101011",130 => "01101001",131 => "00110110",132 => "01001110",133 => "10010001",134 => "00001101",135 => "01110011",136 => "10001000",137 => "10011001",138 => "10000111",139 => "01011011",140 => "11110101",141 => "10011001",142 => "00010010",143 => "00001110",144 => "10001110",145 => "11110010",146 => "01011100",147 => "00110110",148 => "01111110",149 => "01111010",150 => "00111110",151 => "00011001",152 => "10001100",153 => "11010001",154 => "11100001",155 => "00011000",156 => "10000010",157 => "01111101",158 => "01000000",159 => "11000011",160 => "00001001",161 => "01110011",162 => "01111010",163 => "00100011",164 => "11011000",165 => "11110001",166 => "10011001",167 => "11110101",168 => "00000110",169 => "10010011",170 => "11001111",171 => "11010011",172 => "10101110",173 => "01010101",174 => "00011101",175 => "11100011",176 => "00110100",177 => "10000100",178 => "10111110",179 => "01100100",180 => "10100000",181 => "00101101",182 => "01100110",183 => "01100001",184 => "10011010",185 => "01110011",186 => "11110000",187 => "11100000",188 => "01011101",189 => "01101010",190 => "11000010",191 => "10111001",192 => "10110010",193 => "11110101",194 => "11101100",195 => "11010111",196 => "01000001",197 => "10111011",198 => "11010000",199 => "10101100",200 => "11111111",201 => "01111011",202 => "00110100",203 => "01100110",204 => "00010000",205 => "01010001",206 => "01101101",207 => "01100001",208 => "01001011",209 => "11101111",210 => "11111101",211 => "01011000",212 => "01101110",213 => "11000100",214 => "00001010",215 => "11101100",216 => "01010111",217 => "01111110",218 => "11010111",219 => "00111001",220 => "01111000",221 => "10100001",222 => "01011001",223 => "11000111",224 => "01010011",225 => "10000001",226 => "01110000",227 => "01000000",228 => "10001110",229 => "11111110",230 => "00100101",231 => "01001000",232 => "00101001",233 => "10111001",234 => "01000100",235 => "11001010",236 => "11100000",237 => "00001011",238 => "00001011",239 => "00110000",240 => "00000111",241 => "01010010",242 => "00010111",243 => "00111100",244 => "11011100",245 => "01001010",246 => "00000010",247 => "11100100",248 => "00101011",249 => "10010100",250 => "11000101",251 => "11110000",252 => "01101101",253 => "11100101",254 => "11101111",255 => "01101011",256 => "01010101",257 => "11100101",258 => "10011000",259 => "10011111",260 => "00110110",261 => "11010011",262 => "11110011",263 => "10001100",264 => "00000001",265 => "00110111",266 => "10000000",267 => "11011011",268 => "01110111",269 => "01101111",270 => "01100001",271 => "00000001",272 => "00010010",273 => "01001110",274 => "10000011",275 => "01111010",276 => "00100011",277 => "00110001",278 => "11011111",279 => "11010001",280 => "11101101",281 => "00111010",282 => "00101010",283 => "00110011",284 => "01011000",285 => "10001001",286 => "01000100",287 => "10001001",288 => "01101001",289 => "10110100",290 => "01001100",291 => "11010011",292 => "00001001",293 => "00011110",294 => "01110101",295 => "01010110",296 => "11010111",297 => "10000100",298 => "00110000",299 => "11100110",300 => "00011010",301 => "01100010",302 => "11100001",303 => "01101011",304 => "10010000",305 => "00100011",306 => "10110000",307 => "01011110",308 => "10010010",309 => "01000110",310 => "00001001",311 => "11110111",312 => "00000010",313 => "01001111",314 => "10100110",315 => "01110001",316 => "11001100",317 => "01101000",318 => "11001011",319 => "00001110",320 => "01110010",321 => "01101011",322 => "10101101",323 => "10011101",324 => "10001001",325 => "00111000",326 => "10011101",327 => "10101010",328 => "01000101",329 => "01110000",330 => "10111010",331 => "01000101",332 => "00111001",333 => "10001101",334 => "00011011",335 => "00101100",336 => "01011100",337 => "00011100",338 => "10000100",339 => "11011101",340 => "11111100",341 => "11111111",342 => "00110000",343 => "11011110",344 => "10000101",345 => "00001101",346 => "11111101",347 => "10011011",348 => "10111101",349 => "11101011",350 => "01001001",351 => "01100000",352 => "00101011",353 => "01010000",354 => "01000010",355 => "00000001",356 => "01000010",357 => "10000001",358 => "00110101",359 => "01101110",360 => "00110111",361 => "11110011",362 => "00010111",363 => "00000010",364 => "10010110",365 => "11001110",366 => "00011110",367 => "00101101",368 => "10110101",369 => "11011110",370 => "10111001",371 => "00101001",372 => "00011111",373 => "10100000",374 => "01100110",375 => "01000000",376 => "00100011",377 => "00001100",378 => "11011011",379 => "10010010",380 => "01101011",381 => "00001000",382 => "00110010",383 => "01000000",384 => "01001011",385 => "01000100",386 => "01001101",387 => "00111101",388 => "10000001",389 => "01000101",390 => "10010111",391 => "10001101",392 => "11111011",393 => "11010000",394 => "01010010",395 => "11011001",396 => "00101011",397 => "11010110",398 => "00111011",399 => "11111101",400 => "01000100",401 => "01011001",402 => "11000101",403 => "11010010",404 => "00010000",405 => "11001011",406 => "11000111",407 => "11010010",408 => "10111000",409 => "01110100",410 => "10011100",411 => "01111110",412 => "10111010",413 => "00101011",414 => "01111000",415 => "01011000",416 => "01000011",417 => "11100010",418 => "10100010",419 => "00101001",420 => "11111110",421 => "10100101",422 => "10111111",423 => "00000111",424 => "10110001",425 => "10000010",426 => "01100111",427 => "10100110",428 => "00110100",429 => "01011101",430 => "00110010",431 => "11101001",432 => "10101111",433 => "10000001",434 => "10001001",435 => "11110110",436 => "11000101",437 => "01110000",438 => "10111101",439 => "01110101",440 => "00110111",441 => "11111110",442 => "01110000",443 => "10001001",444 => "11011010",445 => "00101100",446 => "11101101",447 => "10010000",448 => "11110110",449 => "01010011",450 => "11011001",451 => "11010100",452 => "10110110",453 => "01110001",454 => "01001001",455 => "00111010",456 => "01101100",457 => "11111000",458 => "10000001",459 => "10111010",460 => "11010100",461 => "00110000",462 => "01101001",463 => "00010101",464 => "01011001",465 => "01001010",466 => "00010010",467 => "01101000",468 => "01000100",469 => "11110111",470 => "10010110",471 => "11001011",472 => "00010000",473 => "01010000",474 => "10110110",475 => "11011010",476 => "10000010",477 => "01100001",478 => "11100110",479 => "01110000",480 => "10010010",481 => "01101000",482 => "00111010",483 => "00000111",484 => "01001101",485 => "11010111",486 => "11111011",487 => "01010111",488 => "11010110",489 => "10111000",490 => "10011001",491 => "11011010",492 => "10000101",493 => "11011010",494 => "10010100",495 => "00100111",496 => "01011101",497 => "10010100",498 => "10010110",499 => "01011110",500 => "00011110",501 => "11011101",502 => "10011111",503 => "01010101",504 => "11111011",505 => "01001111",506 => "00101110",507 => "11101110",508 => "10001001",509 => "01110100",510 => "11011110",511 => "00101111",512 => "00000000",513 => "10001101",514 => "10011000",515 => "01110011",516 => "00101000",517 => "10000101",518 => "01110111",519 => "00101000",520 => "11100011",521 => "11001011",522 => "10001100",523 => "00100011",524 => "01111110",525 => "01000001",526 => "01110111",527 => "11101000",528 => "10111010",529 => "11101011",530 => "00001011",531 => "01111000",532 => "01111000",533 => "01010100",534 => "01111001",535 => "10111110",536 => "11001001",537 => "11000001",538 => "00010001",539 => "11000101",540 => "10000101",541 => "00000100",542 => "01110000",543 => "10010100",544 => "00101001",545 => "10010001",546 => "10110000",547 => "00110010",548 => "11000110",549 => "00111000",550 => "11101100",551 => "10001100",552 => "01010101",553 => "10000000",554 => "00111101",555 => "01110111",556 => "01011000",557 => "11101001",558 => "00010111",559 => "01101111",560 => "10010101",561 => "10110111",562 => "10100101",563 => "01010101",564 => "00000001",565 => "11101010",566 => "00000011",567 => "11000101",568 => "11011101",569 => "00100111",570 => "01100011",571 => "00101011",572 => "11111011",573 => "01000010",574 => "11010011",575 => "01010111",576 => "10100110",577 => "01110011",578 => "00001011",579 => "00000100",580 => "10100011",581 => "01001001",582 => "01000100",583 => "01110000",584 => "00100101",585 => "01101100",586 => "11100110",587 => "01001111",588 => "01001101",589 => "00111110",590 => "00110101",591 => "11111001",592 => "10011111",593 => "00000001",594 => "00001101",595 => "11101000",596 => "10011001",597 => "00100110",598 => "10110011",599 => "11101111",600 => "10100001",601 => "11010000",602 => "10011001",603 => "10011100",604 => "01100111",605 => "00110110",606 => "10000111",607 => "00011010",608 => "00000010",609 => "10011100",610 => "11101100",611 => "10100011",612 => "11011111",613 => "00001111",614 => "10010000",615 => "10100000",616 => "01110110",617 => "00110010",618 => "11001010",619 => "00111101",620 => "11001111",621 => "00110110",622 => "00010111",623 => "00001010",624 => "10101011",625 => "01110010",626 => "01001010",627 => "10111110",628 => "11111001",629 => "01100100",630 => "00001011",631 => "10011110",632 => "01000110",633 => "01001000",634 => "11010100",635 => "00001100",636 => "01000100",637 => "10010011",638 => "11010111",639 => "01011000",640 => "01010100",641 => "00100001",642 => "10010100",643 => "00111000",644 => "01011011",645 => "10110110",646 => "10010101",647 => "01011110",648 => "00001011",649 => "10001000",650 => "10111001",651 => "00001001",652 => "10110010",653 => "11001100",654 => "11100001",655 => "11000101",656 => "01011101",657 => "10100111",658 => "10101100",659 => "00000011",660 => "00000110",661 => "00111110",662 => "01010010",663 => "01011000",664 => "10100011",665 => "10110010",666 => "10110000",667 => "10100001",668 => "00011001",669 => "01111101",670 => "10101010",671 => "01100110",672 => "00000101",673 => "10000111",674 => "00100001",675 => "11010111",676 => "11000110",677 => "11101000",678 => "00011011",679 => "11010111",680 => "01100111",681 => "11000011",682 => "10101110",683 => "01101000",684 => "11001010",685 => "00001111",686 => "10110101",687 => "01000111",688 => "00100011",689 => "11010001",690 => "00011111",691 => "00101011",692 => "01101111",693 => "01110111",694 => "01010100",695 => "01110001",696 => "11110110",697 => "01101001",698 => "00011011",699 => "11011001",700 => "01100101",701 => "10010100",702 => "00110010",703 => "10111000",704 => "11110000",705 => "10010001",706 => "00001110",707 => "10100101",708 => "01110111",709 => "00010000",710 => "01111100",711 => "00101111",712 => "00010000",713 => "10001110",714 => "01100000",715 => "10010110",716 => "10010010",717 => "01010011",718 => "01100101",719 => "00011100",720 => "10001100",721 => "11110110",722 => "00000000",723 => "10011110",724 => "01111010",725 => "01011100",726 => "11010110",727 => "01111010",728 => "10001111",729 => "11101001",730 => "01100100",731 => "10110010",732 => "10100101",733 => "11100110",734 => "01101110",735 => "01100000",736 => "10101101",737 => "00100000",738 => "00111011",739 => "11111011",740 => "00010010",741 => "11001011",742 => "01011011",743 => "01001011",744 => "01000110",745 => "10010000",746 => "01001010",747 => "01000001",748 => "11001001",749 => "01100111",750 => "10011010",751 => "10001110",752 => "11000100",753 => "11001011",754 => "01110101",755 => "10110000",756 => "10111110",757 => "00010111",758 => "10100010",759 => "10010001",760 => "01100100",761 => "00111111",762 => "00100100",763 => "00001000",764 => "01010110",765 => "01011100",766 => "00101000",767 => "10111010",768 => "00001001",769 => "10001000",770 => "01111000",771 => "11101011",772 => "00110000",773 => "00100000",774 => "01000000",775 => "00101000",776 => "11011010",777 => "10011010",778 => "01000000",779 => "00100101",780 => "11110011",781 => "10110101",782 => "00011001",783 => "01100000",784 => "11110111",785 => "10101111",786 => "01000101",787 => "01001100",788 => "11100000",789 => "10110101",790 => "00011110",791 => "01001011",792 => "11011010",793 => "11100010",794 => "00011001",795 => "00101110",796 => "00001011",797 => "10101100",798 => "10101110",799 => "01101100",800 => "10110011",801 => "00011010",802 => "00011111",803 => "01101110",804 => "01000010",805 => "01100010",806 => "10110111",807 => "01111101",808 => "11011011",809 => "10011010",810 => "11110111",811 => "00001100",812 => "10000000",813 => "01010010",814 => "10110110",815 => "01101111",816 => "01101100",817 => "00001101",818 => "01101100",819 => "11100100",820 => "11000100",821 => "11000110",822 => "10010001",823 => "11101011",824 => "00000110",825 => "10001101",826 => "11011100",827 => "11001110",828 => "00100101",829 => "01111011",830 => "10011111",831 => "10100111",832 => "01111110",833 => "10011101",834 => "00001100",835 => "01101101",836 => "00011011",837 => "00010101",838 => "11001110",839 => "00000010",840 => "10000111",841 => "10010111",842 => "00011001",843 => "11010000",844 => "10000111",845 => "11010110",846 => "11111010",847 => "10010100",848 => "01110101",849 => "10001110",850 => "01111111",851 => "01000001",852 => "11101011",853 => "00010000",854 => "11010011",855 => "01111001",856 => "01001000",857 => "11101000",858 => "01001010",859 => "00101111",860 => "00001100",861 => "10000010",862 => "10001100",863 => "10101000",864 => "11100011",865 => "01010000",866 => "00110011",867 => "10111111",868 => "11010001",869 => "11000101",870 => "10100010",871 => "11100001",872 => "00001111",873 => "00011101",874 => "01111111",875 => "11100101",876 => "01010110",877 => "00110110",878 => "11110010",879 => "00101111",880 => "00011111",881 => "00011111",882 => "01011101",883 => "00010001",884 => "10011001",885 => "11001010",886 => "10000110",887 => "10110010",888 => "01101110",889 => "10000000",890 => "10000000",891 => "10110101",892 => "10011001",893 => "00100101",894 => "01001101",895 => "00000111",896 => "01001100",897 => "01111100",898 => "10111100",899 => "01111000",900 => "01101101",901 => "00001011",902 => "11011010",903 => "11101101",904 => "11100000",905 => "11111100",906 => "10111101",907 => "01001111",908 => "00110011",909 => "00100001",910 => "00001110",911 => "01111001",912 => "01100010",913 => "10011011",914 => "01101001",915 => "00101001",916 => "10111111",917 => "10101000",918 => "10000001",919 => "10101110",920 => "01100110",921 => "10100111",922 => "01101000",923 => "01111000",924 => "01100011",925 => "10001110",926 => "11111010",927 => "11101001",928 => "10011100",929 => "11000101",930 => "01111010",931 => "00010101",932 => "10010101",933 => "11110001",934 => "10000001",935 => "11011001",936 => "10100100",937 => "00010100",938 => "00101110",939 => "00111000",940 => "01111110",941 => "10010101",942 => "00111000",943 => "11111111",944 => "10100011",945 => "11000000",946 => "11000101",947 => "00111101",948 => "01001100",949 => "11011001",950 => "01110001",951 => "00000011",952 => "01101011",953 => "01001000",954 => "11111000",955 => "00100101",956 => "01110110",957 => "00111101",958 => "01001100",959 => "00000100",960 => "00001000",961 => "01011111",962 => "01111101",963 => "00101011",964 => "11000010",965 => "11000110",966 => "10101011",967 => "00001110",968 => "00011011",969 => "00010011",970 => "10110001",971 => "11110010",972 => "01000011",973 => "01111001",974 => "11001100",975 => "00100011",976 => "01010101",977 => "10000101",978 => "10000110",979 => "00111101",980 => "10100000",981 => "11101101",982 => "00100001",983 => "10100110",984 => "00011100",985 => "01011010",986 => "01101111",987 => "00110001",988 => "10001010",989 => "10100111",990 => "01011111",991 => "11011001",992 => "10100011",993 => "11100000",994 => "00000000",995 => "10001101",996 => "11011000",997 => "01101100",998 => "11111111",999 => "11000100",1000 => "11111100",1001 => "01110110",1002 => "11010011",1003 => "01110001",1004 => "00001001",1005 => "10001100",1006 => "10110010",1007 => "10101000",1008 => "10100010",1009 => "01111100",1010 => "10100101",1011 => "01110100",1012 => "11011110",1013 => "00101100",1014 => "00100100",1015 => "10110010",1016 => "10010101",1017 => "01111111",1018 => "11010000",1019 => "01011001",1020 => "01011010",1021 => "11011101",1022 => "11111000",1023 => "00001010",1024 => "10000000",1025 => "01000110",1026 => "00011010",1027 => "00101010",1028 => "10110010",1029 => "00000111",1030 => "11000100",1031 => "11001010",1032 => "10001110",1033 => "01000010",1034 => "11010101",1035 => "00110101",1036 => "01110111",1037 => "00110011",1038 => "11101110",1039 => "11011000",1040 => "11111000",1041 => "10001110",1042 => "10111101",1043 => "01011011",1044 => "10000000",1045 => "01100000",1046 => "00101110",1047 => "10011011",1048 => "10000010",1049 => "01110001",1050 => "00011011",1051 => "00011010",1052 => "00110100",1053 => "00011011",1054 => "11110000",1055 => "00001010",1056 => "10000110",1057 => "00000111",1058 => "00101110",1059 => "00101001",1060 => "11011110",1061 => "10111100",1062 => "01111001",1063 => "10011010",1064 => "10010101",1065 => "11010000",1066 => "01010001",1067 => "01000110",1068 => "10110001",1069 => "00110110",1070 => "10101011",1071 => "10110011",1072 => "01000101",1073 => "10111101",1074 => "00110000",1075 => "11100110",1076 => "11010100",1077 => "11011011",1078 => "01001011",1079 => "00000111",1080 => "11000001",1081 => "00110001",1082 => "11101111",1083 => "00111000",1084 => "10100011",1085 => "11001010",1086 => "00001101",1087 => "10010001",1088 => "11001111",1089 => "01101000",1090 => "10010100",1091 => "10111011",1092 => "10111110",1093 => "00011100",1094 => "10110111",1095 => "01011101",1096 => "01001101",1097 => "11001111",1098 => "01010001",1099 => "00000100",1100 => "01001000",1101 => "11111100",1102 => "11111110",1103 => "10101111",1104 => "00110110",1105 => "10111000",1106 => "01101111",1107 => "10010000",1108 => "11010110",1109 => "00110110",1110 => "01100111",1111 => "11101000",1112 => "01010110",1113 => "10100011",1114 => "11110111",1115 => "00111011",1116 => "10101111",1117 => "01000110",1118 => "10001000",1119 => "10101011",1120 => "10001001",1121 => "00100100",1122 => "10100110",1123 => "10101110",1124 => "01111101",1125 => "00010111",1126 => "01111110",1127 => "01011001",1128 => "00010010",1129 => "00011011",1130 => "00011010",1131 => "01101000",1132 => "11111011",1133 => "10101111",1134 => "11100010",1135 => "00101011",1136 => "00000110",1137 => "10011110",1138 => "11011000",1139 => "10011101",1140 => "11000010",1141 => "00010111",1142 => "11100100",1143 => "00100110",1144 => "10011010",1145 => "00011111",1146 => "11011000",1147 => "11001001",1148 => "01000001",1149 => "10011110",1150 => "11110011",1151 => "11001111",1152 => "00111111",1153 => "00111101",1154 => "01110110",1155 => "00011000",1156 => "11001011",1157 => "10111101",1158 => "11011001",1159 => "00001100",1160 => "11100100",1161 => "11000100",1162 => "10010001",1163 => "11000010",1164 => "11110111",1165 => "00110011",1166 => "00000000",1167 => "10011010",1168 => "11000000",1169 => "00011100",1170 => "00010000",1171 => "11011011",1172 => "01001101",1173 => "10111011",1174 => "00010111",1175 => "10010001",1176 => "00101111",1177 => "00111110",1178 => "11100110",1179 => "00101111",1180 => "00100010",1181 => "10010000",1182 => "11011100",1183 => "01110100",1184 => "10010111",1185 => "10011010",1186 => "01110101",1187 => "10011101",1188 => "01110111",1189 => "10000000",1190 => "00100110",1191 => "01001011",1192 => "01111100",1193 => "10111111",1194 => "11001010",1195 => "00110110",1196 => "10010011",1197 => "00010000",1198 => "01110101",1199 => "10111010",1200 => "01010110",1201 => "10000011",1202 => "00101100",1203 => "10001101",1204 => "01101100",1205 => "10010011",1206 => "00010101",1207 => "11101111",1208 => "10111110",1209 => "00011000",1210 => "01101001",1211 => "10010010",1212 => "10011100",1213 => "10101100",1214 => "11010111",1215 => "11100100",1216 => "10101101",1217 => "11110010",1218 => "01000111",1219 => "10111100",1220 => "10101001",1221 => "01011111",1222 => "00011010",1223 => "11110111",1224 => "10000010",1225 => "01100011",1226 => "11011110",1227 => "10000000",1228 => "11011100",1229 => "11111010",1230 => "11100110",1231 => "01110001",1232 => "01001111",1233 => "11100010",1234 => "00010111",1235 => "10001100",1236 => "11110101",1237 => "10001000",1238 => "01111010",1239 => "11110010",1240 => "01101110",1241 => "10101101",1242 => "10110010",1243 => "11100111",1244 => "10011100",1245 => "10011111",1246 => "00110010",1247 => "10010101",1248 => "10101011",1249 => "10100001",1250 => "00100111",1251 => "01101110",1252 => "00010101",1253 => "11011101",1254 => "11100110",1255 => "01111011",1256 => "01011100",1257 => "00011101",1258 => "10011111",1259 => "11001000",1260 => "01111110",1261 => "00111011",1262 => "00100000",1263 => "10101000",1264 => "10100001",1265 => "10101110",1266 => "01110101",1267 => "00100001",1268 => "11110001",1269 => "01011101",1270 => "01100111",1271 => "00001101",1272 => "00010011",1273 => "00010000",1274 => "10011011",1275 => "01101101",1276 => "00101001",1277 => "10110011",1278 => "11011010",1279 => "10100001",1280 => "00100010",1281 => "00100000",1282 => "00001111",1283 => "10100010",1284 => "00111000",1285 => "11001111",1286 => "00101001",1287 => "10010001",1288 => "01101110",1289 => "11010100",1290 => "11100101",1291 => "01101110",1292 => "10001110",1293 => "11101010",1294 => "01101001",1295 => "10110011",1296 => "10110000",1297 => "11011101",1298 => "01110100",1299 => "11101100",1300 => "00110110",1301 => "10110011",1302 => "10110010",1303 => "01111011",1304 => "00011100",1305 => "10111110",1306 => "01001011",1307 => "01101010",1308 => "10010110",1309 => "10101111",1310 => "00100111",1311 => "01110001",1312 => "00010010",1313 => "10010111",1314 => "11001011",1315 => "10011101",1316 => "00110011",1317 => "11110011",1318 => "11110100",1319 => "10101000",1320 => "11100111",1321 => "01001111",1322 => "01110101",1323 => "11001111",1324 => "00111000",1325 => "10001000",1326 => "01100110",1327 => "11000011",1328 => "10111100",1329 => "00111000",1330 => "01111100",1331 => "01100101",1332 => "11110011",1333 => "00010110",1334 => "01111101",1335 => "10111111",1336 => "01101001",1337 => "11010000",1338 => "11011000",1339 => "11001101",1340 => "01110011",1341 => "11001101",1342 => "11000111",1343 => "01001011",1344 => "11111110",1345 => "01001111",1346 => "01001010",1347 => "01110001",1348 => "11110001",1349 => "10001111",1350 => "00000011",1351 => "10010011",1352 => "01100001",1353 => "11101001",1354 => "11001100",1355 => "10100101",1356 => "00111110",1357 => "10000000",1358 => "01001010",1359 => "01110010",1360 => "11100001",1361 => "11100001",1362 => "01100001",1363 => "10101100",1364 => "00111000",1365 => "10110100",1366 => "11000110",1367 => "01011000",1368 => "11001100",1369 => "00010111",1370 => "00110100",1371 => "00101101",1372 => "11100111",1373 => "00000011",1374 => "11001111",1375 => "00011101",1376 => "10110101",1377 => "10111110",1378 => "10100100",1379 => "11110101",1380 => "00010101",1381 => "01110000",1382 => "11101001",1383 => "10011100",1384 => "00011111",1385 => "11111010",1386 => "00110101",1387 => "10001001",1388 => "01111011",1389 => "00011101",1390 => "00100001",1391 => "11001111",1392 => "11001000",1393 => "10111101",1394 => "10001111",1395 => "01100001",1396 => "11011110",1397 => "00101100",1398 => "00000111",1399 => "11111110",1400 => "11100111",1401 => "11110110",1402 => "11001110",1403 => "01111100",1404 => "11010001",1405 => "10000101",1406 => "10000010",1407 => "11001001",1408 => "01110101",1409 => "00001110",1410 => "11111000",1411 => "10100000",1412 => "00100101",1413 => "01101001",1414 => "00100000",1415 => "00111110",1416 => "00010100",1417 => "00100011",1418 => "11010011",1419 => "10001100",1420 => "01000010",1421 => "01001011",1422 => "00011010",1423 => "00010100",1424 => "10000010",1425 => "11110000",1426 => "11101110",1427 => "11000000",1428 => "11111011",1429 => "00010011",1430 => "11001110",1431 => "10010010",1432 => "00110100",1433 => "00001000",1434 => "01111001",1435 => "11000100",1436 => "00110101",1437 => "11001011",1438 => "01101011",1439 => "11000101",1440 => "00100000",1441 => "00110110",1442 => "11010101",1443 => "10011011",1444 => "10010101",1445 => "11011011",1446 => "01111001",1447 => "10101100",1448 => "00001111",1449 => "00001101",1450 => "11110111",1451 => "11110101",1452 => "11011111",1453 => "10111110",1454 => "10001010",1455 => "00110000",1456 => "00110111",1457 => "01111111",1458 => "00101111",1459 => "01001001",1460 => "11001101",1461 => "01111111",1462 => "11101101",1463 => "00111101",1464 => "00100110",1465 => "01001110",1466 => "10101010",1467 => "00011110",1468 => "01101000",1469 => "00110001",1470 => "10000110",1471 => "11000100",1472 => "11011101",1473 => "10000001",1474 => "01010000",1475 => "11110110",1476 => "10011111",1477 => "11111010",1478 => "11000000",1479 => "01011111",1480 => "10111010",1481 => "10000100",1482 => "10010110",1483 => "11000010",1484 => "10011010",1485 => "01010101",1486 => "00110110",1487 => "11111001",1488 => "01010101",1489 => "10011110",1490 => "10001101",1491 => "10001100",1492 => "01110010",1493 => "10001010",1494 => "10001110",1495 => "00110100",1496 => "01101011",1497 => "00010110",1498 => "01000101",1499 => "00001010",1500 => "00101010",1501 => "11011001",1502 => "01100100",1503 => "10110101",1504 => "00010000",1505 => "10111010",1506 => "00000100",1507 => "10100000",1508 => "10011011",1509 => "10001010",1510 => "11011100",1511 => "00011100",1512 => "00111011",1513 => "00011100",1514 => "11111000",1515 => "10011001",1516 => "11100101",1517 => "01011011",1518 => "10101110",1519 => "10011000",1520 => "11010111",1521 => "11000011",1522 => "10000110",1523 => "00110100",1524 => "10101110",1525 => "01101100",1526 => "01100101",1527 => "11000000",1528 => "11000000",1529 => "10101000",1530 => "10010110",1531 => "00011100",1532 => "01101010",1533 => "00000100",1534 => "10010111",1535 => "10110100",1536 => "00010000",1537 => "01111110",1538 => "01010111",1539 => "00110011",1540 => "01110111",1541 => "10111010",1542 => "11001101",1543 => "11010011",1544 => "01001001",1545 => "01001100",1546 => "01000100",1547 => "01010101",1548 => "10100101",1549 => "11111010",1550 => "00010000",1551 => "10001011",1552 => "01000110",1553 => "11010111",1554 => "00011001",1555 => "10100010",1556 => "00110000",1557 => "00100011",1558 => "01010110",1559 => "01010001",1560 => "10010001",1561 => "10110110",1562 => "11111100",1563 => "00111110",1564 => "00111110",1565 => "10101111",1566 => "11011011",1567 => "00110111",1568 => "00110110",1569 => "01000110",1570 => "00011010",1571 => "11010000",1572 => "11011111",1573 => "11000100",1574 => "11101010",1575 => "00101010",1576 => "11110001",1577 => "10010011",1578 => "11010001",1579 => "01001110",1580 => "00110101",1581 => "00100010",1582 => "11011101",1583 => "11110100",1584 => "11000100",1585 => "11111101",1586 => "11001001",1587 => "00000111",1588 => "01110011",1589 => "01000010",1590 => "10111011",1591 => "11011011",1592 => "01010101",1593 => "00111101",1594 => "11001000",1595 => "00011111",1596 => "01101001",1597 => "00111110",1598 => "01101110",1599 => "11110010",1600 => "10010011",1601 => "01100110",1602 => "11001011",1603 => "11100000",1604 => "11100011",1605 => "10000000",1606 => "00111111",1607 => "11101101",1608 => "01000000",1609 => "10001000",1610 => "11111101",1611 => "01001111",1612 => "00110010",1613 => "01111010",1614 => "01010110",1615 => "01011110",1616 => "10001100",1617 => "10010100",1618 => "10010111",1619 => "00111000",1620 => "00101100",1621 => "10101010",1622 => "01000001",1623 => "00111100",1624 => "01001011",1625 => "01001111",1626 => "10100110",1627 => "01001001",1628 => "10011100",1629 => "10100011",1630 => "01001011",1631 => "01111110",1632 => "01011011",1633 => "00010101",1634 => "11011001",1635 => "00110001",1636 => "00101010",1637 => "10000000",1638 => "11101000",1639 => "00111110",1640 => "01001101",1641 => "10010100",1642 => "00000111",1643 => "01001001",1644 => "01110101",1645 => "00101100",1646 => "11100100",1647 => "11111111",1648 => "01100100",1649 => "00110111",1650 => "01000111",1651 => "01011000",1652 => "00101011",1653 => "11101011",1654 => "10101101",1655 => "11000010",1656 => "00101000",1657 => "00101001",1658 => "11101010",1659 => "00100000",1660 => "10000000",1661 => "00010011",1662 => "10010001",1663 => "10001001",1664 => "11001101",1665 => "00001101",1666 => "01101100",1667 => "11000100",1668 => "01001001",1669 => "11100010",1670 => "00010100",1671 => "01011000",1672 => "01101011",1673 => "00000100",1674 => "11011010",1675 => "11111100",1676 => "01110101",1677 => "10101010",1678 => "01110100",1679 => "11110110",1680 => "11010101",1681 => "11011001",1682 => "01101010",1683 => "10011000",1684 => "10000000",1685 => "11001100",1686 => "00101000",1687 => "11011001",1688 => "01000100",1689 => "11000101",1690 => "01011110",1691 => "01111011",1692 => "11100011",1693 => "01110101",1694 => "11000100",1695 => "00101111",1696 => "01001101",1697 => "01110100",1698 => "00010100",1699 => "01011001",1700 => "00001100",1701 => "00101100",1702 => "00110011",1703 => "01001001",1704 => "11001000",1705 => "00000010",1706 => "10010101",1707 => "00101011",1708 => "01000011",1709 => "11111111",1710 => "01000001",1711 => "01001100",1712 => "01110010",1713 => "11001011",1714 => "10000000",1715 => "01011001",1716 => "11010011",1717 => "01000100",1718 => "10010111",1719 => "01000000",1720 => "11001001",1721 => "10000111",1722 => "10001001",1723 => "10011010",1724 => "11101001",1725 => "00110101",1726 => "10111110",1727 => "10000001",1728 => "00101001",1729 => "00011111",1730 => "00001001",1731 => "10001110",1732 => "00011001",1733 => "10101000",1734 => "10100011",1735 => "00001111",1736 => "01101110",1737 => "11000100",1738 => "01111001",1739 => "01010010",1740 => "00001110",1741 => "01001100",1742 => "11001011",1743 => "10101000",1744 => "11011111",1745 => "00101000",1746 => "11001010",1747 => "00010111",1748 => "10110110",1749 => "11010110",1750 => "11101000",1751 => "11011001",1752 => "00101111",1753 => "00100000",1754 => "01001011",1755 => "11110110",1756 => "10001111",1757 => "10001101",1758 => "11111101",1759 => "11011101",1760 => "00101000",1761 => "10100001",1762 => "00010110",1763 => "01011101",1764 => "00101011",1765 => "11111101",1766 => "01000010",1767 => "10110111",1768 => "10000101",1769 => "11101011",1770 => "10001010",1771 => "10101000",1772 => "10110110",1773 => "10111100",1774 => "00101111",1775 => "11000101",1776 => "11110011",1777 => "11011001",1778 => "11001111",1779 => "00101101",1780 => "10010110",1781 => "01000010",1782 => "11101010",1783 => "10111111",1784 => "01011011",1785 => "10101011",1786 => "11110011",1787 => "11001001",1788 => "01100101",1789 => "10101010",1790 => "11011010",1791 => "01001101",1792 => "00011100",1793 => "10111001",1794 => "00110101",1795 => "00001100",1796 => "11101101",1797 => "10110111",1798 => "00000100",1799 => "01010011",1800 => "01111110",1801 => "00111000",1802 => "00010101",1803 => "10010101",1804 => "00001000",1805 => "10111011",1806 => "00011110",1807 => "00001010",1808 => "11000100",1809 => "10100010",1810 => "10010001",1811 => "00010010",1812 => "10010100",1813 => "01111111",1814 => "01110011",1815 => "11010111",1816 => "10110011",1817 => "01110000",1818 => "11110001",1819 => "11110010",1820 => "01100110",1821 => "10100111",1822 => "00111011",1823 => "11111111",1824 => "11001011",1825 => "11101110",1826 => "10000000",1827 => "00000011",1828 => "01000000",1829 => "10111011",1830 => "10100011",1831 => "01001001",1832 => "11110101",1833 => "00001001",1834 => "11011010",1835 => "11010000",1836 => "10011011",1837 => "01000100",1838 => "01101100",1839 => "11100001",1840 => "01001011",1841 => "01010100",1842 => "11000101",1843 => "10110110",1844 => "10100001",1845 => "01001111",1846 => "00010001",1847 => "11110001",1848 => "00101011",1849 => "11110010",1850 => "00010001",1851 => "11110100",1852 => "11110000",1853 => "01100000",1854 => "11011010",1855 => "10100010",1856 => "01111000",1857 => "11010010",1858 => "00001000",1859 => "11001011",1860 => "00101110",1861 => "00001111",1862 => "11100011",1863 => "01000110",1864 => "01111000",1865 => "01011100",1866 => "10001010",1867 => "01101001",1868 => "10111001",1869 => "10101001",1870 => "00010001",1871 => "00101111",1872 => "11011110",1873 => "00000000",1874 => "00011100",1875 => "00010001",1876 => "10110001",1877 => "11110100",1878 => "00001110",1879 => "01010010",1880 => "10000011",1881 => "00101010",1882 => "10111000",1883 => "00001011",1884 => "10010111",1885 => "11011001",1886 => "01110010",1887 => "00111100",1888 => "00101101",1889 => "01000111",1890 => "00110100",1891 => "10110100",1892 => "10100110",1893 => "11100100",1894 => "01001011",1895 => "00110110",1896 => "01101111",1897 => "00100100",1898 => "01111101",1899 => "11001111",1900 => "01011111",1901 => "11110101",1902 => "00100100",1903 => "01001110",1904 => "10011010",1905 => "10101000",1906 => "11000111",1907 => "10100000",1908 => "01001010",1909 => "10010111",1910 => "10100100",1911 => "10010110",1912 => "00010000",1913 => "00111111",1914 => "10111001",1915 => "10011110",1916 => "11110010",1917 => "10010001",1918 => "11110111",1919 => "00000110",1920 => "11011110",1921 => "11001001",1922 => "10001101",1923 => "10110011",1924 => "00011100",1925 => "11111110",1926 => "00000010",1927 => "10000000",1928 => "10100011",1929 => "01000010",1930 => "00110001",1931 => "11000001",1932 => "11010010",1933 => "01010011",1934 => "11010111",1935 => "10000111",1936 => "11010010",1937 => "00001011",1938 => "00100100",1939 => "11000101",1940 => "10111100",1941 => "10111100",1942 => "01111001",1943 => "11111010",1944 => "11001100",1945 => "10000100",1946 => "01011110",1947 => "00010000",1948 => "00111101",1949 => "00111000",1950 => "01010001",1951 => "10011101",1952 => "01011000",1953 => "11101111",1954 => "11100110",1955 => "00110001",1956 => "00101100",1957 => "11100101",1958 => "11110110",1959 => "01000000",1960 => "00101100",1961 => "11100111",1962 => "01100010",1963 => "10111100",1964 => "11011110",1965 => "01010111",1966 => "00101000",1967 => "00000001",1968 => "10011100",1969 => "11001110",1970 => "10010001",1971 => "11010110",1972 => "10111101",1973 => "00001011",1974 => "10111100",1975 => "10001111",1976 => "11001110",1977 => "11101001",1978 => "10001100",1979 => "00101011",1980 => "11110101",1981 => "00001100",1982 => "10010001",1983 => "01100101",1984 => "10110110",1985 => "00000100",1986 => "11011010",1987 => "10000100",1988 => "00011011",1989 => "11011010",1990 => "11010011",1991 => "00100100",1992 => "11010111",1993 => "00111000",1994 => "10011011",1995 => "00100010",1996 => "00010010",1997 => "01010011",1998 => "10010001",1999 => "10000011",2000 => "01100011",2001 => "00001111",2002 => "00010011",2003 => "10010101",2004 => "11001100",2005 => "00100111",2006 => "01001111",2007 => "00011000",2008 => "01101001",2009 => "00010001",2010 => "10010101",2011 => "01010000",2012 => "11001111",2013 => "11111100",2014 => "11101010",2015 => "00111000",2016 => "00110101",2017 => "00000000",2018 => "11100001",2019 => "11101110",2020 => "01110110",2021 => "00011100",2022 => "00111010",2023 => "10000100",2024 => "00000011",2025 => "11111011",2026 => "11101010",2027 => "10111110",2028 => "00001111",2029 => "11110110",2030 => "11010010",2031 => "01111000",2032 => "10110101",2033 => "10110100",2034 => "11100101",2035 => "11110011",2036 => "01011000",2037 => "11111010",2038 => "01111100",2039 => "11110000",2040 => "11000001",2041 => "00100111",2042 => "00001010",2043 => "01100010",2044 => "10001101",2045 => "10011111",2046 => "10110010",2047 => "00111110",2048 => "10011011",2049 => "01011100",2050 => "10111011",2051 => "00000001",2052 => "11110111",2053 => "01010001",2054 => "11010000",2055 => "00000000",2056 => "11111100",2057 => "00011111",2058 => "10010100",2059 => "01000111",2060 => "10000011",2061 => "10000110",2062 => "11111011",2063 => "01001011",2064 => "01110110",2065 => "00100100",2066 => "01001100",2067 => "01111110",2068 => "11111100",2069 => "11011000",2070 => "10000010",2071 => "11011110",2072 => "00100111",2073 => "01010111",2074 => "11100110",2075 => "11001000",2076 => "11101001",2077 => "11001001",2078 => "10101110",2079 => "10000010",2080 => "00000011",2081 => "00110100",2082 => "01111011",2083 => "11110110",2084 => "10000101",2085 => "01100101",2086 => "11101100",2087 => "00001111",2088 => "11100000",2089 => "01100101",2090 => "10101101",2091 => "00101010",2092 => "00110001",2093 => "01111010",2094 => "11110001",2095 => "01010110",2096 => "10011010",2097 => "10100011",2098 => "11000010",2099 => "01101000",2100 => "00010011",2101 => "01010101",2102 => "00100000",2103 => "10110111",2104 => "11101111",2105 => "01100011",2106 => "10111000",2107 => "01101100",2108 => "01100010",2109 => "00110011",2110 => "11111100",2111 => "10011110",2112 => "00101011",2113 => "01111110",2114 => "10111111",2115 => "01011101",2116 => "10110001",2117 => "00011110",2118 => "10111110",2119 => "10010110",2120 => "11101011",2121 => "11010001",2122 => "00101011",2123 => "00010011",2124 => "01000101",2125 => "01010101",2126 => "11100111",2127 => "00011100",2128 => "01111110",2129 => "10111110",2130 => "11110011",2131 => "11111010",2132 => "00100010",2133 => "11101101",2134 => "00010011",2135 => "01000011",2136 => "00111001",2137 => "10011010",2138 => "01001011",2139 => "11010000",2140 => "10101001",2141 => "00111100",2142 => "01001010",2143 => "01001001",2144 => "01010111",2145 => "01110001",2146 => "00100001",2147 => "00010010",2148 => "01011111",2149 => "00101011",2150 => "01000001",2151 => "00010111",2152 => "10000100",2153 => "00010011",2154 => "11100011",2155 => "01001001",2156 => "01010001",2157 => "11101110",2158 => "11101011",2159 => "00000111",2160 => "01100101",2161 => "11001010",2162 => "10000010",2163 => "10110110",2164 => "00010011",2165 => "10011001",2166 => "10110101",2167 => "11101110",2168 => "00011110",2169 => "10110001",2170 => "00111000",2171 => "00101010",2172 => "01110010",2173 => "01110101",2174 => "10110010",2175 => "10010000",2176 => "10011001",2177 => "11001111",2178 => "01001011",2179 => "10101111",2180 => "00101001",2181 => "00110100",2182 => "01001010",2183 => "00011001",2184 => "11100000",2185 => "10011000",2186 => "11001101",2187 => "11111001",2188 => "10110011",2189 => "10010111",2190 => "10011010",2191 => "10111111",2192 => "10010101",2193 => "01100011",2194 => "10011010",2195 => "00010100",2196 => "00100110",2197 => "11000110",2198 => "00011000",2199 => "10101111",2200 => "10100101",2201 => "10011001",2202 => "11111001",2203 => "01010011",2204 => "01001110",2205 => "11101101",2206 => "00110010",2207 => "10000001",2208 => "01100001",2209 => "01101111",2210 => "11011000",2211 => "11100000",2212 => "00000000",2213 => "01011001",2214 => "00000000",2215 => "10110001",2216 => "10111100",2217 => "11000010",2218 => "10101010",2219 => "11011110",2220 => "10111101",2221 => "11111111",2222 => "01100110",2223 => "10101000",2224 => "11111110",2225 => "00110100",2226 => "11010100",2227 => "01011001",2228 => "10111100",2229 => "01100101",2230 => "10011111",2231 => "01110010",2232 => "00111100",2233 => "10000101",2234 => "01110011",2235 => "01101111",2236 => "01100001",2237 => "11001011",2238 => "11001110",2239 => "10000111",2240 => "10100001",2241 => "00111000",2242 => "11001001",2243 => "01100000",2244 => "10101000",2245 => "00001111",2246 => "11111011",2247 => "11100111",2248 => "10110010",2249 => "00010101",2250 => "01111100",2251 => "10011010",2252 => "11010011",2253 => "01011000",2254 => "00011111",2255 => "10101101",2256 => "01001010",2257 => "10110001",2258 => "10100101",2259 => "01010101",2260 => "01111100",2261 => "00110010",2262 => "01011001",2263 => "11111100",2264 => "10011010",2265 => "00010110",2266 => "10001100",2267 => "11111000",2268 => "10100010",2269 => "10000101",2270 => "00111111",2271 => "10111100",2272 => "01001010",2273 => "01110110",2274 => "10001101",2275 => "10010101",2276 => "11001011",2277 => "01100100",2278 => "11110001",2279 => "00000011",2280 => "10101000",2281 => "11010001",2282 => "11101001",2283 => "10111001",2284 => "10100101",2285 => "11011010",2286 => "11001111",2287 => "00110011",2288 => "11111110",2289 => "10011111",2290 => "11011110",2291 => "10101001",2292 => "01010011",2293 => "10010000",2294 => "10111110",2295 => "11110100",2296 => "10100111",2297 => "11001100",2298 => "00001010",2299 => "00110101",2300 => "00110000",2301 => "10100001",2302 => "11010111",2303 => "10011100",2304 => "10000010",2305 => "01000110",2306 => "01011111",2307 => "10111110",2308 => "11000011",2309 => "11000000",2310 => "00110111",2311 => "11001010",2312 => "11011101",2313 => "11010110",2314 => "00111101",2315 => "01010111",2316 => "10011101",2317 => "11101011",2318 => "10000011",2319 => "01010110",2320 => "00100000",2321 => "00111000",2322 => "11000111",2323 => "10111001",2324 => "01101000",2325 => "00000011",2326 => "11100101",2327 => "10111000",2328 => "11111010",2329 => "10000110",2330 => "10011110",2331 => "00010101",2332 => "11001110",2333 => "01000011",2334 => "01011110",2335 => "11011100",2336 => "00111010",2337 => "01010001",2338 => "01100110",2339 => "11010011",2340 => "00001110",2341 => "11101001",2342 => "11100100",2343 => "01010001",2344 => "00101110",2345 => "00001100",2346 => "10011011",2347 => "11110111",2348 => "10101111",2349 => "10000110",2350 => "01000001",2351 => "10111000",2352 => "11011011",2353 => "10101111",2354 => "00110100",2355 => "10000001",2356 => "11111010",2357 => "11000110",2358 => "11010111",2359 => "00100010",2360 => "10010001",2361 => "11100000",2362 => "00110011",2363 => "11101100",2364 => "00100111",2365 => "10000011",2366 => "11101101",2367 => "01110100",2368 => "01001110",2369 => "01011001",2370 => "01000100",2371 => "01000110",2372 => "11000010",2373 => "00000100",2374 => "00110101",2375 => "00001010",2376 => "00011110",2377 => "00110010",2378 => "11110011",2379 => "01000101",2380 => "00001110",2381 => "10111000",2382 => "10010011",2383 => "01011000",2384 => "00010000",2385 => "10011100",2386 => "11011110",2387 => "00111000",2388 => "10101101",2389 => "11100010",2390 => "00001011",2391 => "11110011",2392 => "10001100",2393 => "01110111",2394 => "11100101",2395 => "10111001",2396 => "00110100",2397 => "00001100",2398 => "00110000",2399 => "10001011",2400 => "10000100",2401 => "10011000",2402 => "10100001",2403 => "10010011",2404 => "01101000",2405 => "00111010",2406 => "11010000",2407 => "11011100",2408 => "11110011",2409 => "10111110",2410 => "10110100",2411 => "00110010",2412 => "01100000",2413 => "01110011",2414 => "11010001",2415 => "10011010",2416 => "10100001",2417 => "00000101",2418 => "01101000",2419 => "01011111",2420 => "10111011",2421 => "11111100",2422 => "01011011",2423 => "10100001",2424 => "00101110",2425 => "10111100",2426 => "11010001",2427 => "11000111",2428 => "11100000",2429 => "10110101",2430 => "00001011",2431 => "10100100",2432 => "10101010",2433 => "10000011",2434 => "01001000",2435 => "10000000",2436 => "01010100",2437 => "01010011",2438 => "00111110",2439 => "10101011",2440 => "01100101",2441 => "10001010",2442 => "11100111",2443 => "11001011",2444 => "11100111",2445 => "10010110",2446 => "10000010",2447 => "01101100",2448 => "11101101",2449 => "10110000",2450 => "01010100",2451 => "00101101",2452 => "01000000",2453 => "10001101",2454 => "00101011",2455 => "11101110",2456 => "00001000",2457 => "01111001",2458 => "10101100",2459 => "11010110",2460 => "11100010",2461 => "01111110",2462 => "00001000",2463 => "00110011",2464 => "11010011",2465 => "11001110",2466 => "11100001",2467 => "01011101",2468 => "10110011",2469 => "11010001",2470 => "11111111",2471 => "11111000",2472 => "10011101",2473 => "11110010",2474 => "10101101",2475 => "10100110",2476 => "01110100",2477 => "10010111",2478 => "01010111",2479 => "01010010",2480 => "11101011",2481 => "00000000",2482 => "00110111",2483 => "11100110",2484 => "00010011",2485 => "01011101",2486 => "00001011",2487 => "00011101",2488 => "01100100",2489 => "10011100",2490 => "01010001",2491 => "10011100",2492 => "00110000",2493 => "01111100",2494 => "00110101",2495 => "01111101",2496 => "10100011",2497 => "10110000",2498 => "01010101",2499 => "00011001",2500 => "11100011",2501 => "00110101",2502 => "11111011",2503 => "10010111",2504 => "00101011",2505 => "11110101",2506 => "11001010",2507 => "10111100",2508 => "01000100",2509 => "11000011",2510 => "10100111",2511 => "00100111",2512 => "01100000",2513 => "10000100",2514 => "00010001",2515 => "01001110",2516 => "11100100",2517 => "11100010",2518 => "01110111",2519 => "00111100",2520 => "10000111",2521 => "01100101",2522 => "10110111",2523 => "10110011",2524 => "00011010",2525 => "11110010",2526 => "01001101",2527 => "01100011",2528 => "00111000",2529 => "00000110",2530 => "01010111",2531 => "01101001",2532 => "11000011",2533 => "01110000",2534 => "01000001",2535 => "00101111",2536 => "11100001",2537 => "10001000",2538 => "10000110",2539 => "00110000",2540 => "11010110",2541 => "10001001",2542 => "11100100",2543 => "01111101",2544 => "11000001",2545 => "11101110",2546 => "00011011",2547 => "00010010",2548 => "01010000",2549 => "11011011",2550 => "01111000",2551 => "10101100",2552 => "00001101",2553 => "00110110",2554 => "10111000",2555 => "00001001",2556 => "11000011",2557 => "10110111",2558 => "01010001",2559 => "01101011",2560 => "10111000",2561 => "10001101",2562 => "11101110",2563 => "10011111",2564 => "11000011",2565 => "11011010",2566 => "10111010",2567 => "11011101",2568 => "10001010",2569 => "11010001",2570 => "01111111",2571 => "11100000",2572 => "01011111",2573 => "11111100",2574 => "00100110",2575 => "11011010",2576 => "10101110",2577 => "00111111",2578 => "10001001",2579 => "01000101",2580 => "01000000",2581 => "11010001",2582 => "01011011",2583 => "01011101",2584 => "01001000",2585 => "10101010",2586 => "01111001",2587 => "11100100",2588 => "00101101",2589 => "10110111",2590 => "11101011",2591 => "11001100",2592 => "01110100",2593 => "01111011",2594 => "01100011",2595 => "11100101",2596 => "01101010",2597 => "01111001",2598 => "10001110",2599 => "01110000",2600 => "00110000",2601 => "11110100",2602 => "11110110",2603 => "10011101",2604 => "00101101",2605 => "11110011",2606 => "11000101",2607 => "11100110",2608 => "10100010",2609 => "01110110",2610 => "10011110",2611 => "01011010",2612 => "11101001",2613 => "01101100",2614 => "00111000",2615 => "11001011",2616 => "01111100",2617 => "01111011",2618 => "11000001",2619 => "10001111",2620 => "10101010",2621 => "01010110",2622 => "10110000",2623 => "00100011",2624 => "01110111",2625 => "00001010",2626 => "10000111",2627 => "10110010",2628 => "00110100",2629 => "10110010",2630 => "00101111",2631 => "01110000",2632 => "01001100",2633 => "11101000",2634 => "01010110",2635 => "11010110",2636 => "11010111",2637 => "00111001",2638 => "11111010",2639 => "01101010",2640 => "01011101",2641 => "10111110",2642 => "10111010",2643 => "00111010",2644 => "00000000",2645 => "10110101",2646 => "01000010",2647 => "10101010",2648 => "00111000",2649 => "11101010",2650 => "11011011",2651 => "11001000",2652 => "01000100",2653 => "00000000",2654 => "10111100",2655 => "10110101",2656 => "11011001",2657 => "10000110",2658 => "01000010",2659 => "11010010",2660 => "00011011",2661 => "10001101",2662 => "01100110",2663 => "11001111",2664 => "11010111",2665 => "00010100",2666 => "10001001",2667 => "11100011",2668 => "01011110",2669 => "00111000",2670 => "01010110",2671 => "00010101",2672 => "01001110",2673 => "11110000",2674 => "00101000",2675 => "01101011",2676 => "00000111",2677 => "00100011",2678 => "00001000",2679 => "00000001",2680 => "10001010",2681 => "00010111",2682 => "01111100",2683 => "11100011",2684 => "10011111",2685 => "11110001",2686 => "01101001",2687 => "11100111",2688 => "11111101",2689 => "11111111",2690 => "00000000",2691 => "01000011",2692 => "00011011",2693 => "00100010",2694 => "10000010",2695 => "10101000",2696 => "11011101",2697 => "01001000",2698 => "00111101",2699 => "00101001",2700 => "11101100",2701 => "10100101",2702 => "10100110",2703 => "10111011",2704 => "01100000",2705 => "11010011",2706 => "10000010",2707 => "11100010",2708 => "00011110",2709 => "00101100",2710 => "00000111",2711 => "01000101",2712 => "01100101",2713 => "00110001",2714 => "11000110",2715 => "00000011",2716 => "10111110",2717 => "11000001",2718 => "11111111",2719 => "11101001",2720 => "11011001",2721 => "10101001",2722 => "00110111",2723 => "10110100",2724 => "00001101",2725 => "10110010",2726 => "01000001",2727 => "11011100",2728 => "10001010",2729 => "11101110",2730 => "01001110",2731 => "00101010",2732 => "10110001",2733 => "11110110",2734 => "11111010",2735 => "10010110",2736 => "10111111",2737 => "01011100",2738 => "11100110",2739 => "00000001",2740 => "11000011",2741 => "11001101",2742 => "00010100",2743 => "11011010",2744 => "00101100",2745 => "01010011",2746 => "11110111",2747 => "01110101",2748 => "11100110",2749 => "11011001",2750 => "01000100",2751 => "00000000",2752 => "00011011",2753 => "10111000",2754 => "11110111",2755 => "10111111",2756 => "00010000",2757 => "10011001",2758 => "11100110",2759 => "01110000",2760 => "01011011",2761 => "01010101",2762 => "00101100",2763 => "00110010",2764 => "01000011",2765 => "10111110",2766 => "10101011",2767 => "00011000",2768 => "01110000",2769 => "11101101",2770 => "10001110",2771 => "00110010",2772 => "01010100",2773 => "10011010",2774 => "00110011",2775 => "11011000",2776 => "00001010",2777 => "01100000",2778 => "11011101",2779 => "01110001",2780 => "00100000",2781 => "00000011",2782 => "10011001",2783 => "00101010",2784 => "10000100",2785 => "11011100",2786 => "00011010",2787 => "11011001",2788 => "01110100",2789 => "10001001",2790 => "01101100",2791 => "10000010",2792 => "10100000",2793 => "10111100",2794 => "10011110",2795 => "11000010",2796 => "00000001",2797 => "10001100",2798 => "01011100",2799 => "10101010",2800 => "11111100",2801 => "00011111",2802 => "00000100",2803 => "11110000",2804 => "00000001",2805 => "10100100",2806 => "11010000",2807 => "01110011",2808 => "01001110",2809 => "11100000",2810 => "00111010",2811 => "00100011",2812 => "11100001",2813 => "11001011",2814 => "01010001",2815 => "11001101",2816 => "01110110",2817 => "00001000",2818 => "00001100",2819 => "11011011",2820 => "00011000",2821 => "01011110",2822 => "00010011",2823 => "11101011",2824 => "11100101",2825 => "00100011",2826 => "00110100",2827 => "00010010",2828 => "10100010",2829 => "00000011",2830 => "00000110",2831 => "10011010",2832 => "11111110",2833 => "10000110",2834 => "01101111",2835 => "00011010",2836 => "01100100",2837 => "11110111",2838 => "10100101",2839 => "00000011",2840 => "11110100",2841 => "01011010",2842 => "01000101",2843 => "01011010",2844 => "11110010",2845 => "00010001",2846 => "01010101",2847 => "01001100",2848 => "10011000",2849 => "11110000",2850 => "01011111",2851 => "11000010",2852 => "01111111",2853 => "10011000",2854 => "01110010",2855 => "11001100",2856 => "00110101",2857 => "00110001",2858 => "11110001",2859 => "01000001",2860 => "00011010",2861 => "00101011",2862 => "10101011",2863 => "10110110",2864 => "00111010",2865 => "00000100",2866 => "01010110",2867 => "10100110",2868 => "10110000",2869 => "11001011",2870 => "00110001",2871 => "00100011",2872 => "00000001",2873 => "00001111",2874 => "11010000",2875 => "11111000",2876 => "00011010",2877 => "01001100",2878 => "01101100",2879 => "00011011",2880 => "01000000",2881 => "01110010",2882 => "00011100",2883 => "00110101",2884 => "11000110",2885 => "10010101",2886 => "01110101",2887 => "10101011",2888 => "11010111",2889 => "11111001",2890 => "11101111",2891 => "01011110",2892 => "10100000",2893 => "11110100",2894 => "11000000",2895 => "00110001",2896 => "11101010",2897 => "01011101",2898 => "01110101",2899 => "00000110",2900 => "01111000",2901 => "10011111",2902 => "10101111",2903 => "01101100",2904 => "01111011",2905 => "10111010",2906 => "11000000",2907 => "11000001",2908 => "01110001",2909 => "00100001",2910 => "00010010",2911 => "00111101",2912 => "01110011",2913 => "11000001",2914 => "00100000",2915 => "00111111",2916 => "11010110",2917 => "00001011",2918 => "11101010",2919 => "11010101",2920 => "11000000",2921 => "01010011",2922 => "01000010",2923 => "10001111",2924 => "01101100",2925 => "01100101",2926 => "00001001",2927 => "01000101",2928 => "01000011",2929 => "10000011",2930 => "01100011",2931 => "00110100",2932 => "11101111",2933 => "11100101",2934 => "11100101",2935 => "01001000",2936 => "10011000",2937 => "01110100",2938 => "11001110",2939 => "00101001",2940 => "00010101",2941 => "11110010",2942 => "01110110",2943 => "11100100",2944 => "01101111",2945 => "11101101",2946 => "01010001",2947 => "11010100",2948 => "11100110",2949 => "00011011",2950 => "10111001",2951 => "11011010",2952 => "01100101",2953 => "11001100",2954 => "01110000",2955 => "00100011",2956 => "11100001",2957 => "10000100",2958 => "00101011",2959 => "01010001",2960 => "01111110",2961 => "10011010",2962 => "11111001",2963 => "10111000",2964 => "00001001",2965 => "01111101",2966 => "00010111",2967 => "01011011",2968 => "11101000",2969 => "11110000",2970 => "01111001",2971 => "00000111",2972 => "00111101",2973 => "00111110",2974 => "10110001",2975 => "00000101",2976 => "00011100",2977 => "10000101",2978 => "10000000",2979 => "10010111",2980 => "10101111",2981 => "01111000",2982 => "11101001",2983 => "10011111",2984 => "01110100",2985 => "11010011",2986 => "10000010",2987 => "00111011",2988 => "11100001",2989 => "01010010",2990 => "01001011",2991 => "11110001",2992 => "11101110",2993 => "11000111",2994 => "10001000",2995 => "00111110",2996 => "01001101",2997 => "01111000",2998 => "10100101",2999 => "00011011",3000 => "11110101",3001 => "01100111",3002 => "01100100",3003 => "01110000",3004 => "01010100",3005 => "10011111",3006 => "00000011",3007 => "01010111",3008 => "10010010",3009 => "11101100",3010 => "00100111",3011 => "10010000",3012 => "01110110",3013 => "01011111",3014 => "00011110",3015 => "01111111",3016 => "10011110",3017 => "10010110",3018 => "01101010",3019 => "10100100",3020 => "11001011",3021 => "10001100",3022 => "11011100",3023 => "10011001",3024 => "01011101",3025 => "00110001",3026 => "00011110",3027 => "11110110",3028 => "11100101",3029 => "10101110",3030 => "11000001",3031 => "10000001",3032 => "00010001",3033 => "10010100",3034 => "11001101",3035 => "01000110",3036 => "01010001",3037 => "11111101",3038 => "10000011",3039 => "00010001",3040 => "00110110",3041 => "11100010",3042 => "11101001",3043 => "11100010",3044 => "11011010",3045 => "01010000",3046 => "11101100",3047 => "10010100",3048 => "10100100",3049 => "01110010",3050 => "00111111",3051 => "11001000",3052 => "11001111",3053 => "00011110",3054 => "11001110",3055 => "10100110",3056 => "10001001",3057 => "00110001",3058 => "01001000",3059 => "10011100",3060 => "11000010",3061 => "01001100",3062 => "11000101",3063 => "00100111",3064 => "11011110",3065 => "10111110",3066 => "01110100",3067 => "00000111",3068 => "00100111",3069 => "00110001",3070 => "01000111",3071 => "01001100",3072 => "01000111",3073 => "01100101",3074 => "00010101",3075 => "10110001",3076 => "01111011",3077 => "01111000",3078 => "10000011",3079 => "00101100",3080 => "11101110",3081 => "11110100",3082 => "11001110",3083 => "11010010",3084 => "10011011",3085 => "00011001",3086 => "11111011",3087 => "00011111",3088 => "00100100",3089 => "00100101",3090 => "11100011",3091 => "10011110",3092 => "10011010",3093 => "00100001",3094 => "11111010",3095 => "11100000",3096 => "11101010",3097 => "00010111",3098 => "01100001",3099 => "00000000",3100 => "01110110",3101 => "00100000",3102 => "10010010",3103 => "11010110",3104 => "11011110",3105 => "11010101",3106 => "01001101",3107 => "01110101",3108 => "10100100",3109 => "00110001",3110 => "01100101",3111 => "11111011",3112 => "11001001",3113 => "00000000",3114 => "10011000",3115 => "11000111",3116 => "11111110",3117 => "10111000",3118 => "11001100",3119 => "00111101",3120 => "00101011",3121 => "00011111",3122 => "11111011",3123 => "01101011",3124 => "11100100",3125 => "01110001",3126 => "00110000",3127 => "10000101",3128 => "11000010",3129 => "10010000",3130 => "00010111",3131 => "01100101",3132 => "00000001",3133 => "11100011",3134 => "00000010",3135 => "10111010",3136 => "11010000",3137 => "10101011",3138 => "00000100",3139 => "11011100",3140 => "00000011",3141 => "01001100",3142 => "01110100",3143 => "01110000",3144 => "11100100",3145 => "10110110",3146 => "11111111",3147 => "11110100",3148 => "01011100",3149 => "10001100",3150 => "10011110",3151 => "01110011",3152 => "11111101",3153 => "00111100",3154 => "11101011",3155 => "10101011",3156 => "11000011",3157 => "00100100",3158 => "01101100",3159 => "10011111",3160 => "00010001",3161 => "00110101",3162 => "01011100",3163 => "01101101",3164 => "11001010",3165 => "01010000",3166 => "00100010",3167 => "01010110",3168 => "00001110",3169 => "00100100",3170 => "10111010",3171 => "01010010",3172 => "10010000",3173 => "01001110",3174 => "01001101",3175 => "01101001",3176 => "00011011",3177 => "10110110",3178 => "00101110",3179 => "01101010",3180 => "00001101",3181 => "01001011",3182 => "00101111",3183 => "01110101",3184 => "10011100",3185 => "11001100",3186 => "01000001",3187 => "01110011",3188 => "01010010",3189 => "10100011",3190 => "01100101",3191 => "01010111",3192 => "00110110",3193 => "01000000",3194 => "00101101",3195 => "00011011",3196 => "01101111",3197 => "01011011",3198 => "10101000",3199 => "10000110",3200 => "11010011",3201 => "00000111",3202 => "11010110",3203 => "11011101",3204 => "10101100",3205 => "10100110",3206 => "11110110",3207 => "11011010",3208 => "00100100",3209 => "01101110",3210 => "01110111",3211 => "01110110",3212 => "00101000",3213 => "11010010",3214 => "11111000",3215 => "01000100",3216 => "11111101",3217 => "00110100",3218 => "01000110",3219 => "10010000",3220 => "01010011",3221 => "11111011",3222 => "10111100",3223 => "01010101",3224 => "01001010",3225 => "00000000",3226 => "01000111",3227 => "10101110",3228 => "01011111",3229 => "10010011",3230 => "10110111",3231 => "10001001",3232 => "00100111",3233 => "10100101",3234 => "10101001",3235 => "00000110",3236 => "11000100",3237 => "01000000",3238 => "11001101",3239 => "01010010",3240 => "00110111",3241 => "10110101",3242 => "10111111",3243 => "10101011",3244 => "10100001",3245 => "10101111",3246 => "10100010",3247 => "10001100",3248 => "11000101",3249 => "10111110",3250 => "00001010",3251 => "01000001",3252 => "11101011",3253 => "01011100",3254 => "00111100",3255 => "00100010",3256 => "00101000",3257 => "10010010",3258 => "11111110",3259 => "00100001",3260 => "11001100",3261 => "01010111",3262 => "01011101",3263 => "10100110",3264 => "11111110",3265 => "01010110",3266 => "10001110",3267 => "01111101",3268 => "01010000",3269 => "01100111",3270 => "00010100",3271 => "01000010",3272 => "10101010",3273 => "10010110",3274 => "11011010",3275 => "11011111",3276 => "00110011",3277 => "11000101",3278 => "10010001",3279 => "00101010",3280 => "01110011",3281 => "11111010",3282 => "00111111",3283 => "10111010",3284 => "10011011",3285 => "11010100",3286 => "01011001",3287 => "01010011",3288 => "00000001",3289 => "11100101",3290 => "00111111",3291 => "11010011",3292 => "00101101",3293 => "10110001",3294 => "10110101",3295 => "01010110",3296 => "01110101",3297 => "00000101",3298 => "11011010",3299 => "01001000",3300 => "11010011",3301 => "00100000",3302 => "10001111",3303 => "00111010",3304 => "01100100",3305 => "00111010",3306 => "10111001",3307 => "00101011",3308 => "00010011",3309 => "11101010",3310 => "11011101",3311 => "11101010",3312 => "11110011",3313 => "10110010",3314 => "01101011",3315 => "01111000",3316 => "01011110",3317 => "01111000",3318 => "00000110",3319 => "00011011",3320 => "00101010",3321 => "10010010",3322 => "01100011",3323 => "11000110",3324 => "10100100",3325 => "01101000",3326 => "00100011",3327 => "01110111",3328 => "10110100",3329 => "10101001",3330 => "11101011",3331 => "11001100",3332 => "01001000",3333 => "00011101",3334 => "00100100",3335 => "10101001",3336 => "11001001",3337 => "10111010",3338 => "11111111",3339 => "01000010",3340 => "10101110",3341 => "00011101",3342 => "11010011",3343 => "10111111",3344 => "10011011",3345 => "00011101",3346 => "01101001",3347 => "01010010",3348 => "01010100",3349 => "01000000",3350 => "00110000",3351 => "11111111",3352 => "10110001",3353 => "11100110",3354 => "10010011",3355 => "01001011",3356 => "11011111",3357 => "00010011",3358 => "01100000",3359 => "01110011",3360 => "10111011",3361 => "10101000",3362 => "11001000",3363 => "01111110",3364 => "01110001",3365 => "10001010",3366 => "10010110",3367 => "00000100",3368 => "10010000",3369 => "11100111",3370 => "11001111",3371 => "10010001",3372 => "01101100",3373 => "10110100",3374 => "11110000",3375 => "10111111",3376 => "10000100",3377 => "11010011",3378 => "11100000",3379 => "10000001",3380 => "10110100",3381 => "10100100",3382 => "10011101",3383 => "00011011",3384 => "11111010",3385 => "10100000",3386 => "11110110",3387 => "00111010",3388 => "00001010",3389 => "01111100",3390 => "11110010",3391 => "01010111",3392 => "00110111",3393 => "01011111",3394 => "00010110",3395 => "00011010",3396 => "10111110",3397 => "11110100",3398 => "10010011",3399 => "01100101",3400 => "11001111",3401 => "11100111",3402 => "10011000",3403 => "11011100",3404 => "10000100",3405 => "10100000",3406 => "00101110",3407 => "00110100",3408 => "01010011",3409 => "01011111",3410 => "01100001",3411 => "11001011",3412 => "01101110",3413 => "00111010",3414 => "11100011",3415 => "11111000",3416 => "11010101",3417 => "11111011",3418 => "00011111",3419 => "11000100",3420 => "11110010",3421 => "00101110",3422 => "10100010",3423 => "01010001",3424 => "01010101",3425 => "00001000",3426 => "10000010",3427 => "11111111",3428 => "10101110",3429 => "11100010",3430 => "00111010",3431 => "01001001",3432 => "11100110",3433 => "10110000",3434 => "10101001",3435 => "01100000",3436 => "01100011",3437 => "10111000",3438 => "00101110",3439 => "00010011",3440 => "01111011",3441 => "11111110",3442 => "11100010",3443 => "00101000",3444 => "11000111",3445 => "01001111",3446 => "01000001",3447 => "11000101",3448 => "00011111",3449 => "01001110",3450 => "01110100",3451 => "01111010",3452 => "00101110",3453 => "11111110",3454 => "00100101",3455 => "00101001",3456 => "00110011",3457 => "11010011",3458 => "00101101",3459 => "01100100",3460 => "00001010",3461 => "01011100",3462 => "10111001",3463 => "00001011",3464 => "01111000",3465 => "10100001",3466 => "01100101",3467 => "00111100",3468 => "10111110",3469 => "01010101",3470 => "11110010",3471 => "10111010",3472 => "01111001",3473 => "01110110",3474 => "01010011",3475 => "10010010",3476 => "01100010",3477 => "00000001",3478 => "00010101",3479 => "11110111",3480 => "01000101",3481 => "11001110",3482 => "00110110",3483 => "10000101",3484 => "01000001",3485 => "10111011",3486 => "01010001",3487 => "11101001",3488 => "10111100",3489 => "01111111",3490 => "00011110",3491 => "10010100",3492 => "11001101",3493 => "01100100",3494 => "11110110",3495 => "11100110",3496 => "11110101",3497 => "01100100",3498 => "01111110",3499 => "00100111",3500 => "01111110",3501 => "11000010",3502 => "10010101",3503 => "10010000",3504 => "10111110",3505 => "11001100",3506 => "00011000",3507 => "11100111",3508 => "11100000",3509 => "11110011",3510 => "01011100",3511 => "10000110",3512 => "01100100",3513 => "01001111",3514 => "01111001",3515 => "00110111",3516 => "00000110",3517 => "10111110",3518 => "11111001",3519 => "11110100",3520 => "11010111",3521 => "11011110",3522 => "10100010",3523 => "01010000",3524 => "00101011",3525 => "11001110",3526 => "11001101",3527 => "00110000",3528 => "11000100",3529 => "10111000",3530 => "00000110",3531 => "11100100",3532 => "11101011",3533 => "11011010",3534 => "01111011",3535 => "01100101",3536 => "01000111",3537 => "00000110",3538 => "10001101",3539 => "11100001",3540 => "11101111",3541 => "10110001",3542 => "10011111",3543 => "11000101",3544 => "10111000",3545 => "01100100",3546 => "00100000",3547 => "10100000",3548 => "00010010",3549 => "00010000",3550 => "00110110",3551 => "11111000",3552 => "10000010",3553 => "11100000",3554 => "11101110",3555 => "11001101",3556 => "11110110",3557 => "10000101",3558 => "00110111",3559 => "00010111",3560 => "11101011",3561 => "00111101",3562 => "00110011",3563 => "00010100",3564 => "10010100",3565 => "00101110",3566 => "01111111",3567 => "11101001",3568 => "11110110",3569 => "01111011",3570 => "01000101",3571 => "00110111",3572 => "11110000",3573 => "11010101",3574 => "11110111",3575 => "11100001",3576 => "10100000",3577 => "01111100",3578 => "11101101",3579 => "10110110",3580 => "01100011",3581 => "10000000",3582 => "11100000",3583 => "01101110",3584 => "00011101",3585 => "11001010",3586 => "01001111",3587 => "01110000",3588 => "11011011",3589 => "11100000",3590 => "01010001",3591 => "11111011",3592 => "00011011",3593 => "11111111",3594 => "00001010",3595 => "11001001",3596 => "11010101",3597 => "11001000",3598 => "10001001",3599 => "01001011",3600 => "11001011",3601 => "01001100",3602 => "01011101",3603 => "00101110",3604 => "10001101",3605 => "01000000",3606 => "00011001",3607 => "00100001",3608 => "01000101",3609 => "00000100",3610 => "00101100",3611 => "11100011",3612 => "11011010",3613 => "00101001",3614 => "00010001",3615 => "10111100",3616 => "10100110",3617 => "10011100",3618 => "01101111",3619 => "00111111",3620 => "11101001",3621 => "01110111",3622 => "10010100",3623 => "01110110",3624 => "00000010",3625 => "01110101",3626 => "00111110",3627 => "00100001",3628 => "01111100",3629 => "00101000",3630 => "01000100",3631 => "10010001",3632 => "00101111",3633 => "11001100",3634 => "00100010",3635 => "01110110",3636 => "00100010",3637 => "10000010",3638 => "01110110",3639 => "00111110",3640 => "00110100",3641 => "10011001",3642 => "10100001",3643 => "10011010",3644 => "11010000",3645 => "00010100",3646 => "10100011",3647 => "00010011",3648 => "10001110",3649 => "01001100",3650 => "01000010",3651 => "11100111",3652 => "10011000",3653 => "11101000",3654 => "10000010",3655 => "00001101",3656 => "01011100",3657 => "01010111",3658 => "01010101",3659 => "11010001",3660 => "11001000",3661 => "00110101",3662 => "11100110",3663 => "00011010",3664 => "01100111",3665 => "10111111",3666 => "00110011",3667 => "01101011",3668 => "10100111",3669 => "00111101",3670 => "10010110",3671 => "11101010",3672 => "10001101",3673 => "00101100",3674 => "10010101",3675 => "11011011",3676 => "11101110",3677 => "11010010",3678 => "00011100",3679 => "00000110",3680 => "00110010",3681 => "11111010",3682 => "01011110",3683 => "00100101",3684 => "10111101",3685 => "10010011",3686 => "00111101",3687 => "11000100",3688 => "10101101",3689 => "10110111",3690 => "01011010",3691 => "11001101",3692 => "01110101",3693 => "11000111",3694 => "01011100",3695 => "10010101",3696 => "01001010",3697 => "11110000",3698 => "11001011",3699 => "11011110",3700 => "00110010",3701 => "10101111",3702 => "01111101",3703 => "10010001",3704 => "01010001",3705 => "00001001",3706 => "01111101",3707 => "10001000",3708 => "11111111",3709 => "10111111",3710 => "10011100",3711 => "01010101",3712 => "10111100",3713 => "11111101",3714 => "01011110",3715 => "01101001",3716 => "00111001",3717 => "10111000",3718 => "00111010",3719 => "00110000",3720 => "00001011",3721 => "10110011",3722 => "01101010",3723 => "01000111",3724 => "10101101",3725 => "01001101",3726 => "00010010",3727 => "11011101",3728 => "11111000",3729 => "10001011",3730 => "00000111",3731 => "11001111",3732 => "10101011",3733 => "00101101",3734 => "11011100",3735 => "10001111",3736 => "01001100",3737 => "01001110",3738 => "11100001",3739 => "01000110",3740 => "10111101",3741 => "01110011",3742 => "10000000",3743 => "10100001",3744 => "11010111",3745 => "00001111",3746 => "01101000",3747 => "11101100",3748 => "00101011",3749 => "10111110",3750 => "11000110",3751 => "10001101",3752 => "11010010",3753 => "11100000",3754 => "11111010",3755 => "01110101",3756 => "11111001",3757 => "00010001",3758 => "10111000",3759 => "10101100",3760 => "01111110",3761 => "10000000",3762 => "01110010",3763 => "00110010",3764 => "01001101",3765 => "01011111",3766 => "01000001",3767 => "01010000",3768 => "01010101",3769 => "11110000",3770 => "01000000",3771 => "00010110",3772 => "11001101",3773 => "00010111",3774 => "00011000",3775 => "01001000",3776 => "01001010",3777 => "10011010",3778 => "10001010",3779 => "10100000",3780 => "10001110",3781 => "10111000",3782 => "01000110",3783 => "00100010",3784 => "11010010",3785 => "10110101",3786 => "01010001",3787 => "00011001",3788 => "11100111",3789 => "01001000",3790 => "11000001",3791 => "00000010",3792 => "11100110",3793 => "01001000",3794 => "11000001",3795 => "11001011",3796 => "01110010",3797 => "01110110",3798 => "01000111",3799 => "00111010",3800 => "01010000",3801 => "00000100",3802 => "11010111",3803 => "10011010",3804 => "11001000",3805 => "11111000",3806 => "00110000",3807 => "11011011",3808 => "01100011",3809 => "00111110",3810 => "11100000",3811 => "11110011",3812 => "10110111",3813 => "10011010",3814 => "10001000",3815 => "10100101",3816 => "01101011",3817 => "11110111",3818 => "11010011",3819 => "11001101",3820 => "00101100",3821 => "01001011",3822 => "00110010",3823 => "11110110",3824 => "11110011",3825 => "01110001",3826 => "01110111",3827 => "01111101",3828 => "01100111",3829 => "00001000",3830 => "01111010",3831 => "11110101",3832 => "01010101",3833 => "01110100",3834 => "00101011",3835 => "00100001",3836 => "01110100",3837 => "11010000",3838 => "00000111",3839 => "11101011",3840 => "01010001",3841 => "01000011",3842 => "11101111",3843 => "11010101",3844 => "10000110",3845 => "01010100",3846 => "01100001",3847 => "00011001",3848 => "01101101",3849 => "10100111",3850 => "11100010",3851 => "00001010",3852 => "01111000",3853 => "00110010",3854 => "11011001",3855 => "00101000",3856 => "11001100",3857 => "00011110",3858 => "11011001",3859 => "11011110",3860 => "10100001",3861 => "11011110",3862 => "01010100",3863 => "11110110",3864 => "11000000",3865 => "00101101",3866 => "00111101",3867 => "11011110",3868 => "11110100",3869 => "11101000",3870 => "00111111",3871 => "11001000",3872 => "00001100",3873 => "11111001",3874 => "11111110",3875 => "10000011",3876 => "00111100",3877 => "00000110",3878 => "00011111",3879 => "00110011",3880 => "11010010",3881 => "11010010",3882 => "10111110",3883 => "11100111",3884 => "00100110",3885 => "00100101",3886 => "01000111",3887 => "11000110",3888 => "10100000",3889 => "10100100",3890 => "11010101",3891 => "10000001",3892 => "11010101",3893 => "10110001",3894 => "11011001",3895 => "00000001",3896 => "01101111",3897 => "10100100",3898 => "01001101",3899 => "00100000",3900 => "11111010",3901 => "11010111",3902 => "01100111",3903 => "10100110",3904 => "10001000",3905 => "00010000",3906 => "10110011",3907 => "00010110",3908 => "10010011",3909 => "01000100",3910 => "10001100",3911 => "01001011",3912 => "10010110",3913 => "00011000",3914 => "00011001",3915 => "01101100",3916 => "11011000",3917 => "11011110",3918 => "11100110",3919 => "10110110",3920 => "00100001",3921 => "11000001",3922 => "00110110",3923 => "10110001",3924 => "01001010",3925 => "01100001",3926 => "00100011",3927 => "00010100",3928 => "00110010",3929 => "01000000",3930 => "01010011",3931 => "00011001",3932 => "01010110",3933 => "11101001",3934 => "01101100",3935 => "11010101",3936 => "11101101",3937 => "01101110",3938 => "01010010",3939 => "10111001",3940 => "10010001",3941 => "11000011",3942 => "00011011",3943 => "00111000",3944 => "11101111",3945 => "11101011",3946 => "10100001",3947 => "01111101",3948 => "00001111",3949 => "01010011",3950 => "01000001",3951 => "11010111",3952 => "11010111",3953 => "00111110",3954 => "10111100",3955 => "11011000",3956 => "11001010",3957 => "00100001",3958 => "00111101",3959 => "10111100",3960 => "11010001",3961 => "01000000",3962 => "00101101",3963 => "01110111",3964 => "11011000",3965 => "11111101",3966 => "01111011",3967 => "11111001",3968 => "00011001",3969 => "01001000",3970 => "01011001",3971 => "11110110",3972 => "11100111",3973 => "01111011",3974 => "00001100",3975 => "00101011",3976 => "10001110",3977 => "00011000",3978 => "01010010",3979 => "00001010",3980 => "11001100",3981 => "11101100",3982 => "00100111",3983 => "00110101",3984 => "10001110",3985 => "11011100",3986 => "01000000",3987 => "01010001",3988 => "00011100",3989 => "11001100",3990 => "01000100",3991 => "11110000",3992 => "11010111",3993 => "00111011",3994 => "10010111",3995 => "00001001",3996 => "00100110",3997 => "00011101",3998 => "01111100",3999 => "10111010",4000 => "10100000",4001 => "11011011",4002 => "11011011",4003 => "00101100",4004 => "01001101",4005 => "01110100",4006 => "01111100",4007 => "10011111",4008 => "01100000",4009 => "00110100",4010 => "01010111",4011 => "01001110",4012 => "01000010",4013 => "01001100",4014 => "10101100",4015 => "10110110",4016 => "00000101",4017 => "00101011",4018 => "01111100",4019 => "10111001",4020 => "01010010",4021 => "11001100",4022 => "00010011",4023 => "01001011",4024 => "01111001",4025 => "10101101",4026 => "00011001",4027 => "11000100",4028 => "01111110",4029 => "01101101",4030 => "01110011",4031 => "10000000",4032 => "00010010",4033 => "11100001",4034 => "01111111",4035 => "01111101",4036 => "11100100",4037 => "01011010",4038 => "00100110",4039 => "11100101",4040 => "11000110",4041 => "10111001",4042 => "10110010",4043 => "00010010",4044 => "11111100",4045 => "11011011",4046 => "00011011",4047 => "01111000",4048 => "00000000",4049 => "10110100",4050 => "11110110",4051 => "11110100",4052 => "00111011",4053 => "10001011",4054 => "01110100",4055 => "01001111",4056 => "11000001",4057 => "11100111",4058 => "10110011",4059 => "11001001",4060 => "01001111",4061 => "01101110",4062 => "11110010",4063 => "00110011",4064 => "11110011",4065 => "10100111",4066 => "11010110",4067 => "11110110",4068 => "11011111",4069 => "00010000",4070 => "00101111",4071 => "10010000",4072 => "11110001",4073 => "10000111",4074 => "00100011",4075 => "00010010",4076 => "00110000",4077 => "11000111",4078 => "00000001",4079 => "01000100",4080 => "11110111",4081 => "01111101",4082 => "11000000",4083 => "11101100",4084 => "01001111",4085 => "11000011",4086 => "01111100",4087 => "10000101",4088 => "11111010",4089 => "11100001",4090 => "10100001",4091 => "00101011",4092 => "10001111",4093 => "01010001",4094 => "00111001",4095 => "00111110",4096 => "01100100",4097 => "01010110",4098 => "11000001",4099 => "01111111",4100 => "01101011",4101 => "11100111",4102 => "01111101",4103 => "10101000",4104 => "01001000",4105 => "11110011",4106 => "01100011",4107 => "10001101",4108 => "01010010",4109 => "00100111",4110 => "11101111",4111 => "01100101",4112 => "00100101",4113 => "11010100",4114 => "00110110",4115 => "00101101",4116 => "10111111",4117 => "10110011",4118 => "00010110",4119 => "11010011",4120 => "10010000",4121 => "00011110",4122 => "11011011",4123 => "10101111",4124 => "01111110",4125 => "10111111",4126 => "01000010",4127 => "00101101",4128 => "00010000",4129 => "11100011",4130 => "10101101",4131 => "10111001",4132 => "10010001",4133 => "10111010",4134 => "00010011",4135 => "00000011",4136 => "10100010",4137 => "00010000",4138 => "11001000",4139 => "11101000",4140 => "11110100",4141 => "11000011",4142 => "10001110",4143 => "00001110",4144 => "01000011",4145 => "01111001",4146 => "11101100",4147 => "10100110",4148 => "11100101",4149 => "00110001",4150 => "00110100",4151 => "10111010",4152 => "00010000",4153 => "11001011",4154 => "11011110",4155 => "01110000",4156 => "00000011",4157 => "00100001",4158 => "01000010",4159 => "10001101",4160 => "01001000",4161 => "00101101",4162 => "11011011",4163 => "01100101",4164 => "11100111",4165 => "00111010",4166 => "00011101",4167 => "01001010",4168 => "01101111",4169 => "11100101",4170 => "00110110",4171 => "11000011",4172 => "01001010",4173 => "00101110",4174 => "11011010",4175 => "01100000",4176 => "11000111",4177 => "01101010",4178 => "00000011",4179 => "00111101",4180 => "10011010",4181 => "00011010",4182 => "10000111",4183 => "11101000",4184 => "01110000",4185 => "10101110",4186 => "01100111",4187 => "01101011",4188 => "00010010",4189 => "10000111",4190 => "00100100",4191 => "11110110",4192 => "11011101",4193 => "11111011",4194 => "10111101",4195 => "00010100",4196 => "01100100",4197 => "01111001",4198 => "11101100",4199 => "11000100",4200 => "10000011",4201 => "10100011",4202 => "01111010",4203 => "01011001",4204 => "11011100",4205 => "10011110",4206 => "00010110",4207 => "01110010",4208 => "10011011",4209 => "10001100",4210 => "00100110",4211 => "00010111",4212 => "01011110",4213 => "01011111",4214 => "11001100",4215 => "01110111",4216 => "00001100",4217 => "01101111",4218 => "01110111",4219 => "10101001",4220 => "01111110",4221 => "11010111",4222 => "00011110",4223 => "11011000",4224 => "01001101",4225 => "00100000",4226 => "00001110",4227 => "10001001",4228 => "01010001",4229 => "01011110",4230 => "01001001",4231 => "01110010",4232 => "01110011",4233 => "01110001",4234 => "01000101",4235 => "01011101",4236 => "00011110",4237 => "01011001",4238 => "00111110",4239 => "01010000",4240 => "11011010",4241 => "11101001",4242 => "10111111",4243 => "11100000",4244 => "00010101",4245 => "01001100",4246 => "11010001",4247 => "10000100",4248 => "01100010",4249 => "10001101",4250 => "11111001",4251 => "11000010",4252 => "01010001",4253 => "10011111",4254 => "01100000",4255 => "01110000",4256 => "00101000",4257 => "10100000",4258 => "10110100",4259 => "01001110",4260 => "01101111",4261 => "01011001",4262 => "01111001",4263 => "11011001",4264 => "01010111",4265 => "10100011",4266 => "10111111",4267 => "00001011",4268 => "10000101",4269 => "01101101",4270 => "01110011",4271 => "11100011",4272 => "00000010",4273 => "00011000",4274 => "10101010",4275 => "10011110",4276 => "00110110",4277 => "11001110",4278 => "00000011",4279 => "00001100",4280 => "10001010",4281 => "00110111",4282 => "01110111",4283 => "01001110",4284 => "01010111",4285 => "00111111",4286 => "01111100",4287 => "11011000",4288 => "10100010",4289 => "00000110",4290 => "11000001",4291 => "01111000",4292 => "10010110",4293 => "01001001",4294 => "00010010",4295 => "10010101",4296 => "11111100",4297 => "00111001",4298 => "01010110",4299 => "11111001",4300 => "00000011",4301 => "01110000",4302 => "01011000",4303 => "00110100",4304 => "11101010",4305 => "00001010",4306 => "11011000",4307 => "10001101",4308 => "10001110",4309 => "01000000",4310 => "00110000",4311 => "10001111",4312 => "00110000",4313 => "00111001",4314 => "11100110",4315 => "00001001",4316 => "10110111",4317 => "10101101",4318 => "00111001",4319 => "00110000",4320 => "01010010",4321 => "00100010",4322 => "00011101",4323 => "10101001",4324 => "00101111",4325 => "11100001",4326 => "11100100",4327 => "00100000",4328 => "11100011",4329 => "10101001",4330 => "01100011",4331 => "01110110",4332 => "10000011",4333 => "00111101",4334 => "11010000",4335 => "01100110",4336 => "00111100",4337 => "00101101",4338 => "00011101",4339 => "01100111",4340 => "00111011",4341 => "01110111",4342 => "11010100",4343 => "01111111",4344 => "11010101",4345 => "11111000",4346 => "10101011",4347 => "10011101",4348 => "10100011",4349 => "01010001",4350 => "11111101",4351 => "11000001",4352 => "10110011",4353 => "11000101",4354 => "11111011",4355 => "01001101",4356 => "10000010",4357 => "00111101",4358 => "00100100",4359 => "11100011",4360 => "00100101",4361 => "10000101",4362 => "11101110",4363 => "00011110",4364 => "00010000",4365 => "10110001",4366 => "00101100",4367 => "00011010",4368 => "10101010",4369 => "00101000",4370 => "10010101",4371 => "11011110",4372 => "01001111",4373 => "10111000",4374 => "10101111",4375 => "11001111",4376 => "01010111",4377 => "00001110",4378 => "10101001",4379 => "00010101",4380 => "10010011",4381 => "01011001",4382 => "00010000",4383 => "10001100",4384 => "00110100",4385 => "00000010",4386 => "11010101",4387 => "10011110",4388 => "11001011",4389 => "00101001",4390 => "00110111",4391 => "00001011",4392 => "00100101",4393 => "00011110",4394 => "01001001",4395 => "11011101",4396 => "00001101",4397 => "11101010",4398 => "10110010",4399 => "10100011",4400 => "00101100",4401 => "00000010",4402 => "00100011",4403 => "10010111",4404 => "10000010",4405 => "01110010",4406 => "01101111",4407 => "01000001",4408 => "10101110",4409 => "11110111",4410 => "01111010",4411 => "10100010",4412 => "10101000",4413 => "00111000",4414 => "10111010",4415 => "11101000",4416 => "10101101",4417 => "10011110",4418 => "10000011",4419 => "10001100",4420 => "10110111",4421 => "11000100",4422 => "01010011",4423 => "01001100",4424 => "00000111",4425 => "01100011",4426 => "01011110",4427 => "11110110",4428 => "10011101",4429 => "11001101",4430 => "10000010",4431 => "00110011",4432 => "10001100",4433 => "11111011",4434 => "01001011",4435 => "10100001",4436 => "01101111",4437 => "01100100",4438 => "00001000",4439 => "01100000",4440 => "11000000",4441 => "10101110",4442 => "10100000",4443 => "00100010",4444 => "10101100",4445 => "10111101",4446 => "10111101",4447 => "10110011",4448 => "11010001",4449 => "01110011",4450 => "10111010",4451 => "11010001",4452 => "01010001",4453 => "01000111",4454 => "01010111",4455 => "01001001",4456 => "11011011",4457 => "01101010",4458 => "00111011",4459 => "10001001",4460 => "11010101",4461 => "00101111",4462 => "10100111",4463 => "00111110",4464 => "11100011",4465 => "10000101",4466 => "11101111",4467 => "01000011",4468 => "11101010",4469 => "00011000",4470 => "00001010",4471 => "00111100",4472 => "11101011",4473 => "10001111",4474 => "01100110",4475 => "10001011",4476 => "01000011",4477 => "01010000",4478 => "01011100",4479 => "01001111",4480 => "01101010",4481 => "11010001",4482 => "00010010",4483 => "00010010",4484 => "00101101",4485 => "10101010",4486 => "01011010",4487 => "10000101",4488 => "11011110",4489 => "11010100",4490 => "11110101",4491 => "10011100",4492 => "11000001",4493 => "01010100",4494 => "10100101",4495 => "11001101",4496 => "11100111",4497 => "01011100",4498 => "01000110",4499 => "10001110",4500 => "00101101",4501 => "01110010",4502 => "01100001",4503 => "11100100",4504 => "10110111",4505 => "01001000",4506 => "00111011",4507 => "11111010",4508 => "01001001",4509 => "11010101",4510 => "10111001",4511 => "10001110",4512 => "00110011",4513 => "11000011",4514 => "01001011",4515 => "01001000",4516 => "10000101",4517 => "01101110",4518 => "00111011",4519 => "00111001",4520 => "11010111",4521 => "11100111",4522 => "11100100",4523 => "11010001",4524 => "01011110",4525 => "10111101",4526 => "10110111",4527 => "10001001",4528 => "11110011",4529 => "00100000",4530 => "00000111",4531 => "00101011",4532 => "00101111",4533 => "10010001",4534 => "10100010",4535 => "11100010",4536 => "00001110",4537 => "11110000",4538 => "11110101",4539 => "01001110",4540 => "00100101",4541 => "00100000",4542 => "00001110",4543 => "01011000",4544 => "10000100",4545 => "00111011",4546 => "01010010",4547 => "11001110",4548 => "10000110",4549 => "00000011",4550 => "01100100",4551 => "01101000",4552 => "01101110",4553 => "10111110",4554 => "00011101",4555 => "01101101",4556 => "00100001",4557 => "01000000",4558 => "01011111",4559 => "10010100",4560 => "10010011",4561 => "00010010",4562 => "11100110",4563 => "00110011",4564 => "11010010",4565 => "01100000",4566 => "10010100",4567 => "10110001",4568 => "11110101",4569 => "00101000",4570 => "10110111",4571 => "10001000",4572 => "01101001",4573 => "01000111",4574 => "00110001",4575 => "00100000",4576 => "10111101",4577 => "01110110",4578 => "10101011",4579 => "00110101",4580 => "01110100",4581 => "11101111",4582 => "01000011",4583 => "11100010",4584 => "00011110",4585 => "01001110",4586 => "10001100",4587 => "10010000",4588 => "11011000",4589 => "00111011",4590 => "10011001",4591 => "01001000",4592 => "00000110",4593 => "00101111",4594 => "00111010",4595 => "01111100",4596 => "00101100",4597 => "10101101",4598 => "10001001",4599 => "11010101",4600 => "01101111",4601 => "11000101",4602 => "10001010",4603 => "11110010",4604 => "01101010",4605 => "01001100",4606 => "00100011",4607 => "01000110",4608 => "11000010",4609 => "10000011",4610 => "01111001",4611 => "01100110",4612 => "00111001",4613 => "01111101",4614 => "11011111",4615 => "00001011",4616 => "00000100",4617 => "00101100",4618 => "01010001",4619 => "11000001",4620 => "00011110",4621 => "10100110",4622 => "01100001",4623 => "11011110",4624 => "11111001",4625 => "01100000",4626 => "11000101",4627 => "01000100",4628 => "00111101",4629 => "00101110",4630 => "10110011",4631 => "10010111",4632 => "10011000",4633 => "11001110",4634 => "11010111",4635 => "00110010",4636 => "01000111",4637 => "11000110",4638 => "01111101",4639 => "01011111",4640 => "00100011",4641 => "11011001",4642 => "01111111",4643 => "01111110",4644 => "10001100",4645 => "11001100",4646 => "11010110",4647 => "01100110",4648 => "00011111",4649 => "11000111",4650 => "11010011",4651 => "01001000",4652 => "00010100",4653 => "11101001",4654 => "11110101",4655 => "11011011",4656 => "10111001",4657 => "10010010",4658 => "01000101",4659 => "00101101",4660 => "01000111",4661 => "10011000",4662 => "10101100",4663 => "00000000",4664 => "11011111",4665 => "01100010",4666 => "01010001",4667 => "11001001",4668 => "00100000",4669 => "00111000",4670 => "00111010",4671 => "11010110",4672 => "01000011",4673 => "01011011",4674 => "00000101",4675 => "01010011",4676 => "01101001",4677 => "00110111",4678 => "01001010",4679 => "00010101",4680 => "10110010",4681 => "11111111",4682 => "00000011",4683 => "00010001",4684 => "00100101",4685 => "01110011",4686 => "00001111",4687 => "01110000",4688 => "10111011",4689 => "11110111",4690 => "10101101",4691 => "00110011",4692 => "11100110",4693 => "01110011",4694 => "00001001",4695 => "01111100",4696 => "01110110",4697 => "11101010",4698 => "00101001",4699 => "00101011",4700 => "11000011",4701 => "01111011",4702 => "10000000",4703 => "10001001",4704 => "11111001",4705 => "01000000",4706 => "00111100",4707 => "00100001",4708 => "01111010",4709 => "10101100",4710 => "10111000",4711 => "10101110",4712 => "00110110",4713 => "11000010",4714 => "11111111",4715 => "00010000",4716 => "11101100",4717 => "11110010",4718 => "01110101",4719 => "10001011",4720 => "01011101",4721 => "11001110",4722 => "10000000",4723 => "10001111",4724 => "00101010",4725 => "11100000",4726 => "00010110",4727 => "11111100",4728 => "00100110",4729 => "11111110",4730 => "10111111",4731 => "00000000",4732 => "11010000",4733 => "01111110",4734 => "01000001",4735 => "10000010",4736 => "01110110",4737 => "00000010",4738 => "10011000",4739 => "00101111",4740 => "11110011",4741 => "10000000",4742 => "10010101",4743 => "10101011",4744 => "00001000",4745 => "10011110",4746 => "00010010",4747 => "01001100",4748 => "00101000",4749 => "10010100",4750 => "00001001",4751 => "00100111",4752 => "10100011",4753 => "11011101",4754 => "00110111",4755 => "11100100",4756 => "00000110",4757 => "00010101",4758 => "00011001",4759 => "10111111",4760 => "00110011",4761 => "01000110",4762 => "11110011",4763 => "00010000",4764 => "11010000",4765 => "11100011",4766 => "01010110",4767 => "10101001",4768 => "10110100",4769 => "01111111",4770 => "01000100",4771 => "00111010",4772 => "01001010",4773 => "11111100",4774 => "01010111",4775 => "11010101",4776 => "00111110",4777 => "10101111",4778 => "11101001",4779 => "00011010",4780 => "10000000",4781 => "01100100",4782 => "01000010",4783 => "01000110",4784 => "01100000",4785 => "00000100",4786 => "10111001",4787 => "01010000",4788 => "01010010",4789 => "10001101",4790 => "10101010",4791 => "11010000",4792 => "10111010",4793 => "00000101",4794 => "00000110",4795 => "11100101",4796 => "01110111",4797 => "10111000",4798 => "11000101",4799 => "01111110",4800 => "01100101",4801 => "01111000",4802 => "11100110",4803 => "00010001",4804 => "01010101",4805 => "01111101",4806 => "10010010",4807 => "00000010",4808 => "00101010",4809 => "00000111",4810 => "11101001",4811 => "10010011",4812 => "00100000",4813 => "00111100",4814 => "00010000",4815 => "11011001",4816 => "01111111",4817 => "11100001",4818 => "00101100",4819 => "00010100",4820 => "01110101",4821 => "11010001",4822 => "01110010",4823 => "10111100",4824 => "00110101",4825 => "01111011",4826 => "10000100",4827 => "11101010",4828 => "10010000",4829 => "10011100",4830 => "00011010",4831 => "01110001",4832 => "01000010",4833 => "00011101",4834 => "11011110",4835 => "11100011",4836 => "01011001",4837 => "01111000",4838 => "00011000",4839 => "10101001",4840 => "01100110",4841 => "00000000",4842 => "11010010",4843 => "11001101",4844 => "11100110",4845 => "10011111",4846 => "00101101",4847 => "01001011",4848 => "01110000",4849 => "11001110",4850 => "10010000",4851 => "01000101",4852 => "01100001",4853 => "00001100",4854 => "00010100",4855 => "01011010",4856 => "11101000",4857 => "00101000",4858 => "00011000",4859 => "11001010",4860 => "10010011",4861 => "00100010",4862 => "11001111",4863 => "11101011",4864 => "01111001",4865 => "00010000",4866 => "01001011",4867 => "10000111",4868 => "00100001",4869 => "00011011",4870 => "01100101",4871 => "01111010",4872 => "11010000",4873 => "10100101",4874 => "10010110",4875 => "11111111",4876 => "01000110",4877 => "00011011",4878 => "00111111",4879 => "10001110",4880 => "11000111",4881 => "01000111",4882 => "01110011",4883 => "01100110",4884 => "11000000",4885 => "01100000",4886 => "11100111",4887 => "00011111",4888 => "01001100",4889 => "01110001",4890 => "10110101",4891 => "00000010",4892 => "10110001",4893 => "00100101",4894 => "01000010",4895 => "00000101",4896 => "11001100",4897 => "11100100",4898 => "10010110",4899 => "01111011",4900 => "00101100",4901 => "11010110",4902 => "10111011",4903 => "11001001",4904 => "01100000",4905 => "00100011",4906 => "01011110",4907 => "01101101",4908 => "11101101",4909 => "11000010",4910 => "01010010",4911 => "00100011",4912 => "01001010",4913 => "01010010",4914 => "10001110",4915 => "11010110",4916 => "10110000",4917 => "10101110",4918 => "01101100",4919 => "10111111",4920 => "00100100",4921 => "11011000",4922 => "01010011",4923 => "01100010",4924 => "00011011",4925 => "11110011",4926 => "01110110",4927 => "11111000",4928 => "11100101",4929 => "01111011",4930 => "01001100",4931 => "11011111",4932 => "10011010",4933 => "11100110",4934 => "11001001",4935 => "11001101",4936 => "10101110",4937 => "00111101",4938 => "01101000",4939 => "11111111",4940 => "00010100",4941 => "11010001",4942 => "10110010",4943 => "10000000",4944 => "10001101",4945 => "01101110",4946 => "00110101",4947 => "10100101",4948 => "11110100",4949 => "01100010",4950 => "01011000",4951 => "00001011",4952 => "00101001",4953 => "11001010",4954 => "00101000",4955 => "10011111",4956 => "10100011",4957 => "01111100",4958 => "11000011",4959 => "00001111",4960 => "01010111",4961 => "11000110",4962 => "00000111",4963 => "00111010",4964 => "01110101",4965 => "00000101",4966 => "11000111",4967 => "10011111",4968 => "01000000",4969 => "11111000",4970 => "11001101",4971 => "00000110",4972 => "00000010",4973 => "11100000",4974 => "10001100",4975 => "10010010",4976 => "01110111",4977 => "10001101",4978 => "11101011",4979 => "11001001",4980 => "01101000",4981 => "00010001",4982 => "00101111",4983 => "01011100",4984 => "11011010",4985 => "11101011",4986 => "10000011",4987 => "10011011",4988 => "01001010",4989 => "01010110",4990 => "00100111",4991 => "01001010",4992 => "01111110",4993 => "00000001",4994 => "10101110",4995 => "00001111",4996 => "00000001",4997 => "11100011",4998 => "01000010",4999 => "10000100",5000 => "00111111",5001 => "00110010",5002 => "10011101",5003 => "11010111",5004 => "00110000",5005 => "00010101",5006 => "11111001",5007 => "00011010",5008 => "10000110",5009 => "10100110",5010 => "11100100",5011 => "00111100",5012 => "00110000",5013 => "01001011",5014 => "11101011",5015 => "00001110",5016 => "00010000",5017 => "10111111",5018 => "00001111",5019 => "01010011",5020 => "11000101",5021 => "00111010",5022 => "01111011",5023 => "11110111",5024 => "00111001",5025 => "11100110",5026 => "10010000",5027 => "01011001",5028 => "00010110",5029 => "01010001",5030 => "01010100",5031 => "00001110",5032 => "00010110",5033 => "10001001",5034 => "00101000",5035 => "01101000",5036 => "00110100",5037 => "11101010",5038 => "11000100",5039 => "11000110",5040 => "00010101",5041 => "01010011",5042 => "10110111",5043 => "01001101",5044 => "01000011",5045 => "01011110",5046 => "00000001",5047 => "11111001",5048 => "01100010",5049 => "00011011",5050 => "10010111",5051 => "00101101",5052 => "11001010",5053 => "01100111",5054 => "00011000",5055 => "10010011",5056 => "01101111",5057 => "11101110",5058 => "11000011",5059 => "10000111",5060 => "00010111",5061 => "00001000",5062 => "11111011",5063 => "11100111",5064 => "10100111",5065 => "11010001",5066 => "11011001",5067 => "00001000",5068 => "10100010",5069 => "11000111",5070 => "01010100",5071 => "01100000",5072 => "11100011",5073 => "10011001",5074 => "01101001",5075 => "11100001",5076 => "00110100",5077 => "01000011",5078 => "10011100",5079 => "10110000",5080 => "11110010",5081 => "11011111",5082 => "11101100",5083 => "01011000",5084 => "00100000",5085 => "01000101",5086 => "11100000",5087 => "01101000",5088 => "11110101",5089 => "11001110",5090 => "01101111",5091 => "10101010",5092 => "11100001",5093 => "01000111",5094 => "10101011",5095 => "01100100",5096 => "01100001",5097 => "01111111",5098 => "01000100",5099 => "00111000",5100 => "00010110",5101 => "01101011",5102 => "10111100",5103 => "01010110",5104 => "01101111",5105 => "01010101",5106 => "11110010",5107 => "10100010",5108 => "01010001",5109 => "10100101",5110 => "01101000",5111 => "00100111",5112 => "01001001",5113 => "01010100",5114 => "00101111",5115 => "01101001",5116 => "10101001",5117 => "00001000",5118 => "01010011",5119 => "11101111",5120 => "01011101",5121 => "01001111",5122 => "11011101",5123 => "11010011",5124 => "00011110",5125 => "01100000",5126 => "11001000",5127 => "01100101",5128 => "11101100",5129 => "00101100",5130 => "01100001",5131 => "01100011",5132 => "01101011",5133 => "10101010",5134 => "00110011",5135 => "01011100",5136 => "10101001",5137 => "11011111",5138 => "01101111",5139 => "00101101",5140 => "10101110",5141 => "11111100",5142 => "01010010",5143 => "01101100",5144 => "00100000",5145 => "00110001",5146 => "01100000",5147 => "01101101",5148 => "00010101",5149 => "10011100",5150 => "11011000",5151 => "10000010",5152 => "00100100",5153 => "10000000",5154 => "11111101",5155 => "01001111",5156 => "01000111",5157 => "11101101",5158 => "11100010",5159 => "01111101",5160 => "00101000",5161 => "00100001",5162 => "10010011",5163 => "11110101",5164 => "11000111",5165 => "10100010",5166 => "10101110",5167 => "11011001",5168 => "00001100",5169 => "10010000",5170 => "01101101",5171 => "11100010",5172 => "11101110",5173 => "01111001",5174 => "01010010",5175 => "10101011",5176 => "11100110",5177 => "01011100",5178 => "11100000",5179 => "00010000",5180 => "01010010",5181 => "10000010",5182 => "11111111",5183 => "00100010",5184 => "11101110",5185 => "00001111",5186 => "00100111",5187 => "00110010",5188 => "00000101",5189 => "00000011",5190 => "10110010",5191 => "01011010",5192 => "11100000",5193 => "10101001",5194 => "00010111",5195 => "00100011",5196 => "11011101",5197 => "01001010",5198 => "00010100",5199 => "11110111",5200 => "00011010",5201 => "10000001",5202 => "00001011",5203 => "01101000",5204 => "01000110",5205 => "00011101",5206 => "00010001",5207 => "10001100",5208 => "11010010",5209 => "01100110",5210 => "01111010",5211 => "01110001",5212 => "01111101",5213 => "01000010",5214 => "10100001",5215 => "10110101",5216 => "10111100",5217 => "01111100",5218 => "10010001",5219 => "11101100",5220 => "11110100",5221 => "11110110",5222 => "01001010",5223 => "11011010",5224 => "11111010",5225 => "01001010",5226 => "11100011",5227 => "10011011",5228 => "11011111",5229 => "10001000",5230 => "00010010",5231 => "01011001",5232 => "00001111",5233 => "01000001",5234 => "00101000",5235 => "10110110",5236 => "00011110",5237 => "01011010",5238 => "01000011",5239 => "10100010",5240 => "01101000",5241 => "11011001",5242 => "10011110",5243 => "11010000",5244 => "01110100",5245 => "00110111",5246 => "01011101",5247 => "11101011",5248 => "01100001",5249 => "01100000",5250 => "00100110",5251 => "01101000",5252 => "00111010",5253 => "10001001",5254 => "01001101",5255 => "00000000",5256 => "00001011",5257 => "00101111",5258 => "01111111",5259 => "00111010",5260 => "10011100",5261 => "00101110",5262 => "11111010",5263 => "00001100",5264 => "01101101",5265 => "10011101",5266 => "01000011",5267 => "01100100",5268 => "10011101",5269 => "00000011",5270 => "00001101",5271 => "10100001",5272 => "10011101",5273 => "10011000",5274 => "10000010",5275 => "11010100",5276 => "10001101",5277 => "01110000",5278 => "01111110",5279 => "10111001",5280 => "01000001",5281 => "00110111",5282 => "11111110",5283 => "00000101",5284 => "00000011",5285 => "10100010",5286 => "11101010",5287 => "00101001",5288 => "11111111",5289 => "00000011",5290 => "01111010",5291 => "01001001",5292 => "11000111",5293 => "11111010",5294 => "10011101",5295 => "11101110",5296 => "11110100",5297 => "11110111",5298 => "11001010",5299 => "00001110",5300 => "01010011",5301 => "00110011",5302 => "11111111",5303 => "10111001",5304 => "00010111",5305 => "00110000",5306 => "10010100",5307 => "11000110",5308 => "00010010",5309 => "11011000",5310 => "10010101",5311 => "00001000",5312 => "00111001",5313 => "00011100",5314 => "00011011",5315 => "01101001",5316 => "00100011",5317 => "10100011",5318 => "01110001",5319 => "11101000",5320 => "00100100",5321 => "10110100",5322 => "00001000",5323 => "00000011",5324 => "01101011",5325 => "01001101",5326 => "00010011",5327 => "01001101",5328 => "11101001",5329 => "01101010",5330 => "10111111",5331 => "00101111",5332 => "00010101",5333 => "10000100",5334 => "11100011",5335 => "01111110",5336 => "01110011",5337 => "11100110",5338 => "11000111",5339 => "10010000",5340 => "10010110",5341 => "10100000",5342 => "11101101",5343 => "00001000",5344 => "01001000",5345 => "10101101",5346 => "11110011",5347 => "00011000",5348 => "01111110",5349 => "00000110",5350 => "11011101",5351 => "00001010",5352 => "01000110",5353 => "10110001",5354 => "10001110",5355 => "10110101",5356 => "01110100",5357 => "11000100",5358 => "01100010",5359 => "10110000",5360 => "10000101",5361 => "10011111",5362 => "11000100",5363 => "01110001",5364 => "11110010",5365 => "01100101",5366 => "00100101",5367 => "10101011",5368 => "10101110",5369 => "11100111",5370 => "01010100",5371 => "10011000",5372 => "11100101",5373 => "11100000",5374 => "00100010",5375 => "01110111",5376 => "10011110",5377 => "00101000",5378 => "10101101",5379 => "10101001",5380 => "10001101",5381 => "01100100",5382 => "01101000",5383 => "01001110",5384 => "01100110",5385 => "11110001",5386 => "10001000",5387 => "10100110",5388 => "10110011",5389 => "00101101",5390 => "11010001",5391 => "01001111",5392 => "11000111",5393 => "01001101",5394 => "00000101",5395 => "00011100",5396 => "01001111",5397 => "11011001",5398 => "01100111",5399 => "10110001",5400 => "01001110",5401 => "11100110",5402 => "10000011",5403 => "01000100",5404 => "00000000",5405 => "10111100",5406 => "00010010",5407 => "00110011",5408 => "00110111",5409 => "00100111",5410 => "00100111",5411 => "00001010",5412 => "11010111",5413 => "01101001",5414 => "00000011",5415 => "11101100",5416 => "01110000",5417 => "01110110",5418 => "01010000",5419 => "11000111",5420 => "00011010",5421 => "01111110",5422 => "00011000",5423 => "01010100",5424 => "10100110",5425 => "11101011",5426 => "00011001",5427 => "00111111",5428 => "01101100",5429 => "10000101",5430 => "00000011",5431 => "11100101",5432 => "10011000",5433 => "10100010",5434 => "10001111",5435 => "10001110",5436 => "00100101",5437 => "00010100",5438 => "11011110",5439 => "01011101",5440 => "11100111",5441 => "10000010",5442 => "11110101",5443 => "00110011",5444 => "11111110",5445 => "10101101",5446 => "00101000",5447 => "10010100",5448 => "00100011",5449 => "11110111",5450 => "11101101",5451 => "10101000",5452 => "00000011",5453 => "11100001",5454 => "10010010",5455 => "01110001",5456 => "11010010",5457 => "11010101",5458 => "10001001",5459 => "10001101",5460 => "01001100",5461 => "00110101",5462 => "10000110",5463 => "10111111",5464 => "01000111",5465 => "01110101",5466 => "00111110",5467 => "10110101",5468 => "01101010",5469 => "01110010",5470 => "11110001",5471 => "11001011",5472 => "11111001",5473 => "00001000",5474 => "10101110",5475 => "01111010",5476 => "10101101",5477 => "01110110",5478 => "10001111",5479 => "00010100",5480 => "01100111",5481 => "01010010",5482 => "10111000",5483 => "00001101",5484 => "11101110",5485 => "01111010",5486 => "00101001",5487 => "10111110",5488 => "00010101",5489 => "01110000",5490 => "11001101",5491 => "01000111",5492 => "01101011",5493 => "11010000",5494 => "10101110",5495 => "01100010",5496 => "01101111",5497 => "01011111",5498 => "00010011",5499 => "00110100",5500 => "11111111",5501 => "00011000",5502 => "01101011",5503 => "00010011",5504 => "11110111",5505 => "11101011",5506 => "10111000",5507 => "11010011",5508 => "00011011",5509 => "00111000",5510 => "10001100",5511 => "01110101",5512 => "00010111",5513 => "00101000",5514 => "11011011",5515 => "01101000",5516 => "01010010",5517 => "01011101",5518 => "01001000",5519 => "10110000",5520 => "01101011",5521 => "11010011",5522 => "11110000",5523 => "00011101",5524 => "10100001",5525 => "11101101",5526 => "00111001",5527 => "01010010",5528 => "11010011",5529 => "10100010",5530 => "11111000",5531 => "10000101",5532 => "01100000",5533 => "01111001",5534 => "11001111",5535 => "10111010",5536 => "10011010",5537 => "11111000",5538 => "01111101",5539 => "01111100",5540 => "01010011",5541 => "11000101",5542 => "10011000",5543 => "11111000",5544 => "00000010",5545 => "10111101",5546 => "01110010",5547 => "00101110",5548 => "01111101",5549 => "00000010",5550 => "00000010",5551 => "11010101",5552 => "01000110",5553 => "00000101",5554 => "11000110",5555 => "10011010",5556 => "10001100",5557 => "11110001",5558 => "11000010",5559 => "00110100",5560 => "10110011",5561 => "00000111",5562 => "00010100",5563 => "11110100",5564 => "11011010",5565 => "11010010",5566 => "01010111",5567 => "10000011",5568 => "11111011",5569 => "01001110",5570 => "01110000",5571 => "10001110",5572 => "10001011",5573 => "10011000",5574 => "10110001",5575 => "00100001",5576 => "10110000",5577 => "11100101",5578 => "11100011",5579 => "01010111",5580 => "01100011",5581 => "10110101",5582 => "11011101",5583 => "01110001",5584 => "10011010",5585 => "11101100",5586 => "10101010",5587 => "01001100",5588 => "00011001",5589 => "10101000",5590 => "00001111",5591 => "01110001",5592 => "11100101",5593 => "10011011",5594 => "10001011",5595 => "11001001",5596 => "00010110",5597 => "00010100",5598 => "11101110",5599 => "00110011",5600 => "00000100",5601 => "01110001",5602 => "10000100",5603 => "10010011",5604 => "01100000",5605 => "00100010",5606 => "11010110",5607 => "00011111",5608 => "10010010",5609 => "00000001",5610 => "11111101",5611 => "00001010",5612 => "10000000",5613 => "10010011",5614 => "11101111",5615 => "01111010",5616 => "00111101",5617 => "10010110",5618 => "11010110",5619 => "01111110",5620 => "10100001",5621 => "10101101",5622 => "11010110",5623 => "11101111",5624 => "11101011",5625 => "01001100",5626 => "11010011",5627 => "11111001",5628 => "01011100",5629 => "01000110",5630 => "10110011",5631 => "11111111",5632 => "10001100",5633 => "01001101",5634 => "11010100",5635 => "01111000",5636 => "11010111",5637 => "11110011",5638 => "10110101",5639 => "11111011",5640 => "00000100",5641 => "00001101",5642 => "10010010",5643 => "11010111",5644 => "01100010",5645 => "10101101",5646 => "01111110",5647 => "10011101",5648 => "11110011",5649 => "10011111",5650 => "10000010",5651 => "11011100",5652 => "11110000",5653 => "00001000",5654 => "11011100",5655 => "11101111",5656 => "00011101",5657 => "10010111",5658 => "10001010",5659 => "10100111",5660 => "01111101",5661 => "10110111",5662 => "10111000",5663 => "00010110",5664 => "10101010",5665 => "11011011",5666 => "01100010",5667 => "11111000",5668 => "01000100",5669 => "01101101",5670 => "01010011",5671 => "11001000",5672 => "01110000",5673 => "10100101",5674 => "10011000",5675 => "11100101",5676 => "00001011",5677 => "11100101",5678 => "00111110",5679 => "00101001",5680 => "10111101",5681 => "01010000",5682 => "10101010",5683 => "10010011",5684 => "01000100",5685 => "10111010",5686 => "10110111",5687 => "01101001",5688 => "01100111",5689 => "11010111",5690 => "11100001",5691 => "01011101",5692 => "00110110",5693 => "01110111",5694 => "10100101",5695 => "01000000",5696 => "00000101",5697 => "01111101",5698 => "10100001",5699 => "10101110",5700 => "10101111",5701 => "10111101",5702 => "01100000",5703 => "11011000",5704 => "00000011",5705 => "01110001",5706 => "10110111",5707 => "11110110",5708 => "00010000",5709 => "00100001",5710 => "11101111",5711 => "01111011",5712 => "10101100",5713 => "10101000",5714 => "10100000",5715 => "11100110",5716 => "11100101",5717 => "00001001",5718 => "11101011",5719 => "10010100",5720 => "11011110",5721 => "11001101",5722 => "10110010",5723 => "01011001",5724 => "01110100",5725 => "01111000",5726 => "10011011",5727 => "00111101",5728 => "10011010",5729 => "00001110",5730 => "00111001",5731 => "00011001",5732 => "11111001",5733 => "10111111",5734 => "00100111",5735 => "10100101",5736 => "00100000",5737 => "10100010",5738 => "10110101",5739 => "00100100",5740 => "10100100",5741 => "01110010",5742 => "10101000",5743 => "00100010",5744 => "11001001",5745 => "11010101",5746 => "11111111",5747 => "00100000",5748 => "11001111",5749 => "01100101",5750 => "01101001",5751 => "11010100",5752 => "11010111",5753 => "00101110",5754 => "01110001",5755 => "00010110",5756 => "00110101",5757 => "10000000",5758 => "00010000",5759 => "10001111",5760 => "11001010",5761 => "00011010",5762 => "11001011",5763 => "00001101",5764 => "01011110",5765 => "00001001",5766 => "01000101",5767 => "10100000",5768 => "11101100",5769 => "10101001",5770 => "01100001",5771 => "00110001",5772 => "00111110",5773 => "10000010",5774 => "01001010",5775 => "00000011",5776 => "10101001",5777 => "01110101",5778 => "01010111",5779 => "00110010",5780 => "00111110",5781 => "01010011",5782 => "11001110",5783 => "01001111",5784 => "00010001",5785 => "11001001",5786 => "11000001",5787 => "11000101",5788 => "11010110",5789 => "11100011",5790 => "10000011",5791 => "00001111",5792 => "00100111",5793 => "11111100",5794 => "11000100",5795 => "11100000",5796 => "10101110",5797 => "11010100",5798 => "00100000",5799 => "01100101",5800 => "10110111",5801 => "01111110",5802 => "10110101",5803 => "01011100",5804 => "11010001",5805 => "11110010",5806 => "00111001",5807 => "00010000",5808 => "01111101",5809 => "01110110",5810 => "10000000",5811 => "00000001",5812 => "11110111",5813 => "10010111",5814 => "10101010",5815 => "11110001",5816 => "11011011",5817 => "11000011",5818 => "10110000",5819 => "00100101",5820 => "11001001",5821 => "01001001",5822 => "10001110",5823 => "00010101",5824 => "00000000",5825 => "01110110",5826 => "10001001",5827 => "10000100",5828 => "11001111",5829 => "11100000",5830 => "10001101",5831 => "01100011",5832 => "10100010",5833 => "00100010",5834 => "01000011",5835 => "10000111",5836 => "11010101",5837 => "01110101",5838 => "10001011",5839 => "01010001",5840 => "01100111",5841 => "11111001",5842 => "10000011",5843 => "01100101",5844 => "01001000",5845 => "00110110",5846 => "00110111",5847 => "10110011",5848 => "01100111",5849 => "01111011",5850 => "11000011",5851 => "01111110",5852 => "11011101",5853 => "11111101",5854 => "11111001",5855 => "10110110",5856 => "10111011",5857 => "10110001",5858 => "10010010",5859 => "11001000",5860 => "01100000",5861 => "10010001",5862 => "10100101",5863 => "10111111",5864 => "10110011",5865 => "01010101",5866 => "11001101",5867 => "11000001",5868 => "10011100",5869 => "11101100",5870 => "01100111",5871 => "00111111",5872 => "01110001",5873 => "01001011",5874 => "00001010",5875 => "10110001",5876 => "00010010",5877 => "01011111",5878 => "00011001",5879 => "10000010",5880 => "00001011",5881 => "10101101",5882 => "01011010",5883 => "01001110",5884 => "10011000",5885 => "10011101",5886 => "11101001",5887 => "01010010",5888 => "11010010",5889 => "00011111",5890 => "01111000",5891 => "11101000",5892 => "00101011",5893 => "10000011",5894 => "11010101",5895 => "01100111",5896 => "10101100",5897 => "01100110",5898 => "00101100",5899 => "10010000",5900 => "10010010",5901 => "00111001",5902 => "01111010",5903 => "11110001",5904 => "11010011",5905 => "10010010",5906 => "01010011",5907 => "01000000",5908 => "11001111",5909 => "00010101",5910 => "10110111",5911 => "00011000",5912 => "10101101",5913 => "00011100",5914 => "11001000",5915 => "10111000",5916 => "11110010",5917 => "01110001",5918 => "11101011",5919 => "11111001",5920 => "10000110",5921 => "01000101",5922 => "11011011",5923 => "01011001",5924 => "01010001",5925 => "10110110",5926 => "01111000",5927 => "00111000",5928 => "11101011",5929 => "10110010",5930 => "10110110",5931 => "11001110",5932 => "10000101",5933 => "01100100",5934 => "01111101",5935 => "11000000",5936 => "01000000",5937 => "11001010",5938 => "00111001",5939 => "01110110",5940 => "01010001",5941 => "00100011",5942 => "01000001",5943 => "01010111",5944 => "00100110",5945 => "01100010",5946 => "00111011",5947 => "10101110",5948 => "00100011",5949 => "00010001",5950 => "11100011",5951 => "10011010",5952 => "10010011",5953 => "01000010",5954 => "11110011",5955 => "01000001",5956 => "11111100",5957 => "11011110",5958 => "10110011",5959 => "01011100",5960 => "11001110",5961 => "00110100",5962 => "00000111",5963 => "01110000",5964 => "11100010",5965 => "01000110",5966 => "11101111",5967 => "01010001",5968 => "00110110",5969 => "00100101",5970 => "01101110",5971 => "00100111",5972 => "00111001",5973 => "10011000",5974 => "10000100",5975 => "10010010",5976 => "11101011",5977 => "11100100",5978 => "00100000",5979 => "01110101",5980 => "01011111",5981 => "01000001",5982 => "00111010",5983 => "00011101",5984 => "10010011",5985 => "11100000",5986 => "11110000",5987 => "10000000",5988 => "00100101",5989 => "00100111",5990 => "10110100",5991 => "11100100",5992 => "11111101",5993 => "00010000",5994 => "11110110",5995 => "01101100",5996 => "01111101",5997 => "01000011",5998 => "00101111",5999 => "01011110",6000 => "00010101",6001 => "11111100",6002 => "00110000",6003 => "10101001",6004 => "00101101",6005 => "01011110",6006 => "00011011",6007 => "00110110",6008 => "00110100",6009 => "00000110",6010 => "10110010",6011 => "10010001",6012 => "01111001",6013 => "11110000",6014 => "10000000",6015 => "10011110",6016 => "01011111",6017 => "11001111",6018 => "01000010",6019 => "00010001",6020 => "01011001",6021 => "01100011",6022 => "11000110",6023 => "10011000",6024 => "10001011",6025 => "11001100",6026 => "11010101",6027 => "00110100",6028 => "11101111",6029 => "11100010",6030 => "00101000",6031 => "10111011",6032 => "11001100",6033 => "01010100",6034 => "00001110",6035 => "11010011",6036 => "11101001",6037 => "00000010",6038 => "10011011",6039 => "11011001",6040 => "01100111",6041 => "10000111",6042 => "01001011",6043 => "10101011",6044 => "11000100",6045 => "10011001",6046 => "11010001",6047 => "11010100",6048 => "00111101",6049 => "11001101",6050 => "10011001",6051 => "01100001",6052 => "10000111",6053 => "10110111",6054 => "10110001",6055 => "10011100",6056 => "01000111",6057 => "01010111",6058 => "00001000",6059 => "01010000",6060 => "10110011",6061 => "11111010",6062 => "01101100",6063 => "10100100",6064 => "00011100",6065 => "00001011",6066 => "11100110",6067 => "11011111",6068 => "10111000",6069 => "10010001",6070 => "11000011",6071 => "00000101",6072 => "00100110",6073 => "10000011",6074 => "10001001",6075 => "01111111",6076 => "11101101",6077 => "10111011",6078 => "01011010",6079 => "10000101",6080 => "11110000",6081 => "00110010",6082 => "01101010",6083 => "10010000",6084 => "11101010",6085 => "10011100",6086 => "11111000",6087 => "10001110",6088 => "10110000",6089 => "11110101",6090 => "10100100",6091 => "01101100",6092 => "11001001",6093 => "01001111",6094 => "11000011",6095 => "00100010",6096 => "10110000",6097 => "10010101",6098 => "11011100",6099 => "00110000",6100 => "10111011",6101 => "00010000",6102 => "11010100",6103 => "01110001",6104 => "01110010",6105 => "10111011",6106 => "11100010",6107 => "00101001",6108 => "00000001",6109 => "10110011",6110 => "10100000",6111 => "10010000",6112 => "00000000",6113 => "10011000",6114 => "00011110",6115 => "01011111",6116 => "00010001",6117 => "00000110",6118 => "10110000",6119 => "01111000",6120 => "01111011",6121 => "10101111",6122 => "10101111",6123 => "00010001",6124 => "10010111",6125 => "10101010",6126 => "10001001",6127 => "10101011",6128 => "10001111",6129 => "11101100",6130 => "11101010",6131 => "01101010",6132 => "11111000",6133 => "00111000",6134 => "00010110",6135 => "00110010",6136 => "00110011",6137 => "11000010",6138 => "10111100",6139 => "01000000",6140 => "01001110",6141 => "01011110",6142 => "10001010",6143 => "00111000",6144 => "11110110",6145 => "00010010",6146 => "00100001",6147 => "00001010",6148 => "11110000",6149 => "11100110",6150 => "01100111",6151 => "10000000",6152 => "11101101",6153 => "00111111",6154 => "11010110",6155 => "11101111",6156 => "10100010",6157 => "00001101",6158 => "01000111",6159 => "01111101",6160 => "00100101",6161 => "01111110",6162 => "10010000",6163 => "10010000",6164 => "10101110",6165 => "11101101",6166 => "00011101",6167 => "10000001",6168 => "01011000",6169 => "01001111",6170 => "11000110",6171 => "11011101",6172 => "11110101",6173 => "01000000",6174 => "10101101",6175 => "00011101",6176 => "00101001",6177 => "00001001",6178 => "10001010",6179 => "00011000",6180 => "01110001",6181 => "11010100",6182 => "11101111",6183 => "00111101",6184 => "11110101",6185 => "00110111",6186 => "00010100",6187 => "01010001",6188 => "01011100",6189 => "11001111",6190 => "10001011",6191 => "10100011",6192 => "01000111",6193 => "11111101",6194 => "11111110",6195 => "01011000",6196 => "10111111",6197 => "00001111",6198 => "00101001",6199 => "00110101",6200 => "10010001",6201 => "10001000",6202 => "10110010",6203 => "11101100",6204 => "10000110",6205 => "11010101",6206 => "00110001",6207 => "01010011",6208 => "10010101",6209 => "10001000",6210 => "11101011",6211 => "01111010",6212 => "01111011",6213 => "10001101",6214 => "11101101",6215 => "11011110",6216 => "00001011",6217 => "00001101",6218 => "00001100",6219 => "01001111",6220 => "01111111",6221 => "01010100",6222 => "01101101",6223 => "00011011",6224 => "11111000",6225 => "01000011",6226 => "11001110",6227 => "01110100",6228 => "00010101",6229 => "11111111",6230 => "01110100",6231 => "01001010",6232 => "00100100",6233 => "10001110",6234 => "10001101",6235 => "01001010",6236 => "01000110",6237 => "01001001",6238 => "01011001",6239 => "01110101",6240 => "11100001",6241 => "11110111",6242 => "11111111",6243 => "10110110",6244 => "10100100",6245 => "00010111",6246 => "11010001",6247 => "11011011",6248 => "11111111",6249 => "00111111",6250 => "10001010",6251 => "00000100",6252 => "10000111",6253 => "01100011",6254 => "01110000",6255 => "01001010",6256 => "01010011",6257 => "00000100",6258 => "00101100",6259 => "10010011",6260 => "11010000",6261 => "11000000",6262 => "00100011",6263 => "00111101",6264 => "01100001",6265 => "00101100",6266 => "01110011",6267 => "10110000",6268 => "01110100",6269 => "01100001",6270 => "10111101",6271 => "00011110",6272 => "10011001",6273 => "10010000",6274 => "00000101",6275 => "00001010",6276 => "01100100",6277 => "10100110",6278 => "10111101",6279 => "10011101",6280 => "00010001",6281 => "10011111",6282 => "11111100",6283 => "01001010",6284 => "01001101",6285 => "00010101",6286 => "01000010",6287 => "11110001",6288 => "01010010",6289 => "10010010",6290 => "11111111",6291 => "10010000",6292 => "10101111",6293 => "10001100",6294 => "11001011",6295 => "10001110",6296 => "11100010",6297 => "11001011",6298 => "00101010",6299 => "10100000",6300 => "00100010",6301 => "01010001",6302 => "10100000",6303 => "11010010",6304 => "10010010",6305 => "10111011",6306 => "11100100",6307 => "01010010",6308 => "10011001",6309 => "01011001",6310 => "00011000",6311 => "00010110",6312 => "10100110",6313 => "01110100",6314 => "10111101",6315 => "11011011",6316 => "00100000",6317 => "10110010",6318 => "10001010",6319 => "00000010",6320 => "10100100",6321 => "01110011",6322 => "01101111",6323 => "11000110",6324 => "00010001",6325 => "01111011",6326 => "11101010",6327 => "11010101",6328 => "11001111",6329 => "01101100",6330 => "11000100",6331 => "00010101",6332 => "10010110",6333 => "01010000",6334 => "00010101",6335 => "11100110",6336 => "00010000",6337 => "00110000",6338 => "01110010",6339 => "00010001",6340 => "11111011",6341 => "00111001",6342 => "01011110",6343 => "01101010",6344 => "10011100",6345 => "00010001",6346 => "01011110",6347 => "10001010",6348 => "10110111",6349 => "01100100",6350 => "01100111",6351 => "11010110",6352 => "01100101",6353 => "10101100",6354 => "11011110",6355 => "11101001",6356 => "00110100",6357 => "01011010",6358 => "00100001",6359 => "11100100",6360 => "01011101",6361 => "00101001",6362 => "10001110",6363 => "11011000",6364 => "10011001",6365 => "00010110",6366 => "01110110",6367 => "11110001",6368 => "01011010",6369 => "01101100",6370 => "01000001",6371 => "01101001",6372 => "00000000",6373 => "10100100",6374 => "10001010",6375 => "00110000",6376 => "01100011",6377 => "00111000",6378 => "01101010",6379 => "01001111",6380 => "01100010",6381 => "00001001",6382 => "01100111",6383 => "01101111",6384 => "11110011",6385 => "00001001",6386 => "10111001",6387 => "01100110",6388 => "01001110",6389 => "11011110",6390 => "01101001",6391 => "00001010",6392 => "10011111",6393 => "01010110",6394 => "01010100",6395 => "00000101",6396 => "10000101",6397 => "01011010",6398 => "01001111",6399 => "11001110",6400 => "11011101",6401 => "01000001",6402 => "01011110",6403 => "00100110",6404 => "01010010",6405 => "11101100",6406 => "01000110",6407 => "01001000",6408 => "01100010",6409 => "10110011",6410 => "10001110",6411 => "11011010",6412 => "01010110",6413 => "01001011",6414 => "01000010",6415 => "01101010",6416 => "01001010",6417 => "10000011",6418 => "10111110",6419 => "00100001",6420 => "00110110",6421 => "00101101",6422 => "00101101",6423 => "01010111",6424 => "11110101",6425 => "01111110",6426 => "00011101",6427 => "11000011",6428 => "10011101",6429 => "11100110",6430 => "00110110",6431 => "00010000",6432 => "01100101",6433 => "10100101",6434 => "11111101",6435 => "10100001",6436 => "10001000",6437 => "11011000",6438 => "11101010",6439 => "11101110",6440 => "10011101",6441 => "10111111",6442 => "11110111",6443 => "11001101",6444 => "00101001",6445 => "10110101",6446 => "10011101",6447 => "01011101",6448 => "00000111",6449 => "01111100",6450 => "01101001",6451 => "01110001",6452 => "01000110",6453 => "11111011",6454 => "01110101",6455 => "10001011",6456 => "00011011",6457 => "00100011",6458 => "11111110",6459 => "10011110",6460 => "10110100",6461 => "00001111",6462 => "00000011",6463 => "10010010",6464 => "11011110",6465 => "00001101",6466 => "10111101",6467 => "11001110",6468 => "00110110",6469 => "11011010",6470 => "10000011",6471 => "10100011",6472 => "11100000",6473 => "10100110",6474 => "00111010",6475 => "01100000",6476 => "10101000",6477 => "10011111",6478 => "01001101",6479 => "00110100",6480 => "00100011",6481 => "11000111",6482 => "01110111",6483 => "00110101",6484 => "01010000",6485 => "01000100",6486 => "01001110",6487 => "11100101",6488 => "10000100",6489 => "10110010",6490 => "01011011",6491 => "00111100",6492 => "11100010",6493 => "10011111",6494 => "00110100",6495 => "01010011",6496 => "00111001",6497 => "11110111",6498 => "01111110",6499 => "01111001",6500 => "10011011",6501 => "00001110",6502 => "01010100",6503 => "11101111",6504 => "01000000",6505 => "10001000",6506 => "11001101",6507 => "10101000",6508 => "10010000",6509 => "01010000",6510 => "01111001",6511 => "10111000",6512 => "10100101",6513 => "00011010",6514 => "11010010",6515 => "10101010",6516 => "01010101",6517 => "01010111",6518 => "11001010",6519 => "01111001",6520 => "01110000",6521 => "01010011",6522 => "10101110",6523 => "01110110",6524 => "11001010",6525 => "01100010",6526 => "11100001",6527 => "00010001",6528 => "11001110",6529 => "01110010",6530 => "10111111",6531 => "00110100",6532 => "01000100",6533 => "00001110",6534 => "01101101",6535 => "11110100",6536 => "01011100",6537 => "10111101",6538 => "00111100",6539 => "10101110",6540 => "00101010",6541 => "11000100",6542 => "01001001",6543 => "11111001",6544 => "00111110",6545 => "10010101",6546 => "10010000",6547 => "10100001",6548 => "01111111",6549 => "10001010",6550 => "00011011",6551 => "01101000",6552 => "01111011",6553 => "11001111",6554 => "00111001",6555 => "00001001",6556 => "00010100",6557 => "00110011",6558 => "01010101",6559 => "01110001",6560 => "10111011",6561 => "01101000",6562 => "11000100",6563 => "11100100",6564 => "01010111",6565 => "00001000",6566 => "01010001",6567 => "10101111",6568 => "00011110",6569 => "00111111",6570 => "10010001",6571 => "00101111",6572 => "11011001",6573 => "11011100",6574 => "10001011",6575 => "01101001",6576 => "01001011",6577 => "01001011",6578 => "11000110",6579 => "11000011",6580 => "01001010",6581 => "00110110",6582 => "10111000",6583 => "00111011",6584 => "11110111",6585 => "01100110",6586 => "01010010",6587 => "00111101",6588 => "10011101",6589 => "00010011",6590 => "11000000",6591 => "10000011",6592 => "10010001",6593 => "10100011",6594 => "01011110",6595 => "01000110",6596 => "10000001",6597 => "00011001",6598 => "11101111",6599 => "10111010",6600 => "01101100",6601 => "10101100",6602 => "00101011",6603 => "10111010",6604 => "11011111",6605 => "01100011",6606 => "10010011",6607 => "10000001",6608 => "00101001",6609 => "01101100",6610 => "01010001",6611 => "11001101",6612 => "00111000",6613 => "01001011",6614 => "00100001",6615 => "00000000",6616 => "11100000",6617 => "10111110",6618 => "00100101",6619 => "10010111",6620 => "00011010",6621 => "10100010",6622 => "10110111",6623 => "10010101",6624 => "00110010",6625 => "00110111",6626 => "01111100",6627 => "01010110",6628 => "00111000",6629 => "10001011",6630 => "10001110",6631 => "01000110",6632 => "01000010",6633 => "11110100",6634 => "10010000",6635 => "01001110",6636 => "10000111",6637 => "00100011",6638 => "10001100",6639 => "01111010",6640 => "01010011",6641 => "01011011",6642 => "01011010",6643 => "01001000",6644 => "00100000",6645 => "11001011",6646 => "11100111",6647 => "11100011",6648 => "11011110",6649 => "00110001",6650 => "11011111",6651 => "11101000",6652 => "10000011",6653 => "11001100",6654 => "11101000",6655 => "00011010",6656 => "10010110",6657 => "10000100",6658 => "10110010",6659 => "01011001",6660 => "11011110",6661 => "00010001",6662 => "01010110",6663 => "11011111",6664 => "11011001",6665 => "01010110",6666 => "00101111",6667 => "11010000",6668 => "01111001",6669 => "00001000",6670 => "00100111",6671 => "11101110",6672 => "01101101",6673 => "01001111",6674 => "11100101",6675 => "10010111",6676 => "01011110",6677 => "00011011",6678 => "00101010",6679 => "11001100",6680 => "10011100",6681 => "10110011",6682 => "10001011",6683 => "01001000",6684 => "01010111",6685 => "00001010",6686 => "00011010",6687 => "10100110",6688 => "10100000",6689 => "10101000",6690 => "10011110",6691 => "10011111",6692 => "11100001",6693 => "10101000",6694 => "00110110",6695 => "00100111",6696 => "10001001",6697 => "10001101",6698 => "01010110",6699 => "01101100",6700 => "00001000",6701 => "11100101",6702 => "00001001",6703 => "00110111",6704 => "11011111",6705 => "01101001",6706 => "01110000",6707 => "00110010",6708 => "00111001",6709 => "00010110",6710 => "00100011",6711 => "10110100",6712 => "10000110",6713 => "11100100",6714 => "01110000",6715 => "11111010",6716 => "00110100",6717 => "00011001",6718 => "11010101",6719 => "10010011",6720 => "01001011",6721 => "10000110",6722 => "10010001",6723 => "01101001",6724 => "01000110",6725 => "10000011",6726 => "00001110",6727 => "01010010",6728 => "11001110",6729 => "10010011",6730 => "01000111",6731 => "11001000",6732 => "11010110",6733 => "01011110",6734 => "11110101",6735 => "10011000",6736 => "00010111",6737 => "11101001",6738 => "11111011",6739 => "11100000",6740 => "10011011",6741 => "00000001",6742 => "01001011",6743 => "10010011",6744 => "00010100",6745 => "11000011",6746 => "00100001",6747 => "01101000",6748 => "00101000",6749 => "11110110",6750 => "00111010",6751 => "01010110",6752 => "01101001",6753 => "10011100",6754 => "01111011",6755 => "10000000",6756 => "11101101",6757 => "00110010",6758 => "10101010",6759 => "01011001",6760 => "11011111",6761 => "01010101",6762 => "00001111",6763 => "00111111",6764 => "11000010",6765 => "10000101",6766 => "10111111",6767 => "01110111",6768 => "11010111",6769 => "01010110",6770 => "01101101",6771 => "00000110",6772 => "00111010",6773 => "00010001",6774 => "00011000",6775 => "00010101",6776 => "11001001",6777 => "10011000",6778 => "11101110",6779 => "11010101",6780 => "00100001",6781 => "00100010",6782 => "00001011",6783 => "01110011",6784 => "10111010",6785 => "11101100",6786 => "10011010",6787 => "10110011",6788 => "10111011",6789 => "11100011",6790 => "01101000",6791 => "01111100",6792 => "10000011",6793 => "01001000",6794 => "00011111",6795 => "10010001",6796 => "10111011",6797 => "00101000",6798 => "11110100",6799 => "10010101",6800 => "01000110",6801 => "01110101",6802 => "11000110",6803 => "10100110",6804 => "10000010",6805 => "10011000",6806 => "00010100",6807 => "00010110",6808 => "01010000",6809 => "00011101",6810 => "11001100",6811 => "10011110",6812 => "11010101",6813 => "10001010",6814 => "00010111",6815 => "00010011",6816 => "11000100",6817 => "01011110",6818 => "10001011",6819 => "11100111",6820 => "10001101",6821 => "00001000",6822 => "10010001",6823 => "10000000",6824 => "00100010",6825 => "11011100",6826 => "11111010",6827 => "01001011",6828 => "11100010",6829 => "10011101",6830 => "10001001",6831 => "01110101",6832 => "01101101",6833 => "01111010",6834 => "01010001",6835 => "01100010",6836 => "11001100",6837 => "00100101",6838 => "00010011",6839 => "11110110",6840 => "10110001",6841 => "11000011",6842 => "10101011",6843 => "10111010",6844 => "10010000",6845 => "01001011",6846 => "00010111",6847 => "01110011",6848 => "00100001",6849 => "01111111",6850 => "10001101",6851 => "11101001",6852 => "11001110",6853 => "00101101",6854 => "01100111",6855 => "01010001",6856 => "11000110",6857 => "00101011",6858 => "00000101",6859 => "11111101",6860 => "10110101",6861 => "00010000",6862 => "01110001",6863 => "00101010",6864 => "00110101",6865 => "11010011",6866 => "10100011",6867 => "11011100",6868 => "10001011",6869 => "11110111",6870 => "00000010",6871 => "10100101",6872 => "10011000",6873 => "10101101",6874 => "00010101",6875 => "01110010",6876 => "01100111",6877 => "01011111",6878 => "00010000",6879 => "01111101",6880 => "11110011",6881 => "01110001",6882 => "11101100",6883 => "11010110",6884 => "00101000",6885 => "10101101",6886 => "01110101",6887 => "11011011",6888 => "00101000",6889 => "11000011",6890 => "00010110",6891 => "01000001",6892 => "11001101",6893 => "11111010",6894 => "01111010",6895 => "00110110",6896 => "01110001",6897 => "01010111",6898 => "01001101",6899 => "01110100",6900 => "10000101",6901 => "11001100",6902 => "00100100",6903 => "00001010",6904 => "00011111",6905 => "11001011",6906 => "11110110",6907 => "00001010",6908 => "10001001",6909 => "11101011",6910 => "00110101",6911 => "00000001",6912 => "11011100",6913 => "10111010",6914 => "00110111",6915 => "11101011",6916 => "01001100",6917 => "10100101",6918 => "11001101",6919 => "10110101",6920 => "11100100",6921 => "11111100",6922 => "10110100",6923 => "10111110",6924 => "10101000",6925 => "10011101",6926 => "10110010",6927 => "00100101",6928 => "00110100",6929 => "01101011",6930 => "10110001",6931 => "01100001",6932 => "00111110",6933 => "01010001",6934 => "10010000",6935 => "11100000",6936 => "11111100",6937 => "10011010",6938 => "10010101",6939 => "01001111",6940 => "11110011",6941 => "01010100",6942 => "01010001",6943 => "00000011",6944 => "10001111",6945 => "11011001",6946 => "11111001",6947 => "10101010",6948 => "00111000",6949 => "10111010",6950 => "11110111",6951 => "11001100",6952 => "10101100",6953 => "11010111",6954 => "01111110",6955 => "11100010",6956 => "11000001",6957 => "10101011",6958 => "10110000",6959 => "11001010",6960 => "10011100",6961 => "01000101",6962 => "00010000",6963 => "10000101",6964 => "01001001",6965 => "11001101",6966 => "00101101",6967 => "01110010",6968 => "11111011",6969 => "10011000",6970 => "00000011",6971 => "10001110",6972 => "10011101",6973 => "10001001",6974 => "11100100",6975 => "11000100",6976 => "11000011",6977 => "10001001",6978 => "10001000",6979 => "00010000",6980 => "10100111",6981 => "11010100",6982 => "10010001",6983 => "00000111",6984 => "01100110",6985 => "10101110",6986 => "00110001",6987 => "01001011",6988 => "01101111",6989 => "01001111",6990 => "01001100",6991 => "11100010",6992 => "00101111",6993 => "00011101",6994 => "10110011",6995 => "11100111",6996 => "01101011",6997 => "00001010",6998 => "11101001",6999 => "10100100",7000 => "11110011",7001 => "01100000",7002 => "10110000",7003 => "10001101",7004 => "00001010",7005 => "11101110",7006 => "01100000",7007 => "01110011",7008 => "00010110",7009 => "01001010",7010 => "10100101",7011 => "01001100",7012 => "11011111",7013 => "10000000",7014 => "11011111",7015 => "00001101",7016 => "00101110",7017 => "10001011",7018 => "10110001",7019 => "11111000",7020 => "00000001",7021 => "00101001",7022 => "11101000",7023 => "00011010",7024 => "01011111",7025 => "11101000",7026 => "00111101",7027 => "00010111",7028 => "00100110",7029 => "11110000",7030 => "00111010",7031 => "00011100",7032 => "01010010",7033 => "01001110",7034 => "00010101",7035 => "01100100",7036 => "01000010",7037 => "01101110",7038 => "01100000",7039 => "10101110",7040 => "00001011",7041 => "10101110",7042 => "10010001",7043 => "00100010",7044 => "01110101",7045 => "11011101",7046 => "10111100",7047 => "00010111",7048 => "10111100",7049 => "00110110",7050 => "01111011",7051 => "00100000",7052 => "01111100",7053 => "01111101",7054 => "01010111",7055 => "00110001",7056 => "11101110",7057 => "11000101",7058 => "10001100",7059 => "00001011",7060 => "00101111",7061 => "11000100",7062 => "00111011",7063 => "01100011",7064 => "11110011",7065 => "01101100",7066 => "11111011",7067 => "01110110",7068 => "01110001",7069 => "01101111",7070 => "10011001",7071 => "01101000",7072 => "01001110",7073 => "10000111",7074 => "11101010",7075 => "01000111",7076 => "00110010",7077 => "11010100",7078 => "01100100",7079 => "00101001",7080 => "11111101",7081 => "11101101",7082 => "01101011",7083 => "10001101",7084 => "10110001",7085 => "00001011",7086 => "10110101",7087 => "01101000",7088 => "00001111",7089 => "11110110",7090 => "10111100",7091 => "01111111",7092 => "00001000",7093 => "00110011",7094 => "11110111",7095 => "10000101",7096 => "11001111",7097 => "01111011",7098 => "00110011",7099 => "00000100",7100 => "00111011",7101 => "01010101",7102 => "10101111",7103 => "01000000",7104 => "10001001",7105 => "01010000",7106 => "10010011",7107 => "11010001",7108 => "11100110",7109 => "01101011",7110 => "01011010",7111 => "11011010",7112 => "10001111",7113 => "10000100",7114 => "11010001",7115 => "01101111",7116 => "11010101",7117 => "00010101",7118 => "10100101",7119 => "00001001",7120 => "11001111",7121 => "00101010",7122 => "10000011",7123 => "10100001",7124 => "11101001",7125 => "10111010",7126 => "00010111",7127 => "11110111",7128 => "00011000",7129 => "01100010",7130 => "10001010",7131 => "11110000",7132 => "11011010",7133 => "11010111",7134 => "10111010",7135 => "01001101",7136 => "00111011",7137 => "10100111",7138 => "00011010",7139 => "01000000",7140 => "01011110",7141 => "11001100",7142 => "01011011",7143 => "11110010",7144 => "11000010",7145 => "01010111",7146 => "10101001",7147 => "01111111",7148 => "00000111",7149 => "10000100",7150 => "10010110",7151 => "10100100",7152 => "01001111",7153 => "11110110",7154 => "00111010",7155 => "11010010",7156 => "01101101",7157 => "10000101",7158 => "01000111",7159 => "00000000",7160 => "11110101",7161 => "10110001",7162 => "00011011",7163 => "00101011",7164 => "10001001",7165 => "01010110",7166 => "00001001",7167 => "01011110",7168 => "11100000",7169 => "00000001",7170 => "00110110",7171 => "10010011",7172 => "00110101",7173 => "00011000",7174 => "00101101",7175 => "01000001",7176 => "00111110",7177 => "10010101",7178 => "01011000",7179 => "10110001",7180 => "11100011",7181 => "10100101",7182 => "00100001",7183 => "10111101",7184 => "01001001",7185 => "01000010",7186 => "01001110",7187 => "10110001",7188 => "00011001",7189 => "11111011",7190 => "11100010",7191 => "11101010",7192 => "11101110",7193 => "00100100",7194 => "10000010",7195 => "01100110",7196 => "00110010",7197 => "00111010",7198 => "00010100",7199 => "01001100",7200 => "00110111",7201 => "00001001",7202 => "10001000",7203 => "01001110",7204 => "10100011",7205 => "00000101",7206 => "00000101",7207 => "00000001",7208 => "11010100",7209 => "11111110",7210 => "00010000",7211 => "00110001",7212 => "01101011",7213 => "11011000",7214 => "01111000",7215 => "11001010",7216 => "10110100",7217 => "11011100",7218 => "10111111",7219 => "01100111",7220 => "10010111",7221 => "11110100",7222 => "10000100",7223 => "11001110",7224 => "00010111",7225 => "01111011",7226 => "11111000",7227 => "01011100",7228 => "00110010",7229 => "11000010",7230 => "11100001",7231 => "01110010",7232 => "10011100",7233 => "11110000",7234 => "01011111",7235 => "01110101",7236 => "01101111",7237 => "00001000",7238 => "11111000",7239 => "10111100",7240 => "10011010",7241 => "00110110",7242 => "10010110",7243 => "00000111",7244 => "01101001",7245 => "11010111",7246 => "01101001",7247 => "11010101",7248 => "01001011",7249 => "00100110",7250 => "11011001",7251 => "00101001",7252 => "10010110",7253 => "00000111",7254 => "10000001",7255 => "00101011",7256 => "00111100",7257 => "10101001",7258 => "11001000",7259 => "10001001",7260 => "10100000",7261 => "10000110",7262 => "01101100",7263 => "10001011",7264 => "11010001",7265 => "11111110",7266 => "01111010",7267 => "01011111",7268 => "01101101",7269 => "11110111",7270 => "10011011",7271 => "11011000",7272 => "00010101",7273 => "11010100",7274 => "00101011",7275 => "00110111",7276 => "00110001",7277 => "11100010",7278 => "10001101",7279 => "11100111",7280 => "10000100",7281 => "10100011",7282 => "11111000",7283 => "11001111",7284 => "00000011",7285 => "11100011",7286 => "01010111",7287 => "10001011",7288 => "10101110",7289 => "00111101",7290 => "11100011",7291 => "11011101",7292 => "11001111",7293 => "01110000",7294 => "11000111",7295 => "01111000",7296 => "00000000",7297 => "10011110",7298 => "01111011",7299 => "00001111",7300 => "10101101",7301 => "11010110",7302 => "00110101",7303 => "01001101",7304 => "10110110",7305 => "10001111",7306 => "10100011",7307 => "01100011",7308 => "01010000",7309 => "00010101",7310 => "11000110",7311 => "11001011",7312 => "01001110",7313 => "01101110",7314 => "10001010",7315 => "00011001",7316 => "11000001",7317 => "01100110",7318 => "11110111",7319 => "10011001",7320 => "10110010",7321 => "11011011",7322 => "01010011",7323 => "11000000",7324 => "00100100",7325 => "00110010",7326 => "01011001",7327 => "01111111",7328 => "00000111",7329 => "00010111",7330 => "11100000",7331 => "01011000",7332 => "01101110",7333 => "00001101",7334 => "01101100",7335 => "11111011",7336 => "11000011",7337 => "10001001",7338 => "00101100",7339 => "11000010",7340 => "11111100",7341 => "10100110",7342 => "10111010",7343 => "11010101",7344 => "11101001",7345 => "01110101",7346 => "11000011",7347 => "01010111",7348 => "00111101",7349 => "10011101",7350 => "01000100",7351 => "01010000",7352 => "10001101",7353 => "11100010",7354 => "11100010",7355 => "01001000",7356 => "11101001",7357 => "10111000",7358 => "01111100",7359 => "01111100",7360 => "11010100",7361 => "01010100",7362 => "00010001",7363 => "00000011",7364 => "00000000",7365 => "10000111",7366 => "01110010",7367 => "01001111",7368 => "01000111",7369 => "11000001",7370 => "10110100",7371 => "10110100",7372 => "10101011",7373 => "10100110",7374 => "11010010",7375 => "01000000",7376 => "01011010",7377 => "00100001",7378 => "01000010",7379 => "01010101",7380 => "00001111",7381 => "10000101",7382 => "11100001",7383 => "11011101",7384 => "11000011",7385 => "11011010",7386 => "01100001",7387 => "01011101",7388 => "10101001",7389 => "11110010",7390 => "11110000",7391 => "01000000",7392 => "01111110",7393 => "00010001",7394 => "11000000",7395 => "01110111",7396 => "01000010",7397 => "10101101",7398 => "11010001",7399 => "11101100",7400 => "01100110",7401 => "11100100",7402 => "01101111",7403 => "11001000",7404 => "10011011",7405 => "01001001",7406 => "00100001",7407 => "00010001",7408 => "11101000",7409 => "10001101",7410 => "01101110",7411 => "11010001",7412 => "10110011",7413 => "11001100",7414 => "00001001",7415 => "01101111",7416 => "00101100",7417 => "00100111",7418 => "00110011",7419 => "01100000",7420 => "00111010",7421 => "00001110",7422 => "00111010",7423 => "10100001",7424 => "00100101",7425 => "11010111",7426 => "00111001",7427 => "01000011",7428 => "00010011",7429 => "01000111",7430 => "01101001",7431 => "11010101",7432 => "00011010",7433 => "01110100",7434 => "00001001",7435 => "11100011",7436 => "11011110",7437 => "00110001",7438 => "01101110",7439 => "10100010",7440 => "10100000",7441 => "01010011",7442 => "11000011",7443 => "10100011",7444 => "00110000",7445 => "01100010",7446 => "11010110",7447 => "01111111",7448 => "11110010",7449 => "10001101",7450 => "01010010",7451 => "11011110",7452 => "00010010",7453 => "10000111",7454 => "00111100",7455 => "00101101",7456 => "00001110",7457 => "10011011",7458 => "11010110",7459 => "00110110",7460 => "11011011",7461 => "10110110",7462 => "10011010",7463 => "01101011",7464 => "11101101",7465 => "01110111",7466 => "00010001",7467 => "01110100",7468 => "00011110",7469 => "00111100",7470 => "10011111",7471 => "00010101",7472 => "00001000",7473 => "11010101",7474 => "00000110",7475 => "01101001",7476 => "11001111",7477 => "01010101",7478 => "01011110",7479 => "01011011",7480 => "01111110",7481 => "10001001",7482 => "01011111",7483 => "11001110",7484 => "11000011",7485 => "01000100",7486 => "00111110",7487 => "11001100",7488 => "10100000",7489 => "01110110",7490 => "10010000",7491 => "00001001",7492 => "00001001",7493 => "00100100",7494 => "10111000",7495 => "10000111",7496 => "10001101",7497 => "01001100",7498 => "01010001",7499 => "11110000",7500 => "10111110",7501 => "00101001",7502 => "10000101",7503 => "11111001",7504 => "10111010",7505 => "00001111",7506 => "00000001",7507 => "01001110",7508 => "11110101",7509 => "00011101",7510 => "10100110",7511 => "10111000",7512 => "11100001",7513 => "10101001",7514 => "10011100",7515 => "10001110",7516 => "10000010",7517 => "11111110",7518 => "00101100",7519 => "00011010",7520 => "01111000",7521 => "01001011",7522 => "10000111",7523 => "01001101",7524 => "11010111",7525 => "10001011",7526 => "01100000",7527 => "01010001",7528 => "11000001",7529 => "11000001",7530 => "10101100",7531 => "01000011",7532 => "10111011",7533 => "11011101",7534 => "01000001",7535 => "01011100",7536 => "11110001",7537 => "01001000",7538 => "10111000",7539 => "10111000",7540 => "10000001",7541 => "11010011",7542 => "01111101",7543 => "10001010",7544 => "10011010",7545 => "11111110",7546 => "11011100",7547 => "01000001",7548 => "00011010",7549 => "01111010",7550 => "01000110",7551 => "01110010",7552 => "10010100",7553 => "01101010",7554 => "00111011",7555 => "11011000",7556 => "00110000",7557 => "11000010",7558 => "01100111",7559 => "00100010",7560 => "10001011",7561 => "00010111",7562 => "10010011",7563 => "11001011",7564 => "01100111",7565 => "00000011",7566 => "01000001",7567 => "11011100",7568 => "00001000",7569 => "00001100",7570 => "01011110",7571 => "00101111",7572 => "01101010",7573 => "00001000",7574 => "11110111",7575 => "00000011",7576 => "00100110",7577 => "01110110",7578 => "00011010",7579 => "11111010",7580 => "00100010",7581 => "11001111",7582 => "01010000",7583 => "10111100",7584 => "00101011",7585 => "00111000",7586 => "11010001",7587 => "10111010",7588 => "00110011",7589 => "10111001",7590 => "11001101",7591 => "11100011",7592 => "00010001",7593 => "10011011",7594 => "11001000",7595 => "01001010",7596 => "11010010",7597 => "10100010",7598 => "00000010",7599 => "10010000",7600 => "10111001",7601 => "00100110",7602 => "01111101",7603 => "11010000",7604 => "00001001",7605 => "00011001",7606 => "11111100",7607 => "00010011",7608 => "10100101",7609 => "10011100",7610 => "10001001",7611 => "11000011",7612 => "11101100",7613 => "01010110",7614 => "01101111",7615 => "11000000",7616 => "11001100",7617 => "00111110",7618 => "00101011",7619 => "00011101",7620 => "10101110",7621 => "11011000",7622 => "00001000",7623 => "01110110",7624 => "00010001",7625 => "11101000",7626 => "11100011",7627 => "10001101",7628 => "10110010",7629 => "11011110",7630 => "00010010",7631 => "00010101",7632 => "01010111",7633 => "11110100",7634 => "00100011",7635 => "10110010",7636 => "11001110",7637 => "00101001",7638 => "11000010",7639 => "11110110",7640 => "01100101",7641 => "10000010",7642 => "00111110",7643 => "00101111",7644 => "10000001",7645 => "01111101",7646 => "01101010",7647 => "00101011",7648 => "01100010",7649 => "00111100",7650 => "11110000",7651 => "01100101",7652 => "01101110",7653 => "10100011",7654 => "11001100",7655 => "10000001",7656 => "10100110",7657 => "01101001",7658 => "10110111",7659 => "11000110",7660 => "11011110",7661 => "00001110",7662 => "11000001",7663 => "11101110",7664 => "00010011",7665 => "10001100",7666 => "01100100",7667 => "01000011",7668 => "00111011",7669 => "11101011",7670 => "10110100",7671 => "00100010",7672 => "10000101",7673 => "00100000",7674 => "10101000",7675 => "10101101",7676 => "00101011",7677 => "00110000",7678 => "00110101",7679 => "10001001",7680 => "10110110",7681 => "01111001",7682 => "10110101",7683 => "01111111",7684 => "00010010",7685 => "01111111",7686 => "11111001",7687 => "10010111",7688 => "01100110",7689 => "01001101",7690 => "10100110",7691 => "00101010",7692 => "00000110",7693 => "10111100",7694 => "00000000",7695 => "10001000",7696 => "01000001",7697 => "11000111",7698 => "00010111",7699 => "00100100",7700 => "11010101",7701 => "00110000",7702 => "01001001",7703 => "01100000",7704 => "10001111",7705 => "00011110",7706 => "01011010",7707 => "00100100",7708 => "11100110",7709 => "10010000",7710 => "10011001",7711 => "00100011",7712 => "10101001",7713 => "00011011",7714 => "01101111",7715 => "10111011",7716 => "01101001",7717 => "01101111",7718 => "00011100",7719 => "00101011",7720 => "10011101",7721 => "00010001",7722 => "11011010",7723 => "11010001",7724 => "11011010",7725 => "10110110",7726 => "01100100",7727 => "01000100",7728 => "00001100",7729 => "00111111",7730 => "00110111",7731 => "00001111",7732 => "01010011",7733 => "01111101",7734 => "10010110",7735 => "11001010",7736 => "11100101",7737 => "01001010",7738 => "01011000",7739 => "00011001",7740 => "01010010",7741 => "10011100",7742 => "10101110",7743 => "01110111",7744 => "11111000",7745 => "00101010",7746 => "10111101",7747 => "11010010",7748 => "00001011",7749 => "00001110",7750 => "00011100",7751 => "00111100",7752 => "11110010",7753 => "11000000",7754 => "01001001",7755 => "00100100",7756 => "00110010",7757 => "10001011",7758 => "10111010",7759 => "10000111",7760 => "11011011",7761 => "11101001",7762 => "10000001",7763 => "11111000",7764 => "11111110",7765 => "11010100",7766 => "11000111",7767 => "01111000",7768 => "10110110",7769 => "00001000",7770 => "11100010",7771 => "01101011",7772 => "10100011",7773 => "10101110",7774 => "10001111",7775 => "11011111",7776 => "10011011",7777 => "11110000",7778 => "01111111",7779 => "11110001",7780 => "01011000",7781 => "00111111",7782 => "00111010",7783 => "11101101",7784 => "11010101",7785 => "10001101",7786 => "00110110",7787 => "11111111",7788 => "10001101",7789 => "00000010",7790 => "01101110",7791 => "11111110",7792 => "00001010",7793 => "10011011",7794 => "01110110",7795 => "00010101",7796 => "00101001",7797 => "10011011",7798 => "10011111",7799 => "10001010",7800 => "01100100",7801 => "00001001",7802 => "00100100",7803 => "01011001",7804 => "00000110",7805 => "01000001",7806 => "00111110",7807 => "00110100",7808 => "10111011",7809 => "10001001",7810 => "00011011",7811 => "00010000",7812 => "00110000",7813 => "01010111",7814 => "11010101",7815 => "01100100",7816 => "01100110",7817 => "10011001",7818 => "01101000",7819 => "01110110",7820 => "01111110",7821 => "10001000",7822 => "00001001",7823 => "10001110",7824 => "10110111",7825 => "10110111",7826 => "11010000",7827 => "00010001",7828 => "11110110",7829 => "00010110",7830 => "10100101",7831 => "01110010",7832 => "01010011",7833 => "00110011",7834 => "01100011",7835 => "10000011",7836 => "00111010",7837 => "00000101",7838 => "11110100",7839 => "00111100",7840 => "10101010",7841 => "00010001",7842 => "11010101",7843 => "01111011",7844 => "10001110",7845 => "01010100",7846 => "10010100",7847 => "11100100",7848 => "11111110",7849 => "01001101",7850 => "01100100",7851 => "00010011",7852 => "01110101",7853 => "00000001",7854 => "10110111",7855 => "01000110",7856 => "01101111",7857 => "00100011",7858 => "01110100",7859 => "01111011",7860 => "01100001",7861 => "11011110",7862 => "11000111",7863 => "10100111",7864 => "11101111",7865 => "01101011",7866 => "10000110",7867 => "10000100",7868 => "10011010",7869 => "11011100",7870 => "01101011",7871 => "01011110",7872 => "01100011",7873 => "01111001",7874 => "01101110",7875 => "10011010",7876 => "01001011",7877 => "01111000",7878 => "11111101",7879 => "11100111",7880 => "11001101",7881 => "10111001",7882 => "00110100",7883 => "11101001",7884 => "11011001",7885 => "11110001",7886 => "10111111",7887 => "10000111",7888 => "01100000",7889 => "11110110",7890 => "01100000",7891 => "10101001",7892 => "10110101",7893 => "00010100",7894 => "10011110",7895 => "01000101",7896 => "10001000",7897 => "01101011",7898 => "01101110",7899 => "01110010",7900 => "00001110",7901 => "00011100",7902 => "01101110",7903 => "11101101",7904 => "11100110",7905 => "00101110",7906 => "10100011",7907 => "11101101",7908 => "00001001",7909 => "00011111",7910 => "10101101",7911 => "01100110",7912 => "01011100",7913 => "00100101",7914 => "10001010",7915 => "11000110",7916 => "10100011",7917 => "00010001",7918 => "01101010",7919 => "01101111",7920 => "10110111",7921 => "01111110",7922 => "11100100",7923 => "01010111",7924 => "11101000",7925 => "10010101",7926 => "10110011",7927 => "01110011",7928 => "01011110",7929 => "10010111",7930 => "00000000",7931 => "01001000",7932 => "11101000",7933 => "01111111",7934 => "10111100",7935 => "11011011",7936 => "00111111",7937 => "01110101",7938 => "00101010",7939 => "00100000",7940 => "11011001",7941 => "10110011",7942 => "11010000",7943 => "01100010",7944 => "10000100",7945 => "10000111",7946 => "00000011",7947 => "11100011",7948 => "11110010",7949 => "01101010",7950 => "10100011",7951 => "01100111",7952 => "11011110",7953 => "00010001",7954 => "01100001",7955 => "11100011",7956 => "01000010",7957 => "10100101",7958 => "11011101",7959 => "11011101",7960 => "00011010",7961 => "10100011",7962 => "10110110",7963 => "10000010",7964 => "00010100",7965 => "01000010",7966 => "00101101",7967 => "11110100",7968 => "11001010",7969 => "10010000",7970 => "00110111",7971 => "11001110",7972 => "11000000",7973 => "11101010",7974 => "00110110",7975 => "11001101",7976 => "11011111",7977 => "11101110",7978 => "01001111",7979 => "00100100",7980 => "10011101",7981 => "11001111",7982 => "10101000",7983 => "11001010",7984 => "10000001",7985 => "00010110",7986 => "00100110",7987 => "10111110",7988 => "11101011",7989 => "10100110",7990 => "00100011",7991 => "10001110",7992 => "00100110",7993 => "10001000",7994 => "00110010",7995 => "01011010",7996 => "10000101",7997 => "11111010",7998 => "01100010",7999 => "10001010",8000 => "11001010",8001 => "01100101",8002 => "10111001",8003 => "00010100",8004 => "01101001",8005 => "10000110",8006 => "10111010",8007 => "00111110",8008 => "01001001",8009 => "00100010",8010 => "10001001",8011 => "11101111",8012 => "10111001",8013 => "11110010",8014 => "11011111",8015 => "11001001",8016 => "00101011",8017 => "00000010",8018 => "00011000",8019 => "11101001",8020 => "10111011",8021 => "00001101",8022 => "11111111",8023 => "10101000",8024 => "01111110",8025 => "00010011",8026 => "11011111",8027 => "01101000",8028 => "01101111",8029 => "10011010",8030 => "01101110",8031 => "11101111",8032 => "11001101",8033 => "10001000",8034 => "11000011",8035 => "11000111",8036 => "00010011",8037 => "10110100",8038 => "10011011",8039 => "11010001",8040 => "01011111",8041 => "10001100",8042 => "10000100",8043 => "10010001",8044 => "01010110",8045 => "01110010",8046 => "00101101",8047 => "11001111",8048 => "11001001",8049 => "10101101",8050 => "01001110",8051 => "00100001",8052 => "01011011",8053 => "01101111",8054 => "00000010",8055 => "11110010",8056 => "00100101",8057 => "01010001",8058 => "10111001",8059 => "10100010",8060 => "11110101",8061 => "11010110",8062 => "00010010",8063 => "00110101",8064 => "01101111",8065 => "00111011",8066 => "00010001",8067 => "10001100",8068 => "01000010",8069 => "01101010",8070 => "00001100",8071 => "01111010",8072 => "10110110",8073 => "11110011",8074 => "10100001",8075 => "00100111",8076 => "00110010",8077 => "10111011",8078 => "00000010",8079 => "01101010",8080 => "01110110",8081 => "01101110",8082 => "10100001",8083 => "01001001",8084 => "11111110",8085 => "11111101",8086 => "10110011",8087 => "10101000",8088 => "10110110",8089 => "11110111",8090 => "11110001",8091 => "00000000",8092 => "11111100",8093 => "11000100",8094 => "00000000",8095 => "11101111",8096 => "01011101",8097 => "11000111",8098 => "10011110",8099 => "11001011",8100 => "01111000",8101 => "00000110",8102 => "11100111",8103 => "01100111",8104 => "11010111",8105 => "11110100",8106 => "00010010",8107 => "10001010",8108 => "10100000",8109 => "10101011",8110 => "10001110",8111 => "01110100",8112 => "00000010",8113 => "11101010",8114 => "00010111",8115 => "10011000",8116 => "10000001",8117 => "10010101",8118 => "11011000",8119 => "01111100",8120 => "10101001",8121 => "00101110",8122 => "10110111",8123 => "11011111",8124 => "11001011",8125 => "01011001",8126 => "11110010",8127 => "00101011",8128 => "00011001",8129 => "00111010",8130 => "00101101",8131 => "11010010",8132 => "10111000",8133 => "00101110",8134 => "11111000",8135 => "01101001",8136 => "11000100",8137 => "00000001",8138 => "01101100",8139 => "10001010",8140 => "01011000",8141 => "10101011",8142 => "10000111",8143 => "10010101",8144 => "01000000",8145 => "10010100",8146 => "11001101",8147 => "00001001",8148 => "10010110",8149 => "10010011",8150 => "00111111",8151 => "11001100",8152 => "00100101",8153 => "11101111",8154 => "01000001",8155 => "10000010",8156 => "01000011",8157 => "10000000",8158 => "00101010",8159 => "11110101",8160 => "10111011",8161 => "01110111",8162 => "00010101",8163 => "11100110",8164 => "11001001",8165 => "00111001",8166 => "11000110",8167 => "11001110",8168 => "10110110",8169 => "01000000",8170 => "01101101",8171 => "10000100",8172 => "11111011",8173 => "01000000",8174 => "11010000",8175 => "10010000",8176 => "01100110",8177 => "01000111",8178 => "01101101",8179 => "10011000",8180 => "01101001",8181 => "10100111",8182 => "11011011",8183 => "10101101",8184 => "10000111",8185 => "10111010",8186 => "01011000",8187 => "10011001",8188 => "10101111",8189 => "00100101",8190 => "00000100",8191 => "10000100",8192 => "10100011",8193 => "11011000",8194 => "11110110",8195 => "10100100",8196 => "10000000",8197 => "10000110",8198 => "00011111",8199 => "11111100",8200 => "10100011",8201 => "10001110",8202 => "11011100",8203 => "00011011",8204 => "00100111",8205 => "11000001",8206 => "00111110",8207 => "11000001",8208 => "11101110",8209 => "11101100",8210 => "10100101",8211 => "00011000",8212 => "01101111",8213 => "01101011",8214 => "10011100",8215 => "00000001",8216 => "10001111",8217 => "10001100",8218 => "00101001",8219 => "01010100",8220 => "01001101",8221 => "11001111",8222 => "00010001",8223 => "01110010",8224 => "00111110",8225 => "11001011",8226 => "10010001",8227 => "01101101",8228 => "00001000",8229 => "10001001",8230 => "10001001",8231 => "01011111",8232 => "00011111",8233 => "00111100",8234 => "00011110",8235 => "01011010",8236 => "10010111",8237 => "11001010",8238 => "11000110",8239 => "00011011",8240 => "00110000",8241 => "01010111",8242 => "01101111",8243 => "10111001",8244 => "11110011",8245 => "11111010",8246 => "00000011",8247 => "11111110",8248 => "00000011",8249 => "00000101",8250 => "01000111",8251 => "01011010",8252 => "00010101",8253 => "00100011",8254 => "10101111",8255 => "00110010",8256 => "11110000",8257 => "00011010",8258 => "00101010",8259 => "01100011",8260 => "00010000",8261 => "10111101",8262 => "11000011",8263 => "10100010",8264 => "10001110",8265 => "11000000",8266 => "00110010",8267 => "01010001",8268 => "11101111",8269 => "00101110",8270 => "10100000",8271 => "10001000",8272 => "10100011",8273 => "10010110",8274 => "01010001",8275 => "00101101",8276 => "10011100",8277 => "10100100",8278 => "11011100",8279 => "01011101",8280 => "11111001",8281 => "11101010",8282 => "11000011",8283 => "11011011",8284 => "11101001",8285 => "01010000",8286 => "01011010",8287 => "01000111",8288 => "10111100",8289 => "10000111",8290 => "10011111",8291 => "10111100",8292 => "11001110",8293 => "11010100",8294 => "00101100",8295 => "10101110",8296 => "00010001",8297 => "01111101",8298 => "11010010",8299 => "11100111",8300 => "00101000",8301 => "01011100",8302 => "11110011",8303 => "11011000",8304 => "00100101",8305 => "01010100",8306 => "00101100",8307 => "11100100",8308 => "11011111",8309 => "11111110",8310 => "00100010",8311 => "01101001",8312 => "10000000",8313 => "00100111",8314 => "00011111",8315 => "00111011",8316 => "01111000",8317 => "01100010",8318 => "11100011",8319 => "01000011",8320 => "00101110",8321 => "01101111",8322 => "01110011",8323 => "00010011",8324 => "11011010",8325 => "01001010",8326 => "01101000",8327 => "00011011",8328 => "10001101",8329 => "00010101",8330 => "00011100",8331 => "11101100",8332 => "01011011",8333 => "00111110",8334 => "00011101",8335 => "01101011",8336 => "01111110",8337 => "11010111",8338 => "01101100",8339 => "10000010",8340 => "01000100",8341 => "01101111",8342 => "01011001",8343 => "10100101",8344 => "11111010",8345 => "00011001",8346 => "01101010",8347 => "11011000",8348 => "00000100",8349 => "01010010",8350 => "01101100",8351 => "00011010",8352 => "11010011",8353 => "11011011",8354 => "10011010",8355 => "11101000",8356 => "01100000",8357 => "10010001",8358 => "11110010",8359 => "00010010",8360 => "10000010",8361 => "00010000",8362 => "10101000",8363 => "11101110",8364 => "00101011",8365 => "00011000",8366 => "10111010",8367 => "00100110",8368 => "00001001",8369 => "00011010",8370 => "10000111",8371 => "00101001",8372 => "00110011",8373 => "11001010",8374 => "11111110",8375 => "11111111",8376 => "00100000",8377 => "00111011",8378 => "00011011",8379 => "00000100",8380 => "10110111",8381 => "11010010",8382 => "11011001",8383 => "00010110",8384 => "11111111",8385 => "11000000",8386 => "01110010",8387 => "00011010",8388 => "11001001",8389 => "01001000",8390 => "10000000",8391 => "01000010",8392 => "01110101",8393 => "11101001",8394 => "00001010",8395 => "01110111",8396 => "01011101",8397 => "00010011",8398 => "10000101",8399 => "11100101",8400 => "01111011",8401 => "10100000",8402 => "11000100",8403 => "11010100",8404 => "01011111",8405 => "10100011",8406 => "10110100",8407 => "01001000",8408 => "11010011",8409 => "11000110",8410 => "10110011",8411 => "01101101",8412 => "01001010",8413 => "00101010",8414 => "11001110",8415 => "10110101",8416 => "00011001",8417 => "01111101",8418 => "10100001",8419 => "00111000",8420 => "11000110",8421 => "00010000",8422 => "00101111",8423 => "01110111",8424 => "11000000",8425 => "10011001",8426 => "01110101",8427 => "10110010",8428 => "11110110",8429 => "00101110",8430 => "01000010",8431 => "10000011",8432 => "01110010",8433 => "00001110",8434 => "10010000",8435 => "01110110",8436 => "11011001",8437 => "01101010",8438 => "01001100",8439 => "11101000",8440 => "11111010",8441 => "11000010",8442 => "10101001",8443 => "00110101",8444 => "00100111",8445 => "11100011",8446 => "10111100",8447 => "10000011",8448 => "10110101",8449 => "10001011",8450 => "01100100",8451 => "11110000",8452 => "10101111",8453 => "10110111",8454 => "10111110",8455 => "01111001",8456 => "11011100",8457 => "00110000",8458 => "10101111",8459 => "01110011",8460 => "10100111",8461 => "10100010",8462 => "00010111",8463 => "01101000",8464 => "11111101",8465 => "00111010",8466 => "00110001",8467 => "01011001",8468 => "01110101",8469 => "01111101",8470 => "10100000",8471 => "00000101",8472 => "01011110",8473 => "00101101",8474 => "00011100",8475 => "00000000",8476 => "01011100",8477 => "10111110",8478 => "00010010",8479 => "01011011",8480 => "00101010",8481 => "11001110",8482 => "00001000",8483 => "11100110",8484 => "10101100",8485 => "11010001",8486 => "00101000",8487 => "10110010",8488 => "10111011",8489 => "10110110",8490 => "11100011",8491 => "01000010",8492 => "00101101",8493 => "10011110",8494 => "10011011",8495 => "11011001",8496 => "01000001",8497 => "00010011",8498 => "11100101",8499 => "11100001",8500 => "10001010",8501 => "11000010",8502 => "11101000",8503 => "11111110",8504 => "01111101",8505 => "11001101",8506 => "00011111",8507 => "00101000",8508 => "11010010",8509 => "01001001",8510 => "00110100",8511 => "00111010",8512 => "11110001",8513 => "00000111",8514 => "11101011",8515 => "01010011",8516 => "00001100",8517 => "11111011",8518 => "01000101",8519 => "00001000",8520 => "00100100",8521 => "11000001",8522 => "10101000",8523 => "11111010",8524 => "10100000",8525 => "11001011",8526 => "10010110",8527 => "11011011",8528 => "00000110",8529 => "11000111",8530 => "10010010",8531 => "00001010",8532 => "01101100",8533 => "01100111",8534 => "11010101",8535 => "10101101",8536 => "11010010",8537 => "10110111",8538 => "00000000",8539 => "10000010",8540 => "11001111",8541 => "11100100",8542 => "10010010",8543 => "10000111",8544 => "00110100",8545 => "00100000",8546 => "00111010",8547 => "10101110",8548 => "10110001",8549 => "01110010",8550 => "01010010",8551 => "00111001",8552 => "01110011",8553 => "11001101",8554 => "11111010",8555 => "11100101",8556 => "11011001",8557 => "00110111",8558 => "10001110",8559 => "10000000",8560 => "11111011",8561 => "10011010",8562 => "00010110",8563 => "01010000",8564 => "00000111",8565 => "10101011",8566 => "01110011",8567 => "11010110",8568 => "10011000",8569 => "00110101",8570 => "11010011",8571 => "01111111",8572 => "00110110",8573 => "11111110",8574 => "10010111",8575 => "01110010",8576 => "10010111",8577 => "10100011",8578 => "11000011",8579 => "11000000",8580 => "00110110",8581 => "11101000",8582 => "00010100",8583 => "00000101",8584 => "10011010",8585 => "01000011",8586 => "00001111",8587 => "00110110",8588 => "10010101",8589 => "01011100",8590 => "10101001",8591 => "00111111",8592 => "10111011",8593 => "00010010",8594 => "00101100",8595 => "00001101",8596 => "10100001",8597 => "00011100",8598 => "01100010",8599 => "00101110",8600 => "01100101",8601 => "00010000",8602 => "10101101",8603 => "11101100",8604 => "00000011",8605 => "00100100",8606 => "01011000",8607 => "01011110",8608 => "00101011",8609 => "10010000",8610 => "11111001",8611 => "11111110",8612 => "11000001",8613 => "10001100",8614 => "10000101",8615 => "00000111",8616 => "01010011",8617 => "10000110",8618 => "00101101",8619 => "10000011",8620 => "10111100",8621 => "10111110",8622 => "11001100",8623 => "00110011",8624 => "01010000",8625 => "00001101",8626 => "00100111",8627 => "11101011",8628 => "00101000",8629 => "11011101",8630 => "00100010",8631 => "11110101",8632 => "11100111",8633 => "10111001",8634 => "11101010",8635 => "00001101",8636 => "11101101",8637 => "11110111",8638 => "01000010",8639 => "00000000",8640 => "10001100",8641 => "11110001",8642 => "10001110",8643 => "10000000",8644 => "00110000",8645 => "11111011",8646 => "01000100",8647 => "11110011",8648 => "00011000",8649 => "11111010",8650 => "00001000",8651 => "00101011",8652 => "10010000",8653 => "10001100",8654 => "11010011",8655 => "10101000",8656 => "10001001",8657 => "11111111",8658 => "11000011",8659 => "11011000",8660 => "00100001",8661 => "11110100",8662 => "10010111",8663 => "11000110",8664 => "11101000",8665 => "10010111",8666 => "01100001",8667 => "01000001",8668 => "11000011",8669 => "11001101",8670 => "00001001",8671 => "00111100",8672 => "10100111",8673 => "10100010",8674 => "11110111",8675 => "01010001",8676 => "11100110",8677 => "11101000",8678 => "01100100",8679 => "01001001",8680 => "00010010",8681 => "00000111",8682 => "00110110",8683 => "10001101",8684 => "01101010",8685 => "10000111",8686 => "00111111",8687 => "10001110",8688 => "01010110",8689 => "00010100",8690 => "10111101",8691 => "00100111",8692 => "00110010",8693 => "01001101",8694 => "00100000",8695 => "10111000",8696 => "00010011",8697 => "01111110",8698 => "11010011",8699 => "00111101",8700 => "00111100",8701 => "00010111",8702 => "00000011",8703 => "11011010",8704 => "01000111",8705 => "01110100",8706 => "10100101",8707 => "00110000",8708 => "11001000",8709 => "11001111",8710 => "10100001",8711 => "11101001",8712 => "10000000",8713 => "00110100",8714 => "11100000",8715 => "11110100",8716 => "10000111",8717 => "10011001",8718 => "01111111",8719 => "00110001",8720 => "11111100",8721 => "10101000",8722 => "00001111",8723 => "10100101",8724 => "01001100",8725 => "11000110",8726 => "00101111",8727 => "00100000",8728 => "01101100",8729 => "11001101",8730 => "01100100",8731 => "00010010",8732 => "11011100",8733 => "01100110",8734 => "01100111",8735 => "10011100",8736 => "11000000",8737 => "00001010",8738 => "00000110",8739 => "01011011",8740 => "00001010",8741 => "10011000",8742 => "11011101",8743 => "00110101",8744 => "11111010",8745 => "01011000",8746 => "10110010",8747 => "11111110",8748 => "10111101",8749 => "11000111",8750 => "10100110",8751 => "10001101",8752 => "10100010",8753 => "01100100",8754 => "01010011",8755 => "10100010",8756 => "00110010",8757 => "00100000",8758 => "00110110",8759 => "10001111",8760 => "11111001",8761 => "10110011",8762 => "11001000",8763 => "00111010",8764 => "01101110",8765 => "11000010",8766 => "11100101",8767 => "10010011",8768 => "10011011",8769 => "11111011",8770 => "11011100",8771 => "01010010",8772 => "00111011",8773 => "10011011",8774 => "11111000",8775 => "00001110",8776 => "11010000",8777 => "11010001",8778 => "00010011",8779 => "11111001",8780 => "10000011",8781 => "11101111",8782 => "11011101",8783 => "01111110",8784 => "00010000",8785 => "01110100",8786 => "00001001",8787 => "00100110",8788 => "10100111",8789 => "01011110",8790 => "01110101",8791 => "11101010",8792 => "11111010",8793 => "01001001",8794 => "11010110",8795 => "01101111",8796 => "10101010",8797 => "10011001",8798 => "11100000",8799 => "00101100",8800 => "11100101",8801 => "10111000",8802 => "11101000",8803 => "11000000",8804 => "01010000",8805 => "00111011",8806 => "11110000",8807 => "01011001",8808 => "01100011",8809 => "11100110",8810 => "00001001",8811 => "00001111",8812 => "01000110",8813 => "10110110",8814 => "01000001",8815 => "11011011",8816 => "10110000",8817 => "11110111",8818 => "10010100",8819 => "00000010",8820 => "00101010",8821 => "01100000",8822 => "00000111",8823 => "01101000",8824 => "01101110",8825 => "11001000",8826 => "00100010",8827 => "00011111",8828 => "10000110",8829 => "11101110",8830 => "00011010",8831 => "01010011",8832 => "11100110",8833 => "11111001",8834 => "10111010",8835 => "11110011",8836 => "00111000",8837 => "00001011",8838 => "11011001",8839 => "11111000",8840 => "10101010",8841 => "00100111",8842 => "00010010",8843 => "11001101",8844 => "00000111",8845 => "11101100",8846 => "00110011",8847 => "10000111",8848 => "00000011",8849 => "10010010",8850 => "10011110",8851 => "01110110",8852 => "01010100",8853 => "10111011",8854 => "11010110",8855 => "01000001",8856 => "00101011",8857 => "11010100",8858 => "00111100",8859 => "11101011",8860 => "00011000",8861 => "00101111",8862 => "01000001",8863 => "01110111",8864 => "10011111",8865 => "11111001",8866 => "01000000",8867 => "11010001",8868 => "11010001",8869 => "01010110",8870 => "10001011",8871 => "10010101",8872 => "00011000",8873 => "11100101",8874 => "11110111",8875 => "00010000",8876 => "10101110",8877 => "11110000",8878 => "00001010",8879 => "01101011",8880 => "10111110",8881 => "01011101",8882 => "10011110",8883 => "00101110",8884 => "11101100",8885 => "11100101",8886 => "01111010",8887 => "01000000",8888 => "10101101",8889 => "01010110",8890 => "01110110",8891 => "11000110",8892 => "00010000",8893 => "11111100",8894 => "00000100",8895 => "11011000",8896 => "01100110",8897 => "10011010",8898 => "00110010",8899 => "01111110",8900 => "11011011",8901 => "11010111",8902 => "00101101",8903 => "10000011",8904 => "01100001",8905 => "00010100",8906 => "11100011",8907 => "00101100",8908 => "11001011",8909 => "11001000",8910 => "10100110",8911 => "01010110",8912 => "10010101",8913 => "01011010",8914 => "01011010",8915 => "00011000",8916 => "11010100",8917 => "01101010",8918 => "10000000",8919 => "11010101",8920 => "11011000",8921 => "11110001",8922 => "10110010",8923 => "01111001",8924 => "00000111",8925 => "10110101",8926 => "10111100",8927 => "10010110",8928 => "11101111",8929 => "11110101",8930 => "00010101",8931 => "01100111",8932 => "00001100",8933 => "11001110",8934 => "01100001",8935 => "01101111",8936 => "00001011",8937 => "11000111",8938 => "11010011",8939 => "00001011",8940 => "11101011",8941 => "10100001",8942 => "10010100",8943 => "01100111",8944 => "00110000",8945 => "00000001",8946 => "10100011",8947 => "00101100",8948 => "10010111",8949 => "00110010",8950 => "10110110",8951 => "10100011",8952 => "10110010",8953 => "10101011",8954 => "01111111",8955 => "01100001",8956 => "10000111",8957 => "01111111",8958 => "11110001",8959 => "11010010",8960 => "00000011",8961 => "10001001",8962 => "01010111",8963 => "01111110",8964 => "01100111",8965 => "10001111",8966 => "10100011",8967 => "10001100",8968 => "11011001",8969 => "10010000",8970 => "00101111",8971 => "11110011",8972 => "11110011",8973 => "10010100",8974 => "01100100",8975 => "10111001",8976 => "01110001",8977 => "11111011",8978 => "00110110",8979 => "11010110",8980 => "01100001",8981 => "11011000",8982 => "10010001",8983 => "00100110",8984 => "00100010",8985 => "00100110",8986 => "01010010",8987 => "00001000",8988 => "10101100",8989 => "00110010",8990 => "11011110",8991 => "00101111",8992 => "11000000",8993 => "10000010",8994 => "00011011",8995 => "11010011",8996 => "11001101",8997 => "01111111",8998 => "10001100",8999 => "10010001",9000 => "00011001",9001 => "01010100",9002 => "10011100",9003 => "11000110",9004 => "01000101",9005 => "11011100",9006 => "10100110",9007 => "11001111",9008 => "01111100",9009 => "10011110",9010 => "10000111",9011 => "10100001",9012 => "01000010",9013 => "00000111",9014 => "10001011",9015 => "11000011",9016 => "01101100",9017 => "10101100",9018 => "11110001",9019 => "10000001",9020 => "00011000",9021 => "10000110",9022 => "00011010",9023 => "11111111",9024 => "00010101",9025 => "00000000",9026 => "00001010",9027 => "01011101",9028 => "01101011",9029 => "11010010",9030 => "01011101",9031 => "00111000",9032 => "01100000",9033 => "00101011",9034 => "01010101",9035 => "01111010",9036 => "10011110",9037 => "10011010",9038 => "01010110",9039 => "01110100",9040 => "01101110",9041 => "10000010",9042 => "01111101",9043 => "11011101",9044 => "11111101",9045 => "00100111",9046 => "11101110",9047 => "10101111",9048 => "00000000",9049 => "01110111",9050 => "10110110",9051 => "01011010",9052 => "01010111",9053 => "01001011",9054 => "11110111",9055 => "10000100",9056 => "10001000",9057 => "11110011",9058 => "10000100",9059 => "10100010",9060 => "10101110",9061 => "01011101",9062 => "00100111",9063 => "10100100",9064 => "00111101",9065 => "00011111",9066 => "10110010",9067 => "01011010",9068 => "00111111",9069 => "11110101",9070 => "11100011",9071 => "10011110",9072 => "00010110",9073 => "01111101",9074 => "00010100",9075 => "10110111",9076 => "01001001",9077 => "10001001",9078 => "00000100",9079 => "00011011",9080 => "00101111",9081 => "11011101",9082 => "11100011",9083 => "10011001",9084 => "00101100",9085 => "01100100",9086 => "10100010",9087 => "11001011",9088 => "10011010",9089 => "10000010",9090 => "10010100",9091 => "11101111",9092 => "10100000",9093 => "10110001",9094 => "00101011",9095 => "11010111",9096 => "11101010",9097 => "01000111",9098 => "11100000",9099 => "11011011",9100 => "00100011",9101 => "10110100",9102 => "11011010",9103 => "10100110",9104 => "10001001",9105 => "10001001",9106 => "10010100",9107 => "11010111",9108 => "10101100",9109 => "11111100",9110 => "01001100",9111 => "00001001",9112 => "10001010",9113 => "10110011",9114 => "10111111",9115 => "01111011",9116 => "11010010",9117 => "00101111",9118 => "01101100",9119 => "11111111",9120 => "00110001",9121 => "11001011",9122 => "00101100",9123 => "00011001",9124 => "01111000",9125 => "11101000",9126 => "10111010",9127 => "00111110",9128 => "10101010",9129 => "10011001",9130 => "01010101",9131 => "00111000",9132 => "10010101",9133 => "10000100",9134 => "01101100",9135 => "11100001",9136 => "10111011",9137 => "00000000",9138 => "01000011",9139 => "00101111",9140 => "10110110",9141 => "00100110",9142 => "00100000",9143 => "11001101",9144 => "01011101",9145 => "11101110",9146 => "01101011",9147 => "10100011",9148 => "11100100",9149 => "00100101",9150 => "10111100",9151 => "11000101",9152 => "11110111",9153 => "00100010",9154 => "01010101",9155 => "01000001",9156 => "00110110",9157 => "10111101",9158 => "10111001",9159 => "00000111",9160 => "10001001",9161 => "01010010",9162 => "10000110",9163 => "11101111",9164 => "10101111",9165 => "01001110",9166 => "11101101",9167 => "11011011",9168 => "01110000",9169 => "01010101",9170 => "00010110",9171 => "10101110",9172 => "11101000",9173 => "00010110",9174 => "00100100",9175 => "01100010",9176 => "10100111",9177 => "00110001",9178 => "00111001",9179 => "00000000",9180 => "00111000",9181 => "10100100",9182 => "10110011",9183 => "01001101",9184 => "10100011",9185 => "01001000",9186 => "00001100",9187 => "11110101",9188 => "10011010",9189 => "10010110",9190 => "11110001",9191 => "10101001",9192 => "01001000",9193 => "01001101",9194 => "11011000",9195 => "00000111",9196 => "10000100",9197 => "00111001",9198 => "01100100",9199 => "00001000",9200 => "10101011",9201 => "00100101",9202 => "10101111",9203 => "00010001",9204 => "01110011",9205 => "00011001",9206 => "11011011",9207 => "11001111",9208 => "10010011",9209 => "00010010",9210 => "10100101",9211 => "11011100",9212 => "01011000",9213 => "01100011",9214 => "01101011",9215 => "01111010",9216 => "01011000",9217 => "10101011",9218 => "00000011",9219 => "10011010",9220 => "10101000",9221 => "01001000",9222 => "10011001",9223 => "11010011",9224 => "11100111",9225 => "00000110",9226 => "11001010",9227 => "11101000",9228 => "11000010",9229 => "10110001",9230 => "00101001",9231 => "10110010",9232 => "10111100",9233 => "11101111",9234 => "00100010",9235 => "00001100",9236 => "00001100",9237 => "11011111",9238 => "10000101",9239 => "00101101",9240 => "10001000",9241 => "11010101",9242 => "10000011",9243 => "00000100",9244 => "11110101",9245 => "00100110",9246 => "01111010",9247 => "01001101",9248 => "00011101",9249 => "01010010",9250 => "01010001",9251 => "10111000",9252 => "10011110",9253 => "01110110",9254 => "10001010",9255 => "10010111",9256 => "11001010",9257 => "00011011",9258 => "10111011",9259 => "11010111",9260 => "00001100",9261 => "11011110",9262 => "11011110",9263 => "00101000",9264 => "10000100",9265 => "00111011",9266 => "00010001",9267 => "11110110",9268 => "00100001",9269 => "00010011",9270 => "10000111",9271 => "01101101",9272 => "00000101",9273 => "01110111",9274 => "11010001",9275 => "00110010",9276 => "11111110",9277 => "00010100",9278 => "10010101",9279 => "10000100",9280 => "01001010",9281 => "01110011",9282 => "00001101",9283 => "01111000",9284 => "00100100",9285 => "10100111",9286 => "00011011",9287 => "00001111",9288 => "01010000",9289 => "01100111",9290 => "10100001",9291 => "11111110",9292 => "11100100",9293 => "11001110",9294 => "11011001",9295 => "10111000",9296 => "00011011",9297 => "01011000",9298 => "00101001",9299 => "11001011",9300 => "10001101",9301 => "01010000",9302 => "11111111",9303 => "00111000",9304 => "10000101",9305 => "11101011",9306 => "11010001",9307 => "00010110",9308 => "01101010",9309 => "11000011",9310 => "11000110",9311 => "10111101",9312 => "11001001",9313 => "00110100",9314 => "10010001",9315 => "10000110",9316 => "00101011",9317 => "11111111",9318 => "10111101",9319 => "10100011",9320 => "11101101",9321 => "10001110",9322 => "00000111",9323 => "01000111",9324 => "11101011",9325 => "00001001",9326 => "11100001",9327 => "00111101",9328 => "01010011",9329 => "00111001",9330 => "01000011",9331 => "01011110",9332 => "00011110",9333 => "11011010",9334 => "10010111",9335 => "01100000",9336 => "11011011",9337 => "11100010",9338 => "01001000",9339 => "00110101",9340 => "00100011",9341 => "01101100",9342 => "10011110",9343 => "11001001",9344 => "11011110",9345 => "10000101",9346 => "11101010",9347 => "00111101",9348 => "11111110",9349 => "10110100",9350 => "10010110",9351 => "10100110",9352 => "11101100",9353 => "11100010",9354 => "01110101",9355 => "01010011",9356 => "01001100",9357 => "01111010",9358 => "11111001",9359 => "11111110",9360 => "01111111",9361 => "00110011",9362 => "00111111",9363 => "11000000",9364 => "11011010",9365 => "10000101",9366 => "00101010",9367 => "00110100",9368 => "10000100",9369 => "10101110",9370 => "10001101",9371 => "11110100",9372 => "11110111",9373 => "01110011",9374 => "10110110",9375 => "10011101",9376 => "10110101",9377 => "00101101",9378 => "00001110",9379 => "10010100",9380 => "10100001",9381 => "00010001",9382 => "11011011",9383 => "11010001",9384 => "00111001",9385 => "10101000",9386 => "00000110",9387 => "10100101",9388 => "00101011",9389 => "11100001",9390 => "10001111",9391 => "10001000",9392 => "11110110",9393 => "00011100",9394 => "10100001",9395 => "00000110",9396 => "10110110",9397 => "01111110",9398 => "01001001",9399 => "01010000",9400 => "00010001",9401 => "01010010",9402 => "01101110",9403 => "00110010",9404 => "10011001",9405 => "01011011",9406 => "11100011",9407 => "01111010",9408 => "11010101",9409 => "11001100",9410 => "00111000",9411 => "11111100",9412 => "11011101",9413 => "11011100",9414 => "10001001",9415 => "11000110",9416 => "11100101",9417 => "01010100",9418 => "00010110",9419 => "10111100",9420 => "11111010",9421 => "10011001",9422 => "01011011",9423 => "00111100",9424 => "10111010",9425 => "10101111",9426 => "10100101",9427 => "01100110",9428 => "01101111",9429 => "00110110",9430 => "00100000",9431 => "11100110",9432 => "10101010",9433 => "11110010",9434 => "00000010",9435 => "01111001",9436 => "10001110",9437 => "11110000",9438 => "10010110",9439 => "00111000",9440 => "10010010",9441 => "01111101",9442 => "00100011",9443 => "11110100",9444 => "01100000",9445 => "00101011",9446 => "01111010",9447 => "10111001",9448 => "11000101",9449 => "11110001",9450 => "00000000",9451 => "10000001",9452 => "10010111",9453 => "11010110",9454 => "01011010",9455 => "01011010",9456 => "01011011",9457 => "10010110",9458 => "10011011",9459 => "11010010",9460 => "11000001",9461 => "11000101",9462 => "00011010",9463 => "01111111",9464 => "01111110",9465 => "10100110",9466 => "11110100",9467 => "00000101",9468 => "10101110",9469 => "10110100",9470 => "10011001",9471 => "10111011",9472 => "00011010",9473 => "01100001",9474 => "01110001",9475 => "10010000",9476 => "01111110",9477 => "01111001",9478 => "11110110",9479 => "11011011",9480 => "00100010",9481 => "00000001",9482 => "00001010",9483 => "11000101",9484 => "10110010",9485 => "11110000",9486 => "10000100",9487 => "01001011",9488 => "00101000",9489 => "00010110",9490 => "10001100",9491 => "10001100",9492 => "10011101",9493 => "00010101",9494 => "11011111",9495 => "11101001",9496 => "10010110",9497 => "01011010",9498 => "01010001",9499 => "11100011",9500 => "11001001",9501 => "10100000",9502 => "01101100",9503 => "01000110",9504 => "11010011",9505 => "01110101",9506 => "01011100",9507 => "01000001",9508 => "10010110",9509 => "11000000",9510 => "00011101",9511 => "00001011",9512 => "11100110",9513 => "11000110",9514 => "01011110",9515 => "00111011",9516 => "00001101",9517 => "00100111",9518 => "01000100",9519 => "00011111",9520 => "01111111",9521 => "11110101",9522 => "00000100",9523 => "00111110",9524 => "10111000",9525 => "11010101",9526 => "11001100",9527 => "01111011",9528 => "00101001",9529 => "10000010",9530 => "00110010",9531 => "11111010",9532 => "01011111",9533 => "01101011",9534 => "11001011",9535 => "11101100",9536 => "01011100",9537 => "00011000",9538 => "01101001",9539 => "10110111",9540 => "01000100",9541 => "00100000",9542 => "11001010",9543 => "10011111",9544 => "11001011",9545 => "00110101",9546 => "00110100",9547 => "01110001",9548 => "10001101",9549 => "10110011",9550 => "10111010",9551 => "11101111",9552 => "00011011",9553 => "11111000",9554 => "10011011",9555 => "10111001",9556 => "01000000",9557 => "11101101",9558 => "01111000",9559 => "10001010",9560 => "00110100",9561 => "01111110",9562 => "10101100",9563 => "00010000",9564 => "10001100",9565 => "00000100",9566 => "00010100",9567 => "00001111",9568 => "10111101",9569 => "00110101",9570 => "01100101",9571 => "00010100",9572 => "11111000",9573 => "10010010",9574 => "11111101",9575 => "10011101",9576 => "10001000",9577 => "01001001",9578 => "10011011",9579 => "11001010",9580 => "10100000",9581 => "11000101",9582 => "00011010",9583 => "11111101",9584 => "00110101",9585 => "01101110",9586 => "00111101",9587 => "00111000",9588 => "01111101",9589 => "01100001",9590 => "10100000",9591 => "00110101",9592 => "01010000",9593 => "01001111",9594 => "01011101",9595 => "01111100",9596 => "01011110",9597 => "10001011",9598 => "10010111",9599 => "01100111",9600 => "10101000",9601 => "00000100",9602 => "01111100",9603 => "10100001",9604 => "01011000",9605 => "11101011",9606 => "01011100",9607 => "10001011",9608 => "10001010",9609 => "10110111",9610 => "01110010",9611 => "11001111",9612 => "10010111",9613 => "11011110",9614 => "01000101",9615 => "10110110",9616 => "10001010",9617 => "00000000",9618 => "01111111",9619 => "00001111",9620 => "00001010",9621 => "10110110",9622 => "01110100",9623 => "10010100",9624 => "01001000",9625 => "11100001",9626 => "11111111",9627 => "11000010",9628 => "11111110",9629 => "10101110",9630 => "11010110",9631 => "10010010",9632 => "11101111",9633 => "01110100",9634 => "11101110",9635 => "00010010",9636 => "01111010",9637 => "00100010",9638 => "01001001",9639 => "00101001",9640 => "10000111",9641 => "00100111",9642 => "00000000",9643 => "01101101",9644 => "00100100",9645 => "00101100",9646 => "11100010",9647 => "10011111",9648 => "00110011",9649 => "01000000",9650 => "00111001",9651 => "10011110",9652 => "10110111",9653 => "10100000",9654 => "00010011",9655 => "00000011",9656 => "11010111",9657 => "01011111",9658 => "01010000",9659 => "01100010",9660 => "00110100",9661 => "11111000",9662 => "01000001",9663 => "10100111",9664 => "00010010",9665 => "11111000",9666 => "11011100",9667 => "11101111",9668 => "01111100",9669 => "01001101",9670 => "10100011",9671 => "10010010",9672 => "00011110",9673 => "10011000",9674 => "10011010",9675 => "01000011",9676 => "10011110",9677 => "10100101",9678 => "00000000",9679 => "11010110",9680 => "01010001",9681 => "00011101",9682 => "11011010",9683 => "01011010",9684 => "11100011",9685 => "10001010",9686 => "11011011",9687 => "10100101",9688 => "10110011",9689 => "01011110",9690 => "00110100",9691 => "01010111",9692 => "00111110",9693 => "00010110",9694 => "10100001",9695 => "10100101",9696 => "11100010",9697 => "10101001",9698 => "10001111",9699 => "01111100",9700 => "11111111",9701 => "00010101",9702 => "10010110",9703 => "00110000",9704 => "11110110",9705 => "11101111",9706 => "00000100",9707 => "10111011",9708 => "01101111",9709 => "00110101",9710 => "11111000",9711 => "11100010",9712 => "01011111",9713 => "10111000",9714 => "10000100",9715 => "01101000",9716 => "00010100",9717 => "01011111",9718 => "01000110",9719 => "10010100",9720 => "01001000",9721 => "11100110",9722 => "00011011",9723 => "11001001",9724 => "10000010",9725 => "10100001",9726 => "00110000",9727 => "10000111",9728 => "10001110",9729 => "10010100",9730 => "01011110",9731 => "10011000",9732 => "10100000",9733 => "00010101",9734 => "00001100",9735 => "00001101",9736 => "10111001",9737 => "11010011",9738 => "10111111",9739 => "00000000",9740 => "11110011",9741 => "11010100",9742 => "11010001",9743 => "00001011",9744 => "11010111",9745 => "10001111",9746 => "11111010",9747 => "11010100",9748 => "01001001",9749 => "10110100",9750 => "00100100",9751 => "11010010",9752 => "11101100",9753 => "10110100",9754 => "10001001",9755 => "10101111",9756 => "01101001",9757 => "01110001",9758 => "01101101",9759 => "10110111",9760 => "00111111",9761 => "00101110",9762 => "01011100",9763 => "00010101",9764 => "11101011",9765 => "11010110",9766 => "00010110",9767 => "00011100",9768 => "11111010",9769 => "10011001",9770 => "01111011",9771 => "00011001",9772 => "10000010",9773 => "00111110",9774 => "00110001",9775 => "11101001",9776 => "11110101",9777 => "00111100",9778 => "00110110",9779 => "01001111",9780 => "01001111",9781 => "00111001",9782 => "01000111",9783 => "01111100",9784 => "10111101",9785 => "11010011",9786 => "01000110",9787 => "01111100",9788 => "01100111",9789 => "11000011",9790 => "01100111",9791 => "11001110",9792 => "11010110",9793 => "10000011",9794 => "00101001",9795 => "00001101",9796 => "11000000",9797 => "01011111",9798 => "00110101",9799 => "01101000",9800 => "01101111",9801 => "00111111",9802 => "01001010",9803 => "00011101",9804 => "00110000",9805 => "11111000",9806 => "00111011",9807 => "10101001",9808 => "11100011",9809 => "00011101",9810 => "01101000",9811 => "00011110",9812 => "10110101",9813 => "01101001",9814 => "10000110",9815 => "00110101",9816 => "10111001",9817 => "01101111",9818 => "01011011",9819 => "00010111",9820 => "11111111",9821 => "11101100",9822 => "10000000",9823 => "01110110",9824 => "00101010",9825 => "10111000",9826 => "01000001",9827 => "01100000",9828 => "11100111",9829 => "11100100",9830 => "01111001",9831 => "00110101",9832 => "11110000",9833 => "01001111",9834 => "00110000",9835 => "10111000",9836 => "00000111",9837 => "01010100",9838 => "00101010",9839 => "00111111",9840 => "10011000",9841 => "00000011",9842 => "00110001",9843 => "00010001",9844 => "10110010",9845 => "10110010",9846 => "11101110",9847 => "00111010",9848 => "11110000",9849 => "11101011",9850 => "11000010",9851 => "11001010",9852 => "00111110",9853 => "01000000",9854 => "11010000",9855 => "10101011",9856 => "00000000",9857 => "00011000",9858 => "11111110",9859 => "01111110",9860 => "01011100",9861 => "11110101",9862 => "01010001",9863 => "01011010",9864 => "01111011",9865 => "00110000",9866 => "01110110",9867 => "10110011",9868 => "00000111",9869 => "00101110",9870 => "11000001",9871 => "00110000",9872 => "10001000",9873 => "01000110",9874 => "01010101",9875 => "01000000",9876 => "11101010",9877 => "00010010",9878 => "10100101",9879 => "00101001",9880 => "11110110",9881 => "10010010",9882 => "10000010",9883 => "11011001",9884 => "10011101",9885 => "01111001",9886 => "11100000",9887 => "10101101",9888 => "11011001",9889 => "01101011",9890 => "11010001",9891 => "00101011",9892 => "11011001",9893 => "11111000",9894 => "11110011",9895 => "01010100",9896 => "11001001",9897 => "11000011",9898 => "11010100",9899 => "10011011",9900 => "00101101",9901 => "01110111",9902 => "10111100",9903 => "01010100",9904 => "00101110",9905 => "10000001",9906 => "01011000",9907 => "00011101",9908 => "10101100",9909 => "00011011",9910 => "01101000",9911 => "10111011",9912 => "10101000",9913 => "01101000",9914 => "10000100",9915 => "11010110",9916 => "00010100",9917 => "00000010",9918 => "01000011",9919 => "11010111",9920 => "01010001",9921 => "01000101",9922 => "11100010",9923 => "00000011",9924 => "11001100",9925 => "10011011",9926 => "01110101",9927 => "00111001",9928 => "01110101",9929 => "01110101",9930 => "10001011",9931 => "00000101",9932 => "11011101",9933 => "01001000",9934 => "10000101",9935 => "00010000",9936 => "01001100",9937 => "01101010",9938 => "00000011",9939 => "10000101",9940 => "11010101",9941 => "10111011",9942 => "00011011",9943 => "10010011",9944 => "01110101",9945 => "10000110",9946 => "11100001",9947 => "00111000",9948 => "01000110",9949 => "11101011",9950 => "01111010",9951 => "00101101",9952 => "01101000",9953 => "01101100",9954 => "00100010",9955 => "10110010",9956 => "10000111",9957 => "00011101",9958 => "11100010",9959 => "00000101",9960 => "01000111",9961 => "11110000",9962 => "10010101",9963 => "11110001",9964 => "01011001",9965 => "11010101",9966 => "10100110",9967 => "11000101",9968 => "11000011",9969 => "01110101",9970 => "11100111",9971 => "01000000",9972 => "10010011",9973 => "11101101",9974 => "10000010",9975 => "10100101",9976 => "11111100",9977 => "10011100",9978 => "10110000",9979 => "10110101",9980 => "11010100",9981 => "10011111",9982 => "01101111",9983 => "11000011",9984 => "11000110",9985 => "00110100",9986 => "11111110",9987 => "11001110",9988 => "10011110",9989 => "10011001",9990 => "01000101",9991 => "00011010",9992 => "10100011",9993 => "00000101",9994 => "11000001",9995 => "01111010",9996 => "00101000",9997 => "10010110",9998 => "00101100",9999 => "00100011",10000 => "11101100",10001 => "00010110",10002 => "01100010",10003 => "11111010",10004 => "00010011",10005 => "11011101",10006 => "10001100",10007 => "11010111",10008 => "11001011",10009 => "01101110",10010 => "10010001",10011 => "11100001",10012 => "01111000",10013 => "10111111",10014 => "01111011",10015 => "11111001",10016 => "00101010",10017 => "00001001",10018 => "00101000",10019 => "10111001",10020 => "01110110",10021 => "10011010",10022 => "10011101",10023 => "01111110",10024 => "01101011",10025 => "11100100",10026 => "11011101",10027 => "01110000",10028 => "10111101",10029 => "11010111",10030 => "10101101",10031 => "00001110",10032 => "00111111",10033 => "11110000",10034 => "00010110",10035 => "00001011",10036 => "10110110",10037 => "10001111",10038 => "11001001",10039 => "01001010",10040 => "00101101",10041 => "11001001",10042 => "10110001",10043 => "11000100",10044 => "10000100",10045 => "00111111",10046 => "11101001",10047 => "11101011",10048 => "00011110",10049 => "00111000",10050 => "01110101",10051 => "01000010",10052 => "01001000",10053 => "01010110",10054 => "10001101",10055 => "10000000",10056 => "00010000",10057 => "00100001",10058 => "11000000",10059 => "01001110",10060 => "01110010",10061 => "00000010",10062 => "00000101",10063 => "01110100",10064 => "11101101",10065 => "01111000",10066 => "11000011",10067 => "00110110",10068 => "01101001",10069 => "11000010",10070 => "00000001",10071 => "11001010",10072 => "10110001",10073 => "01110110",10074 => "11100110",10075 => "00001100",10076 => "11010100",10077 => "10101110",10078 => "00100011",10079 => "01111110",10080 => "00111100",10081 => "01110011",10082 => "00111010",10083 => "11111001",10084 => "11110011",10085 => "10101100",10086 => "01110110",10087 => "01010001",10088 => "10101010",10089 => "00101000",10090 => "11001001",10091 => "01110101",10092 => "00000110",10093 => "10110000",10094 => "10111011",10095 => "11010100",10096 => "10100001",10097 => "01111111",10098 => "01101001",10099 => "00110111",10100 => "10011111",10101 => "00000010",10102 => "01111010",10103 => "11101010",10104 => "01110011",10105 => "01101000",10106 => "11000110",10107 => "00111000",10108 => "01010010",10109 => "10101111",10110 => "01001001",10111 => "10100101",10112 => "00100000",10113 => "11000000",10114 => "10110010",10115 => "10001101",10116 => "10011001",10117 => "01100100",10118 => "10110011",10119 => "10001100",10120 => "11000000",10121 => "11100001",10122 => "00010110",10123 => "10011011",10124 => "10001010",10125 => "00011001",10126 => "00100010",10127 => "00111000",10128 => "10001110",10129 => "01111111",10130 => "00111010",10131 => "00111011",10132 => "10111110",10133 => "10011001",10134 => "11111100",10135 => "00011101",10136 => "11010010",10137 => "10101111",10138 => "10111011",10139 => "00101011",10140 => "00000001",10141 => "00000001",10142 => "11011010",10143 => "01100010",10144 => "01101000",10145 => "01000111",10146 => "10011011",10147 => "11110111",10148 => "00011110",10149 => "11010110",10150 => "01001011",10151 => "10000010",10152 => "11010000",10153 => "01111100",10154 => "01110101",10155 => "01011011",10156 => "11101010",10157 => "11010110",10158 => "11110001",10159 => "10110110",10160 => "00011011",10161 => "10000001",10162 => "01000000",10163 => "00110010",10164 => "01110010",10165 => "10010001",10166 => "10111010",10167 => "01111100",10168 => "01100000",10169 => "11111001",10170 => "01000010",10171 => "10011001",10172 => "00000100",10173 => "01000000",10174 => "00001100",10175 => "00011011",10176 => "00110100",10177 => "11101011",10178 => "01000100",10179 => "01111010",10180 => "11011111",10181 => "10010110",10182 => "00010001",10183 => "10001100",10184 => "11111010",10185 => "01001000",10186 => "10101000",10187 => "00110001",10188 => "01101100",10189 => "11110000",10190 => "10111001",10191 => "11000110",10192 => "11101110",10193 => "01101010",10194 => "00101010",10195 => "11111110",10196 => "10111111",10197 => "00001110",10198 => "01000010",10199 => "10101110",10200 => "10110100",10201 => "01111111",10202 => "01011101",10203 => "01010100",10204 => "10101001",10205 => "01101101",10206 => "00000001",10207 => "01101111",10208 => "10001110",10209 => "00100100",10210 => "10100010",10211 => "10001000",10212 => "01011010",10213 => "01011101",10214 => "10111001",10215 => "01110000",10216 => "11111010",10217 => "00101110",10218 => "10000001",10219 => "10100110",10220 => "10001011",10221 => "00101001",10222 => "00101111",10223 => "11100111",10224 => "11111010",10225 => "00000110",10226 => "10100000",10227 => "11110100",10228 => "10011001",10229 => "11111011",10230 => "01111100",10231 => "01111000",10232 => "10110111",10233 => "01010111",10234 => "11011110",10235 => "11001110",10236 => "11100110",10237 => "11100000",10238 => "00010011",10239 => "11011010",10240 => "10100010",10241 => "01100011",10242 => "01000100",10243 => "01000100",10244 => "11011100",10245 => "00001111",10246 => "11010111",10247 => "10111011",10248 => "00000111",10249 => "11001010",10250 => "11100111",10251 => "10100000",10252 => "01011011",10253 => "10100110",10254 => "11001101",10255 => "10000100",10256 => "10101011",10257 => "01000101",10258 => "10001100",10259 => "10011010",10260 => "10010000",10261 => "01000110",10262 => "11011010",10263 => "11100001",10264 => "00001110",10265 => "10010011",10266 => "00001000",10267 => "01001110",10268 => "11111011",10269 => "01001010",10270 => "10111010",10271 => "00010101",10272 => "01111101",10273 => "01110111",10274 => "01011000",10275 => "00110100",10276 => "01000010",10277 => "10000000",10278 => "10001000",10279 => "01111100",10280 => "01011010",10281 => "11001010",10282 => "00111101",10283 => "00100110",10284 => "00101001",10285 => "11101111",10286 => "00111000",10287 => "01000001",10288 => "01101001",10289 => "10100100",10290 => "00111111",10291 => "11010000",10292 => "01011000",10293 => "11001100",10294 => "10011110",10295 => "11110101",10296 => "10110101",10297 => "00101111",10298 => "01110000",10299 => "00111110",10300 => "10011010",10301 => "00100001",10302 => "10100001",10303 => "00000000",10304 => "10110000",10305 => "10001000",10306 => "10100100",10307 => "00100100",10308 => "00111001",10309 => "10001100",10310 => "10111010",10311 => "10110010",10312 => "11010001",10313 => "11001000",10314 => "00000100",10315 => "01100001",10316 => "00110000",10317 => "11111011",10318 => "00010101",10319 => "11010111",10320 => "01100101",10321 => "11011111",10322 => "01100010",10323 => "10101110",10324 => "10011011",10325 => "01110111",10326 => "10001000",10327 => "11101100",10328 => "00111110",10329 => "01111000",10330 => "10111110",10331 => "01110100",10332 => "11111010",10333 => "10011011",10334 => "10010011",10335 => "11101100",10336 => "10001000",10337 => "10100011",10338 => "00011100",10339 => "11000000",10340 => "00001101",10341 => "00101000",10342 => "00000110",10343 => "00000011",10344 => "11000001",10345 => "11000100",10346 => "11011100",10347 => "00110000",10348 => "10000001",10349 => "00111110",10350 => "01101000",10351 => "10101001",10352 => "10100001",10353 => "11000111",10354 => "00110000",10355 => "01010011",10356 => "00011110",10357 => "11010101",10358 => "01111101",10359 => "11100010",10360 => "11110000",10361 => "11111111",10362 => "11000100",10363 => "01110110",10364 => "11010100",10365 => "00001001",10366 => "00001110",10367 => "00110001",10368 => "10100010",10369 => "00011110",10370 => "01000110",10371 => "11010001",10372 => "01001000",10373 => "11110101",10374 => "01111101",10375 => "10001011",10376 => "01101000",10377 => "00100111",10378 => "00001001",10379 => "10110000",10380 => "00101001",10381 => "00111001",10382 => "00101001",10383 => "10010101",10384 => "11000111",10385 => "10110111",10386 => "01011001",10387 => "11111011",10388 => "11111000",10389 => "10111011",10390 => "11110001",10391 => "01100011",10392 => "01100000",10393 => "11110101",10394 => "11010011",10395 => "01001101",10396 => "01110001",10397 => "10100100",10398 => "11101101",10399 => "11110011",10400 => "00010011",10401 => "10111001",10402 => "11111111",10403 => "11000101",10404 => "11000111",10405 => "11111101",10406 => "00011010",10407 => "10011000",10408 => "00000010",10409 => "01010011",10410 => "10000001",10411 => "01011101",10412 => "01110010",10413 => "00011110",10414 => "10010001",10415 => "11110110",10416 => "10110100",10417 => "11001000",10418 => "01010000",10419 => "00111010",10420 => "01110010",10421 => "00011100",10422 => "00111100",10423 => "10011010",10424 => "10000010",10425 => "10100100",10426 => "11010101",10427 => "11100110",10428 => "01010011",10429 => "01001110",10430 => "00001010",10431 => "10111000",10432 => "01101111",10433 => "11111111",10434 => "11100011",10435 => "10001010",10436 => "11111011",10437 => "00101110",10438 => "00000101",10439 => "10101101",10440 => "10110101",10441 => "01010101",10442 => "10001100",10443 => "11101110",10444 => "11011111",10445 => "11100011",10446 => "11000110",10447 => "01010001",10448 => "10111001",10449 => "01110110",10450 => "00110011",10451 => "00110001",10452 => "10111010",10453 => "00001111",10454 => "11100010",10455 => "10010011",10456 => "00100011",10457 => "10100010",10458 => "00111101",10459 => "01100110",10460 => "10110011",10461 => "00111110",10462 => "11100011",10463 => "10101001",10464 => "00000111",10465 => "10110000",10466 => "10011001",10467 => "00110110",10468 => "00000100",10469 => "10010101",10470 => "00001010",10471 => "11001011",10472 => "01001010",10473 => "11111011",10474 => "01111001",10475 => "01011010",10476 => "10101111",10477 => "01110010",10478 => "10100010",10479 => "00000001",10480 => "11101001",10481 => "10100100",10482 => "01111010",10483 => "10111001",10484 => "00001110",10485 => "01100000",10486 => "00101100",10487 => "11011100",10488 => "10001010",10489 => "11010001",10490 => "00000101",10491 => "10111011",10492 => "11100001",10493 => "00100000",10494 => "00100110",10495 => "10001010",10496 => "00100011",10497 => "00100100",10498 => "10100111",10499 => "10101100",10500 => "10000011",10501 => "11110101",10502 => "10010111",10503 => "01100010",10504 => "01000001",10505 => "01101101",10506 => "01100100",10507 => "00101010",10508 => "01101100",10509 => "11111101",10510 => "00000111",10511 => "01011101",10512 => "11010110",10513 => "10100111",10514 => "10101111",10515 => "00001001",10516 => "01100101",10517 => "01000011",10518 => "11101010",10519 => "00001110",10520 => "01001000",10521 => "01100100",10522 => "10010101",10523 => "10010110",10524 => "10011100",10525 => "10110111",10526 => "01101101",10527 => "01000110",10528 => "01111110",10529 => "11111110",10530 => "01001111",10531 => "11110011",10532 => "10111000",10533 => "10001001",10534 => "00110110",10535 => "01111001",10536 => "01111000",10537 => "11100001",10538 => "00001010",10539 => "01101000",10540 => "10000010",10541 => "11100101",10542 => "01110110",10543 => "11111101",10544 => "10011111",10545 => "10101101",10546 => "00010010",10547 => "11000100",10548 => "10001010",10549 => "00101110",10550 => "01011111",10551 => "01111111",10552 => "01010011",10553 => "00011011",10554 => "00010110",10555 => "00011000",10556 => "10010111",10557 => "01001100",10558 => "11011011",10559 => "01010010",10560 => "01110000",10561 => "10011101",10562 => "10110011",10563 => "00100001",10564 => "11111001",10565 => "01010110",10566 => "11110100",10567 => "11101110",10568 => "01010000",10569 => "00001100",10570 => "01110010",10571 => "11110010",10572 => "00110001",10573 => "01010110",10574 => "10001000",10575 => "00010000",10576 => "00110110",10577 => "11111111",10578 => "11011000",10579 => "11010111",10580 => "11111000",10581 => "11001101",10582 => "11110111",10583 => "00010010",10584 => "00001010",10585 => "11001000",10586 => "00010100",10587 => "00011011",10588 => "01101111",10589 => "01110011",10590 => "11001111",10591 => "00011011",10592 => "10000110",10593 => "01011110",10594 => "10101110",10595 => "11011100",10596 => "11100100",10597 => "00101001",10598 => "01101001",10599 => "00010111",10600 => "11001101",10601 => "00010001",10602 => "11010011",10603 => "10101001",10604 => "00111010",10605 => "01011101",10606 => "11100101",10607 => "00001111",10608 => "10000010",10609 => "01000100",10610 => "01110011",10611 => "01100010",10612 => "00000111",10613 => "10111111",10614 => "00000010",10615 => "11111000",10616 => "01000000",10617 => "11111011",10618 => "00111001",10619 => "11111100",10620 => "01011100",10621 => "00110100",10622 => "01011111",10623 => "10011001",10624 => "10010111",10625 => "10001010",10626 => "11110001",10627 => "11011010",10628 => "01100100",10629 => "11101001",10630 => "10111000",10631 => "11000110",10632 => "00100101",10633 => "11011101",10634 => "10000100",10635 => "10000000",10636 => "01010110",10637 => "00000110",10638 => "10000011",10639 => "00011001",10640 => "01001110",10641 => "00000110",10642 => "11111011",10643 => "10000010",10644 => "00100000",10645 => "01101001",10646 => "01110000",10647 => "01111100",10648 => "10011111",10649 => "00100010",10650 => "10111000",10651 => "10101100",10652 => "01111011",10653 => "11010101",10654 => "00010110",10655 => "11100010",10656 => "10100111",10657 => "00101001",10658 => "01001001",10659 => "11111011",10660 => "01010000",10661 => "01101100",10662 => "00000001",10663 => "00010101",10664 => "10000000",10665 => "11100101",10666 => "00100111",10667 => "11100101",10668 => "00011000",10669 => "01111110",10670 => "11011011",10671 => "00011100",10672 => "11100100",10673 => "10010011",10674 => "00001011",10675 => "01111000",10676 => "11000000",10677 => "11101100",10678 => "00011001",10679 => "10011000",10680 => "10101100",10681 => "11111011",10682 => "00001100",10683 => "01110110",10684 => "01011000",10685 => "11101000",10686 => "10101110",10687 => "01111111",10688 => "01111110",10689 => "01111000",10690 => "00011100",10691 => "11110011",10692 => "10110001",10693 => "01011100",10694 => "01010000",10695 => "00110110",10696 => "00110010",10697 => "10001100",10698 => "00000110",10699 => "00011111",10700 => "01001110",10701 => "01000101",10702 => "10111001",10703 => "01100110",10704 => "11101100",10705 => "11111001",10706 => "00001100",10707 => "10001001",10708 => "10100011",10709 => "00010110",10710 => "10000000",10711 => "10001011",10712 => "11011000",10713 => "00110110",10714 => "11100111",10715 => "00101000",10716 => "00000010",10717 => "00100100",10718 => "01100101",10719 => "11111011",10720 => "01101010",10721 => "10001001",10722 => "11111000",10723 => "10101110",10724 => "10001111",10725 => "11100001",10726 => "00110110",10727 => "01101010",10728 => "10111100",10729 => "10110100",10730 => "11100001",10731 => "10101011",10732 => "00101000",10733 => "01000000",10734 => "01111011",10735 => "10000011",10736 => "10000100",10737 => "10100010",10738 => "01000001",10739 => "01100101",10740 => "11000000",10741 => "01001001",10742 => "11101010",10743 => "10100000",10744 => "11100100",10745 => "00001001",10746 => "11100001",10747 => "11110000",10748 => "10010001",10749 => "00001101",10750 => "00100000",10751 => "11001110",10752 => "10010100",10753 => "00001111",10754 => "01001101",10755 => "11110001",10756 => "00110001",10757 => "00011110",10758 => "00000110",10759 => "11101111",10760 => "01001010",10761 => "01010111",10762 => "11100000",10763 => "11100101",10764 => "01101010",10765 => "01100001",10766 => "10100010",10767 => "11011000",10768 => "00001001",10769 => "01101111",10770 => "00000010",10771 => "01011101",10772 => "00001100",10773 => "00010011",10774 => "00011100",10775 => "11000101",10776 => "01101011",10777 => "11110110",10778 => "00110110",10779 => "10000000",10780 => "11000001",10781 => "10111010",10782 => "00111001",10783 => "11101001",10784 => "00011010",10785 => "10000001",10786 => "11001010",10787 => "11111111",10788 => "00011000",10789 => "10110100",10790 => "00110001",10791 => "01011101",10792 => "00001011",10793 => "11010011",10794 => "01110011",10795 => "10000001",10796 => "11011010",10797 => "00101010",10798 => "01110001",10799 => "00010001",10800 => "10010111",10801 => "11010000",10802 => "10011001",10803 => "10111000",10804 => "01010110",10805 => "11100001",10806 => "11000110",10807 => "00000011",10808 => "00010101",10809 => "11010100",10810 => "11000011",10811 => "10011110",10812 => "11101101",10813 => "10101101",10814 => "01111000",10815 => "00001001",10816 => "10010110",10817 => "11111111",10818 => "10100111",10819 => "01001011",10820 => "00111110",10821 => "11110101",10822 => "00101001",10823 => "01101000",10824 => "10001110",10825 => "00100101",10826 => "00000101",10827 => "01101110",10828 => "00000011",10829 => "01110110",10830 => "01000110",10831 => "11001000",10832 => "10000101",10833 => "10001000",10834 => "01011011",10835 => "10010100",10836 => "10101100",10837 => "11100111",10838 => "01110101",10839 => "10111100",10840 => "10101010",10841 => "00100000",10842 => "01010110",10843 => "10001100",10844 => "11000101",10845 => "11101111",10846 => "01001111",10847 => "10000000",10848 => "00011000",10849 => "00010001",10850 => "11111000",10851 => "11010000",10852 => "01111110",10853 => "00110011",10854 => "00111111",10855 => "01101101",10856 => "11110000",10857 => "11010101",10858 => "10010001",10859 => "11110010",10860 => "00000001",10861 => "00010101",10862 => "11100011",10863 => "10001011",10864 => "00100110",10865 => "00011110",10866 => "01011100",10867 => "01001111",10868 => "10001011",10869 => "11001100",10870 => "10101001",10871 => "11110100",10872 => "10100110",10873 => "00011001",10874 => "10011110",10875 => "10011100",10876 => "01100110",10877 => "11011111",10878 => "01100111",10879 => "10100011",10880 => "00001100",10881 => "11000001",10882 => "11100100",10883 => "00011010",10884 => "11011111",10885 => "10111000",10886 => "10000011",10887 => "01010000",10888 => "00000010",10889 => "00100000",10890 => "00110100",10891 => "01001011",10892 => "11110100",10893 => "01000010",10894 => "00010010",10895 => "10011010",10896 => "01001000",10897 => "00001000",10898 => "11010111",10899 => "00001101",10900 => "11001010",10901 => "11101001",10902 => "00111100",10903 => "11111111",10904 => "11101110",10905 => "00001111",10906 => "11000001",10907 => "01100001",10908 => "11100110",10909 => "01011110",10910 => "10111001",10911 => "11011101",10912 => "00010011",10913 => "00010000",10914 => "00100110",10915 => "00100110",10916 => "00111001",10917 => "11111011",10918 => "11101101",10919 => "00110110",10920 => "01000110",10921 => "00010011",10922 => "11011010",10923 => "11110000",10924 => "10110100",10925 => "01000011",10926 => "11001101",10927 => "11100100",10928 => "11110001",10929 => "00000011",10930 => "11110110",10931 => "10101100",10932 => "01001111",10933 => "00101100",10934 => "00111000",10935 => "01001110",10936 => "01010011",10937 => "11101011",10938 => "00000111",10939 => "00100001",10940 => "11011100",10941 => "10001011",10942 => "01100101",10943 => "11110110",10944 => "00100011",10945 => "01010111",10946 => "01001000",10947 => "10001101",10948 => "01010010",10949 => "00100001",10950 => "01011000",10951 => "11000110",10952 => "11111101",10953 => "11011111",10954 => "00010000",10955 => "01011010",10956 => "01010011",10957 => "11011100",10958 => "01010110",10959 => "01010000",10960 => "01000110",10961 => "10111111",10962 => "11110111",10963 => "11010101",10964 => "10100010",10965 => "00000101",10966 => "01101101",10967 => "11100000",10968 => "11100110",10969 => "01110010",10970 => "10111111",10971 => "10011011",10972 => "00000110",10973 => "10111000",10974 => "11001011",10975 => "00010100",10976 => "01011001",10977 => "11101101",10978 => "01100100",10979 => "01010100",10980 => "10011111",10981 => "00110011",10982 => "01000111",10983 => "11100110",10984 => "11010100",10985 => "00011111",10986 => "11001100",10987 => "10011010",10988 => "10100110",10989 => "00111001",10990 => "01110101",10991 => "11110110",10992 => "01010001",10993 => "01001000",10994 => "00100101",10995 => "00100100",10996 => "11011100",10997 => "10110000",10998 => "00001001",10999 => "10110100",11000 => "11111100",11001 => "00100110",11002 => "11111110",11003 => "00011000",11004 => "11101000",11005 => "10011001",11006 => "11000110",11007 => "10110010",11008 => "00010111",11009 => "11101111",11010 => "11100010",11011 => "10100011",11012 => "11100011",11013 => "10010111",11014 => "11111100",11015 => "11111101",11016 => "00010001",11017 => "10111110",11018 => "11011111",11019 => "01110000",11020 => "10111011",11021 => "11000111",11022 => "11101111",11023 => "10011100",11024 => "01100010",11025 => "01011001",11026 => "01100001",11027 => "01111110",11028 => "00101111",11029 => "00010000",11030 => "00011100",11031 => "10111000",11032 => "00001000",11033 => "10111101",11034 => "01110010",11035 => "01000110",11036 => "11101000",11037 => "10001011",11038 => "10011001",11039 => "00011110",11040 => "01111100",11041 => "10111000",11042 => "11010001",11043 => "01101100",11044 => "10111001",11045 => "11110111",11046 => "10000011",11047 => "01001000",11048 => "11101110",11049 => "11010101",11050 => "00111010",11051 => "11010010",11052 => "11000110",11053 => "01001000",11054 => "01011111",11055 => "11111101",11056 => "00100111",11057 => "10100010",11058 => "11011011",11059 => "11101001",11060 => "11011000",11061 => "01100001",11062 => "01110101",11063 => "11001011",11064 => "01001110",11065 => "11011111",11066 => "01011001",11067 => "11001101",11068 => "11111111",11069 => "00111001",11070 => "00011111",11071 => "00001110",11072 => "00100101",11073 => "00010110",11074 => "10011010",11075 => "00000100",11076 => "11010110",11077 => "11001101",11078 => "11000001",11079 => "01110011",11080 => "10001100",11081 => "00000101",11082 => "10101110",11083 => "01000001",11084 => "11100110",11085 => "10010000",11086 => "10010000",11087 => "01101110",11088 => "00111001",11089 => "11101111",11090 => "01010100",11091 => "00000011",11092 => "01001111",11093 => "11110111",11094 => "00101010",11095 => "01010001",11096 => "10001010",11097 => "00000001",11098 => "00001101",11099 => "01010111",11100 => "01110101",11101 => "11000110",11102 => "01000101",11103 => "11110101",11104 => "11010110",11105 => "00001111",11106 => "10000001",11107 => "11111000",11108 => "11001101",11109 => "11111010",11110 => "00010100",11111 => "10010110",11112 => "10000100",11113 => "11001100",11114 => "10011010",11115 => "01101100",11116 => "00001110",11117 => "11110110",11118 => "00101001",11119 => "00011010",11120 => "11111011",11121 => "00111111",11122 => "00110111",11123 => "11001110",11124 => "11100000",11125 => "01011111",11126 => "10010010",11127 => "11010100",11128 => "00011011",11129 => "01010111",11130 => "01001010",11131 => "10010100",11132 => "00010101",11133 => "11011100",11134 => "01001011",11135 => "10001010",11136 => "00000101",11137 => "11101110",11138 => "10111011",11139 => "00110111",11140 => "01101011",11141 => "10110101",11142 => "01101110",11143 => "01100011",11144 => "11010100",11145 => "11000011",11146 => "11110111",11147 => "01101010",11148 => "11111001",11149 => "11011110",11150 => "11110000",11151 => "00000110",11152 => "11101101",11153 => "00110100",11154 => "10101111",11155 => "00000001",11156 => "00010000",11157 => "00100111",11158 => "01100111",11159 => "11011111",11160 => "00000100",11161 => "01010010",11162 => "10010111",11163 => "00011111",11164 => "11001100",11165 => "10000011",11166 => "00010101",11167 => "00110110",11168 => "10111011",11169 => "11010101",11170 => "10010000",11171 => "00110011",11172 => "01011111",11173 => "01110111",11174 => "01011101",11175 => "01110110",11176 => "11110000",11177 => "11001011",11178 => "00111111",11179 => "00001100",11180 => "10000111",11181 => "00000010",11182 => "00100000",11183 => "00101011",11184 => "01010110",11185 => "01001111",11186 => "10111001",11187 => "11011100",11188 => "01010011",11189 => "01000110",11190 => "11001101",11191 => "00010001",11192 => "01101100",11193 => "10000100",11194 => "01111101",11195 => "01101110",11196 => "00010000",11197 => "00010100",11198 => "01010000",11199 => "00101111",11200 => "10011110",11201 => "10011101",11202 => "00110101",11203 => "01111000",11204 => "00100111",11205 => "00100000",11206 => "10010101",11207 => "10010000",11208 => "00010110",11209 => "11010010",11210 => "10010001",11211 => "11010011",11212 => "10001100",11213 => "11010111",11214 => "11110001",11215 => "01011011",11216 => "10010100",11217 => "01010011",11218 => "11110001",11219 => "01001111",11220 => "11101100",11221 => "01111000",11222 => "11001110",11223 => "10110010",11224 => "11010100",11225 => "00001011",11226 => "00101110",11227 => "00000111",11228 => "00111010",11229 => "11011000",11230 => "01010111",11231 => "01100111",11232 => "11110001",11233 => "10110011",11234 => "10010011",11235 => "10000101",11236 => "01001011",11237 => "11001110",11238 => "00111001",11239 => "01110011",11240 => "00110010",11241 => "11001100",11242 => "01011010",11243 => "01001111",11244 => "00111001",11245 => "01000100",11246 => "11111111",11247 => "11010111",11248 => "10110010",11249 => "11000101",11250 => "00101010",11251 => "00101000",11252 => "01011111",11253 => "00110111",11254 => "11101101",11255 => "01001111",11256 => "00001011",11257 => "11111101",11258 => "01000110",11259 => "01111011",11260 => "00100110",11261 => "10110011",11262 => "00110011",11263 => "01001110",11264 => "01111110",11265 => "11100000",11266 => "10010010",11267 => "11101101",11268 => "11100101",11269 => "11000001",11270 => "10101001",11271 => "00001010",11272 => "10001101",11273 => "10101010",11274 => "11110000",11275 => "00000000",11276 => "10111110",11277 => "01011101",11278 => "01101101",11279 => "10001000",11280 => "10111000",11281 => "11001110",11282 => "01011000",11283 => "11110011",11284 => "01100111",11285 => "00111100",11286 => "10010100",11287 => "11011010",11288 => "00101111",11289 => "00010111",11290 => "11100101",11291 => "00001000",11292 => "01000111",11293 => "11010111",11294 => "11010000",11295 => "10000001",11296 => "10111001",11297 => "01110010",11298 => "00001011",11299 => "10001101",11300 => "00111001",11301 => "01110100",11302 => "00000101",11303 => "11101011",11304 => "00000001",11305 => "01001010",11306 => "00000011",11307 => "01011100",11308 => "10110001",11309 => "10100011",11310 => "10111000",11311 => "10011011",11312 => "00010001",11313 => "10000110",11314 => "11010000",11315 => "01010101",11316 => "10110010",11317 => "10101110",11318 => "11111011",11319 => "10110010",11320 => "11110011",11321 => "11011000",11322 => "00101100",11323 => "11011101",11324 => "00100010",11325 => "00100011",11326 => "00000110",11327 => "00111110",11328 => "10110110",11329 => "01010010",11330 => "00010110",11331 => "00010001",11332 => "01110110",11333 => "01001000",11334 => "00100110",11335 => "00101010",11336 => "01000101",11337 => "01101111",11338 => "11001111",11339 => "11011111",11340 => "01101001",11341 => "01100011",11342 => "10100101",11343 => "11000110",11344 => "00010110",11345 => "01010001",11346 => "01101001",11347 => "10101110",11348 => "11100001",11349 => "00010100",11350 => "01111101",11351 => "01000011",11352 => "00001101",11353 => "11100000",11354 => "00101000",11355 => "10001010",11356 => "01111011",11357 => "10100000",11358 => "01111101",11359 => "01110000",11360 => "10010010",11361 => "10100010",11362 => "01111101",11363 => "01001110",11364 => "11010010",11365 => "11111001",11366 => "00000100",11367 => "00011011",11368 => "10010101",11369 => "10001000",11370 => "00001011",11371 => "11111010",11372 => "10010000",11373 => "01011100",11374 => "10101110",11375 => "10110010",11376 => "11111010",11377 => "00101111",11378 => "11011001",11379 => "01111110",11380 => "10100100",11381 => "11101101",11382 => "10001101",11383 => "00110101",11384 => "01001001",11385 => "00011111",11386 => "00010000",11387 => "01011000",11388 => "11010101",11389 => "01101001",11390 => "10000001",11391 => "01001101",11392 => "10111100",11393 => "10010001",11394 => "01100101",11395 => "11110100",11396 => "00011101",11397 => "11111101",11398 => "01110010",11399 => "11101000",11400 => "10101111",11401 => "11011111",11402 => "11001110",11403 => "10001011",11404 => "00000100",11405 => "11011111",11406 => "10011101",11407 => "10011011",11408 => "00011011",11409 => "11110011",11410 => "11101011",11411 => "00011110",11412 => "10101000",11413 => "00101010",11414 => "00111011",11415 => "10011101",11416 => "11110001",11417 => "11000111",11418 => "01010011",11419 => "10011001",11420 => "01001111",11421 => "10001101",11422 => "01000001",11423 => "11001001",11424 => "00010001",11425 => "10010010",11426 => "11101001",11427 => "01011100",11428 => "11110000",11429 => "00101101",11430 => "10010001",11431 => "01000001",11432 => "11011010",11433 => "00001110",11434 => "10101100",11435 => "01101111",11436 => "01101000",11437 => "10101000",11438 => "10111011",11439 => "10111110",11440 => "00000000",11441 => "10100011",11442 => "01000000",11443 => "00100001",11444 => "11110001",11445 => "11100001",11446 => "01001000",11447 => "01000100",11448 => "01100000",11449 => "11100010",11450 => "00011110",11451 => "00000101",11452 => "10101010",11453 => "01101101",11454 => "00001111",11455 => "01010010",11456 => "01010001",11457 => "10010010",11458 => "01101001",11459 => "10111110",11460 => "01001110",11461 => "10011011",11462 => "00010001",11463 => "01001000",11464 => "10110100",11465 => "01010111",11466 => "10110000",11467 => "11101000",11468 => "01111001",11469 => "11111001",11470 => "10000000",11471 => "00110001",11472 => "00110010",11473 => "01001000",11474 => "10101100",11475 => "01111110",11476 => "00010111",11477 => "01011100",11478 => "01100101",11479 => "00100100",11480 => "10011100",11481 => "10000001",11482 => "11011000",11483 => "00011100",11484 => "01000111",11485 => "11111101",11486 => "11110010",11487 => "11001010",11488 => "11010011",11489 => "10100110",11490 => "10001100",11491 => "01010111",11492 => "11101011",11493 => "10101011",11494 => "10001100",11495 => "10100111",11496 => "10110110",11497 => "01010101",11498 => "01101010",11499 => "01111000",11500 => "10001010",11501 => "00100101",11502 => "01011110",11503 => "11000111",11504 => "11010111",11505 => "11110000",11506 => "01011100",11507 => "11101110",11508 => "11010010",11509 => "10110101",11510 => "11000110",11511 => "01110000",11512 => "10001111",11513 => "01011011",11514 => "11100010",11515 => "01110011",11516 => "01110000",11517 => "11010100",11518 => "10100111",11519 => "01000011",11520 => "11111011",11521 => "01101101",11522 => "00110111",11523 => "00111010",11524 => "01000011",11525 => "01000111",11526 => "11111111",11527 => "01111100",11528 => "01111010",11529 => "00110101",11530 => "01110111",11531 => "00100100",11532 => "11101010",11533 => "00010100",11534 => "11100000",11535 => "11001110",11536 => "11011011",11537 => "00100101",11538 => "11100011",11539 => "11110001",11540 => "11110100",11541 => "11101010",11542 => "00011010",11543 => "10111010",11544 => "11010101",11545 => "11011010",11546 => "01011100",11547 => "11011011",11548 => "11110001",11549 => "00001011",11550 => "10101011",11551 => "00100101",11552 => "01100110",11553 => "01001010",11554 => "10110101",11555 => "11100000",11556 => "11111101",11557 => "11101011",11558 => "11111101",11559 => "01001001",11560 => "01011010",11561 => "10010100",11562 => "10100111",11563 => "10011111",11564 => "01100010",11565 => "11011100",11566 => "10001110",11567 => "10111111",11568 => "01000000",11569 => "01000010",11570 => "11111110",11571 => "00011010",11572 => "10011011",11573 => "00101011",11574 => "00110100",11575 => "01000100",11576 => "00110011",11577 => "01100011",11578 => "01111010",11579 => "10101000",11580 => "01000001",11581 => "10111101",11582 => "11100101",11583 => "10101001",11584 => "00000001",11585 => "01011000",11586 => "10011100",11587 => "01011000",11588 => "00101001",11589 => "00010101",11590 => "01110100",11591 => "00010000",11592 => "11101001",11593 => "00100101",11594 => "00010001",11595 => "01110111",11596 => "10101001",11597 => "10011111",11598 => "01000000",11599 => "00001100",11600 => "00101111",11601 => "01000011",11602 => "11010011",11603 => "11001110",11604 => "01001101",11605 => "01111100",11606 => "00110111",11607 => "10001010",11608 => "11110101",11609 => "01001010",11610 => "01111011",11611 => "00000101",11612 => "11001111",11613 => "01011111",11614 => "01001000",11615 => "10101000",11616 => "11100000",11617 => "00011101",11618 => "10110011",11619 => "10100111",11620 => "00101111",11621 => "11010101",11622 => "11100111",11623 => "01110011",11624 => "01001000",11625 => "01111101",11626 => "00010100",11627 => "11100110",11628 => "10011001",11629 => "11110010",11630 => "00011111",11631 => "11001000",11632 => "01011100",11633 => "10100011",11634 => "10001001",11635 => "00010110",11636 => "00011011",11637 => "01110110",11638 => "11110100",11639 => "00100010",11640 => "10101100",11641 => "00011011",11642 => "11010110",11643 => "10111100",11644 => "11010111",11645 => "00001010",11646 => "10010001",11647 => "10111101",11648 => "11111100",11649 => "00010111",11650 => "11110001",11651 => "11000100",11652 => "00000011",11653 => "01111001",11654 => "10100101",11655 => "00101000",11656 => "11110100",11657 => "01000101",11658 => "11110010",11659 => "11011101",11660 => "11001011",11661 => "10001001",11662 => "10110000",11663 => "10100010",11664 => "00111101",11665 => "00010101",11666 => "11101100",11667 => "00100110",11668 => "10110011",11669 => "00011000",11670 => "01110011",11671 => "10000011",11672 => "01000101",11673 => "01001011",11674 => "01010100",11675 => "11111111",11676 => "00110010",11677 => "01101101",11678 => "00110110",11679 => "00001100",11680 => "01100001",11681 => "11000011",11682 => "10001110",11683 => "01000100",11684 => "10001100",11685 => "01101110",11686 => "01110000",11687 => "00011100",11688 => "00000000",11689 => "11110001",11690 => "10110010",11691 => "00001110",11692 => "00011010",11693 => "10100110",11694 => "10111010",11695 => "00001000",11696 => "10011001",11697 => "01011111",11698 => "11011101",11699 => "11111010",11700 => "00110011",11701 => "11001111",11702 => "01100010",11703 => "01010010",11704 => "00100001",11705 => "10011100",11706 => "00010000",11707 => "11000000",11708 => "01100001",11709 => "11111011",11710 => "11000000",11711 => "01110010",11712 => "01010100",11713 => "10110110",11714 => "01010111",11715 => "10110111",11716 => "00001010",11717 => "11011110",11718 => "00111001",11719 => "11001110",11720 => "01000010",11721 => "11100110",11722 => "10011011",11723 => "11101000",11724 => "01111011",11725 => "01111101",11726 => "00110011",11727 => "01001000",11728 => "10001110",11729 => "00001001",11730 => "00111010",11731 => "01101100",11732 => "11101101",11733 => "01010010",11734 => "10001101",11735 => "00110001",11736 => "11000001",11737 => "00010110",11738 => "11010101",11739 => "11100011",11740 => "01100101",11741 => "00110111",11742 => "11010000",11743 => "00011100",11744 => "10101100",11745 => "00010011",11746 => "11100110",11747 => "01100101",11748 => "01011101",11749 => "11001010",11750 => "01100110",11751 => "01101110",11752 => "10111011",11753 => "11001101",11754 => "01110000",11755 => "01000101",11756 => "01100100",11757 => "00101001",11758 => "11110010",11759 => "10000000",11760 => "01110000",11761 => "10010010",11762 => "11010000",11763 => "11011100",11764 => "00101000",11765 => "01111010",11766 => "11011111",11767 => "01110101",11768 => "10111101",11769 => "11111001",11770 => "01100100",11771 => "01101001",11772 => "10111111",11773 => "00100011",11774 => "10001000",11775 => "11011100",11776 => "01011111",11777 => "10001010",11778 => "00011100",11779 => "10000101",11780 => "01011010",11781 => "01010101",11782 => "10001011",11783 => "10011011",11784 => "01111001",11785 => "00110111",11786 => "10010110",11787 => "00011111",11788 => "11100001",11789 => "00111001",11790 => "10010010",11791 => "00100100",11792 => "11011101",11793 => "01100000",11794 => "01000011",11795 => "11000100",11796 => "11011100",11797 => "10000011",11798 => "00000110",11799 => "11100111",11800 => "11111000",11801 => "00001010",11802 => "01001000",11803 => "10001011",11804 => "11001001",11805 => "01101011",11806 => "01110010",11807 => "01110001",11808 => "11000011",11809 => "11100011",11810 => "11100100",11811 => "10111011",11812 => "11011100",11813 => "00110000",11814 => "11011011",11815 => "10000101",11816 => "11001101",11817 => "10100110",11818 => "11100100",11819 => "11001111",11820 => "11010111",11821 => "11110110",11822 => "01011101",11823 => "11001101",11824 => "00100000",11825 => "01011011",11826 => "00001001",11827 => "11110001",11828 => "00100110",11829 => "00010111",11830 => "11000111",11831 => "01111101",11832 => "00101000",11833 => "01100010",11834 => "01100000",11835 => "11011100",11836 => "10101010",11837 => "01000111",11838 => "11111000",11839 => "11100110",11840 => "11101100",11841 => "01010100",11842 => "11110111",11843 => "10000001",11844 => "01110010",11845 => "00011101",11846 => "10011000",11847 => "11001100",11848 => "11100010",11849 => "10000110",11850 => "10010010",11851 => "11110010",11852 => "01011100",11853 => "10100000",11854 => "01100001",11855 => "11011110",11856 => "11100111",11857 => "01101000",11858 => "00101111",11859 => "00101111",11860 => "11111011",11861 => "00101011",11862 => "11110011",11863 => "10110011",11864 => "10011100",11865 => "11001011",11866 => "10011011",11867 => "00000001",11868 => "10101000",11869 => "01100011",11870 => "01000010",11871 => "00011100",11872 => "00001010",11873 => "00001100",11874 => "10111110",11875 => "00111110",11876 => "10100010",11877 => "10110111",11878 => "01110001",11879 => "10110010",11880 => "00011010",11881 => "10011111",11882 => "01100001",11883 => "10111010",11884 => "11000000",11885 => "01000101",11886 => "01101011",11887 => "10011101",11888 => "01111010",11889 => "00011111",11890 => "00000110",11891 => "00011111",11892 => "11010011",11893 => "00111110",11894 => "00000111",11895 => "01101110",11896 => "10011001",11897 => "11011010",11898 => "00111101",11899 => "11111000",11900 => "10101100",11901 => "01000001",11902 => "00011100",11903 => "10011000",11904 => "10100101",11905 => "01000000",11906 => "00110101",11907 => "10110000",11908 => "10111111",11909 => "10011011",11910 => "11110011",11911 => "10001011",11912 => "00010001",11913 => "10111100",11914 => "10111000",11915 => "11010100",11916 => "00100101",11917 => "00000110",11918 => "01011010",11919 => "00000011",11920 => "01000011",11921 => "01010001",11922 => "11100010",11923 => "00111011",11924 => "11110000",11925 => "11111110",11926 => "11101001",11927 => "01100111",11928 => "11001000",11929 => "11001011",11930 => "11101100",11931 => "11111001",11932 => "01000011",11933 => "00101010",11934 => "01111011",11935 => "00010001",11936 => "11010011",11937 => "10110000",11938 => "00010101",11939 => "10100100",11940 => "00010111",11941 => "00000101",11942 => "11001000",11943 => "10000001",11944 => "00011110",11945 => "10001011",11946 => "01100101",11947 => "01010011",11948 => "10011000",11949 => "01111011",11950 => "01100110",11951 => "10110001",11952 => "10000111",11953 => "11111011",11954 => "10011110",11955 => "10101100",11956 => "01101001",11957 => "01000001",11958 => "11110110",11959 => "01001100",11960 => "01010011",11961 => "11000111",11962 => "00110000",11963 => "01110101",11964 => "00110011",11965 => "00101100",11966 => "10011100",11967 => "11011000",11968 => "00010010",11969 => "01000111",11970 => "01011001",11971 => "01000001",11972 => "01101011",11973 => "00111100",11974 => "01010100",11975 => "00000010",11976 => "00101001",11977 => "01011000",11978 => "11101001",11979 => "10011011",11980 => "10010000",11981 => "11101001",11982 => "01100001",11983 => "00011011",11984 => "10100101",11985 => "11100111",11986 => "01101010",11987 => "00110010",11988 => "00100110",11989 => "10100010",11990 => "01011101",11991 => "01010111",11992 => "10110101",11993 => "10110110",11994 => "10101011",11995 => "10000011",11996 => "11010111",11997 => "00010011",11998 => "01000001",11999 => "01100011",12000 => "11001111",12001 => "00011001",12002 => "01001001",12003 => "10000011",12004 => "01111101",12005 => "00110101",12006 => "00011011",12007 => "11001000",12008 => "10111101",12009 => "10000111",12010 => "01010011",12011 => "00000000",12012 => "10101101",12013 => "01010001",12014 => "00111110",12015 => "10000100",12016 => "11101101",12017 => "11111011",12018 => "01001001",12019 => "10101010",12020 => "01000010",12021 => "00111001",12022 => "11010101",12023 => "00010010",12024 => "10110001",12025 => "10001111",12026 => "00110011",12027 => "10100111",12028 => "10000000",12029 => "01101101",12030 => "00001000",12031 => "10111101",12032 => "10011000",12033 => "10110010",12034 => "00011011",12035 => "11101010",12036 => "10110010",12037 => "00110011",12038 => "11001000",12039 => "01010001",12040 => "01110110",12041 => "11011111",12042 => "00000111",12043 => "01001011",12044 => "00001001",12045 => "01100001",12046 => "10001100",12047 => "11101001",12048 => "01010111",12049 => "00100101",12050 => "10101011",12051 => "10100110",12052 => "10100000",12053 => "11010101",12054 => "01001111",12055 => "11000011",12056 => "10111110",12057 => "11010101",12058 => "11101110",12059 => "10000001",12060 => "10101100",12061 => "11001110",12062 => "11111000",12063 => "10010100",12064 => "00011000",12065 => "11010010",12066 => "01111101",12067 => "01101011",12068 => "11110000",12069 => "01001010",12070 => "11111111",12071 => "01111010",12072 => "10101001",12073 => "00010011",12074 => "01011001",12075 => "00110111",12076 => "00111111",12077 => "01001111",12078 => "00000011",12079 => "00011000",12080 => "01111010",12081 => "01100011",12082 => "11110001",12083 => "11001110",12084 => "00001011",12085 => "00111110",12086 => "11110010",12087 => "10011010",12088 => "10100101",12089 => "00111101",12090 => "01110011",12091 => "11001101",12092 => "01010001",12093 => "00101000",12094 => "10000001",12095 => "00110010",12096 => "11000111",12097 => "10111101",12098 => "01011010",12099 => "11011110",12100 => "10111110",12101 => "00010001",12102 => "10101100",12103 => "10011111",12104 => "10011011",12105 => "10110111",12106 => "11011000",12107 => "01100011",12108 => "00100101",12109 => "01010101",12110 => "00110110",12111 => "11101101",12112 => "10110000",12113 => "11010111",12114 => "01111101",12115 => "00010100",12116 => "11001011",12117 => "11011100",12118 => "00110111",12119 => "01110010",12120 => "00110001",12121 => "10101110",12122 => "10010011",12123 => "00001001",12124 => "10010100",12125 => "11011110",12126 => "11011011",12127 => "11111111",12128 => "11001010",12129 => "10001001",12130 => "01000010",12131 => "00011111",12132 => "01111111",12133 => "10001100",12134 => "01001011",12135 => "11100100",12136 => "11000100",12137 => "00110110",12138 => "01000010",12139 => "10111101",12140 => "10010111",12141 => "10100111",12142 => "10010101",12143 => "10110110",12144 => "01011011",12145 => "10100100",12146 => "01110000",12147 => "00000110",12148 => "11110000",12149 => "11011011",12150 => "11001100",12151 => "01011001",12152 => "10000011",12153 => "01100111",12154 => "01010110",12155 => "10011011",12156 => "01000010",12157 => "11000011",12158 => "01010001",12159 => "11110111",12160 => "00011111",12161 => "00111011",12162 => "00101001",12163 => "10110111",12164 => "11100100",12165 => "10101101",12166 => "01000000",12167 => "11011100",12168 => "10010011",12169 => "10011001",12170 => "01111110",12171 => "00001111",12172 => "00011000",12173 => "00001010",12174 => "00011100",12175 => "01000101",12176 => "10101010",12177 => "10010100",12178 => "01010111",12179 => "11100100",12180 => "11100101",12181 => "11100011",12182 => "00000000",12183 => "10000010",12184 => "00110010",12185 => "00100101",12186 => "01101001",12187 => "10000000",12188 => "10111111",12189 => "11101100",12190 => "00100101",12191 => "00100011",12192 => "10111100",12193 => "10101111",12194 => "11100000",12195 => "10011100",12196 => "11100001",12197 => "10010010",12198 => "11011111",12199 => "00011100",12200 => "10001101",12201 => "00101000",12202 => "00100101",12203 => "10111100",12204 => "10011100",12205 => "11111001",12206 => "00111111",12207 => "01101111",12208 => "00111000",12209 => "10101110",12210 => "11000010",12211 => "10000111",12212 => "10111001",12213 => "00010101",12214 => "10011001",12215 => "00011001",12216 => "10011111",12217 => "11010100",12218 => "00000110",12219 => "11000001",12220 => "10011110",12221 => "10011001",12222 => "10010101",12223 => "00010010",12224 => "01010001",12225 => "11001101",12226 => "01100011",12227 => "00011001",12228 => "01000101",12229 => "10111110",12230 => "11000011",12231 => "11000001",12232 => "10000000",12233 => "00110100",12234 => "01110001",12235 => "11010101",12236 => "01001100",12237 => "01011000",12238 => "11110100",12239 => "00101010",12240 => "10001010",12241 => "01111111",12242 => "00001000",12243 => "01001010",12244 => "11100100",12245 => "01000001",12246 => "10100111",12247 => "10010100",12248 => "10110111",12249 => "10011100",12250 => "00001000",12251 => "11000001",12252 => "01010010",12253 => "01010001",12254 => "11011100",12255 => "10100111",12256 => "01010100",12257 => "10110011",12258 => "10111000",12259 => "00100011",12260 => "11000000",12261 => "11101010",12262 => "01110110",12263 => "00001010",12264 => "11010011",12265 => "01100000",12266 => "01000110",12267 => "11000100",12268 => "11110101",12269 => "00011000",12270 => "01011110",12271 => "11101001",12272 => "01100011",12273 => "01111111",12274 => "00101010",12275 => "00110011",12276 => "10011010",12277 => "10100110",12278 => "00101111",12279 => "00010110",12280 => "10100101",12281 => "10101110",12282 => "10000011",12283 => "10011111",12284 => "10110010",12285 => "00100001",12286 => "11110100",12287 => "10101100",12288 => "00110000",12289 => "01001111",12290 => "11100011",12291 => "00101000",12292 => "10111010",12293 => "10001000",12294 => "10101110",12295 => "11000010",12296 => "11010010",12297 => "00101011",12298 => "11111110",12299 => "10010000",12300 => "10001111",12301 => "01010010",12302 => "10110101",12303 => "10001101",12304 => "01011000",12305 => "01110110",12306 => "00000010",12307 => "01110100",12308 => "00111100",12309 => "00110100",12310 => "01100111",12311 => "01010100",12312 => "10111011",12313 => "11100001",12314 => "01000001",12315 => "00100101",12316 => "01100110",12317 => "01011101",12318 => "10010101",12319 => "01110001",12320 => "10000010",12321 => "10010001",12322 => "10010101",12323 => "11101111",12324 => "10111000",12325 => "00110011",12326 => "10000110",12327 => "01111111",12328 => "10101011",12329 => "11000100",12330 => "00000111",12331 => "10000100",12332 => "11100111",12333 => "10101110",12334 => "10000000",12335 => "00110110",12336 => "11001101",12337 => "00100000",12338 => "00000000",12339 => "11111100",12340 => "01000110",12341 => "00010001",12342 => "10110001",12343 => "01011111",12344 => "01000000",12345 => "01011011",12346 => "00111110",12347 => "11110111",12348 => "01001100",12349 => "01111111",12350 => "01101111",12351 => "00010010",12352 => "11111100",12353 => "11101000",12354 => "01101000",12355 => "10110100",12356 => "10011100",12357 => "01000101",12358 => "01100111",12359 => "11110001",12360 => "11010011",12361 => "00001100",12362 => "00001110",12363 => "10001010",12364 => "11011010",12365 => "11100111",12366 => "10111000",12367 => "10111101",12368 => "10010111",12369 => "00100101",12370 => "00100010",12371 => "01100111",12372 => "11100100",12373 => "00101001",12374 => "11101110",12375 => "00010000",12376 => "00010110",12377 => "10110010",12378 => "11010001",12379 => "10100000",12380 => "00000110",12381 => "11010101",12382 => "11100000",12383 => "00010010",12384 => "11001100",12385 => "10011111",12386 => "01101110",12387 => "10000001",12388 => "11110011",12389 => "01001011",12390 => "00011110",12391 => "10011000",12392 => "11100111",12393 => "01010000",12394 => "00010100",12395 => "01000101",12396 => "01111111",12397 => "01111111",12398 => "10010111",12399 => "01110001",12400 => "01110111",12401 => "01011110",12402 => "10101011",12403 => "01110011",12404 => "00010011",12405 => "11100101",12406 => "01100100",12407 => "11101010",12408 => "11100000",12409 => "00001101",12410 => "10111110",12411 => "11011110",12412 => "11110101",12413 => "11000101",12414 => "11100011",12415 => "10101100",12416 => "00010111",12417 => "10010011",12418 => "01100110",12419 => "11010111",12420 => "01101001",12421 => "00100011",12422 => "10010001",12423 => "01100011",12424 => "11000000",12425 => "10101000",12426 => "01111101",12427 => "00001100",12428 => "01111100",12429 => "00010100",12430 => "01111101",12431 => "11110001",12432 => "00110001",12433 => "11010010",12434 => "10000111",12435 => "10110001",12436 => "01111001",12437 => "10011100",12438 => "11010100",12439 => "01000100",12440 => "10101010",12441 => "11111001",12442 => "01010011",12443 => "10100011",12444 => "00011111",12445 => "00110001",12446 => "00000010",12447 => "01011011",12448 => "11100001",12449 => "01110111",12450 => "01011010",12451 => "11110111",12452 => "10011101",12453 => "01101101",12454 => "01000101",12455 => "11111100",12456 => "10100111",12457 => "00001111",12458 => "01111000",12459 => "10101010",12460 => "11011110",12461 => "01100011",12462 => "00011000",12463 => "00001111",12464 => "10101110",12465 => "10000111",12466 => "10011011",12467 => "01011010",12468 => "00100010",12469 => "00101010",12470 => "11100011",12471 => "00001111",12472 => "00100011",12473 => "11011110",12474 => "01110010",12475 => "01110001",12476 => "00110010",12477 => "00111111",12478 => "00111101",12479 => "11001111",12480 => "00011110",12481 => "10001100",12482 => "10111000",12483 => "01101111",12484 => "01010101",12485 => "01101101",12486 => "01110001",12487 => "00100100",12488 => "00010010",12489 => "10010000",12490 => "00111100",12491 => "11001011",12492 => "00110001",12493 => "11100001",12494 => "01111111",12495 => "10010001",12496 => "01110100",12497 => "10000111",12498 => "11111110",12499 => "00111001",12500 => "11101101",12501 => "11010000",12502 => "01100111",12503 => "11001000",12504 => "00110111",12505 => "00000111",12506 => "01110100",12507 => "11111000",12508 => "00001000",12509 => "11000111",12510 => "00111011",12511 => "11100010",12512 => "00011101",12513 => "01000100",12514 => "10110011",12515 => "10010110",12516 => "11010000",12517 => "10100010",12518 => "01001001",12519 => "00011011",12520 => "01011110",12521 => "01111101",12522 => "01010001",12523 => "11111001",12524 => "11001011",12525 => "00101100",12526 => "00000011",12527 => "01101010",12528 => "00001111",12529 => "01001011",12530 => "11110110",12531 => "00000110",12532 => "01011010",12533 => "01100010",12534 => "10101100",12535 => "00010111",12536 => "11001000",12537 => "10111100",12538 => "00000100",12539 => "11010111",12540 => "01110001",12541 => "10000010",12542 => "01111011",12543 => "11000100",12544 => "00010001",12545 => "01001011",12546 => "00111000",12547 => "00010111",12548 => "01010100",12549 => "00001101",12550 => "10111010",12551 => "10111010",12552 => "01001010",12553 => "10011101",12554 => "00101101",12555 => "10111000",12556 => "10110000",12557 => "11110101",12558 => "11111000",12559 => "10000101",12560 => "00011101",12561 => "10011100",12562 => "00011101",12563 => "00101100",12564 => "11101000",12565 => "00001011",12566 => "00011010",12567 => "01001111",12568 => "01101101",12569 => "10111010",12570 => "01011000",12571 => "10010001",12572 => "01000010",12573 => "11001111",12574 => "00000100",12575 => "01011110",12576 => "10111101",12577 => "10010101",12578 => "11010001",12579 => "10100111",12580 => "11011011",12581 => "01101110",12582 => "00001000",12583 => "01000010",12584 => "11101011",12585 => "10110001",12586 => "10010101",12587 => "11110011",12588 => "10001001",12589 => "11100101",12590 => "01111001",12591 => "01110010",12592 => "00011011",12593 => "10101110",12594 => "01100010",12595 => "10101010",12596 => "10000010",12597 => "00101111",12598 => "11010000",12599 => "00110001",12600 => "11111011",12601 => "01010000",12602 => "11110100",12603 => "00111110",12604 => "01011010",12605 => "11010110",12606 => "00111000",12607 => "01101111",12608 => "01100000",12609 => "11100011",12610 => "10011011",12611 => "10110001",12612 => "11100110",12613 => "10110010",12614 => "11111101",12615 => "00110111",12616 => "01011100",12617 => "11001011",12618 => "01100111",12619 => "00011010",12620 => "11110011",12621 => "11000100",12622 => "11011101",12623 => "00010000",12624 => "00100011",12625 => "01101110",12626 => "11000011",12627 => "10111011",12628 => "01011100",12629 => "00001110",12630 => "11011111",12631 => "00101111",12632 => "01111100",12633 => "01001111",12634 => "01011010",12635 => "10011111",12636 => "10010011",12637 => "10010100",12638 => "10000001",12639 => "10000100",12640 => "11010111",12641 => "10110010",12642 => "00011100",12643 => "11001101",12644 => "00011111",12645 => "11000111",12646 => "10111011",12647 => "11101000",12648 => "11100111",12649 => "00001110",12650 => "11000010",12651 => "00000100",12652 => "00000000",12653 => "00000000",12654 => "01110001",12655 => "00010110",12656 => "01110000",12657 => "00101011",12658 => "10100011",12659 => "11000111",12660 => "00111101",12661 => "11001110",12662 => "11100000",12663 => "01001100",12664 => "10111010",12665 => "10101100",12666 => "10101101",12667 => "11000000",12668 => "00000101",12669 => "11101011",12670 => "11100010",12671 => "10100111",12672 => "01100101",12673 => "10110000",12674 => "11111010",12675 => "01010011",12676 => "01000011",12677 => "00010001",12678 => "01111101",12679 => "01011100",12680 => "11110010",12681 => "01110101",12682 => "11001011",12683 => "00010101",12684 => "10001001",12685 => "00100000",12686 => "10111101",12687 => "00100101",12688 => "10001101",12689 => "10101110",12690 => "10111101",12691 => "00000010",12692 => "11110000",12693 => "11011001",12694 => "11111100",12695 => "01110111",12696 => "01110110",12697 => "01101100",12698 => "01111000",12699 => "11110000",12700 => "11111011",12701 => "00111010",12702 => "11010011",12703 => "01010000",12704 => "10010101",12705 => "11011110",12706 => "01101111",12707 => "01111011",12708 => "01001101",12709 => "10101000",12710 => "11100011",12711 => "11010000",12712 => "11101110",12713 => "01000001",12714 => "10110011",12715 => "10111111",12716 => "00100001",12717 => "01001001",12718 => "10110110",12719 => "01001111",12720 => "11010000",12721 => "01000011",12722 => "01110000",12723 => "01010110",12724 => "11000110",12725 => "01110110",12726 => "10011000",12727 => "00110011",12728 => "11000001",12729 => "11110001",12730 => "00000110",12731 => "10101010",12732 => "01101001",12733 => "00000111",12734 => "00010000",12735 => "01000001",12736 => "01010000",12737 => "01001001",12738 => "10101011",12739 => "10101001",12740 => "10001010",12741 => "01111000",12742 => "00010100",12743 => "11110111",12744 => "01011111",12745 => "11010100",12746 => "10110011",12747 => "00010111",12748 => "11010111",12749 => "00011111",12750 => "10000100",12751 => "11000111",12752 => "01100011",12753 => "01000000",12754 => "11001101",12755 => "01101010",12756 => "00000010",12757 => "00111111",12758 => "11100101",12759 => "00000000",12760 => "11001100",12761 => "11100100",12762 => "01011111",12763 => "01110100",12764 => "01111011",12765 => "10011000",12766 => "01111100",12767 => "01000011",12768 => "10010000",12769 => "01101100",12770 => "01100110",12771 => "11001010",12772 => "10000110",12773 => "00010000",12774 => "11111011",12775 => "10100101",12776 => "10001111",12777 => "10101011",12778 => "11100101",12779 => "01110000",12780 => "10110100",12781 => "00111000",12782 => "11010111",12783 => "11001000",12784 => "00001011",12785 => "00010001",12786 => "01010110",12787 => "10100110",12788 => "10110001",12789 => "11101011",12790 => "10010101",12791 => "11010101",12792 => "01000100",12793 => "11010010",12794 => "01001011",12795 => "10001000",12796 => "00100001",12797 => "01001101",12798 => "00011111",12799 => "00101111",12800 => "01101100",12801 => "01100000",12802 => "00101100",12803 => "01101000",12804 => "10010111",12805 => "11010111",12806 => "10001010",12807 => "10011100",12808 => "11110111",12809 => "00110010",12810 => "00101101",12811 => "11101101",12812 => "10000111",12813 => "10111100",12814 => "11110100",12815 => "10100011",12816 => "11001011",12817 => "11100110",12818 => "00001110",12819 => "01100001",12820 => "01100011",12821 => "00100001",12822 => "10110110",12823 => "00011101",12824 => "11011010",12825 => "11001110",12826 => "01101101",12827 => "01111011",12828 => "00110100",12829 => "01110100",12830 => "00110101",12831 => "00110000",12832 => "01000010",12833 => "01010011",12834 => "11000000",12835 => "11000111",12836 => "01001101",12837 => "00101111",12838 => "11000001",12839 => "01001011",12840 => "10101111",12841 => "11000100",12842 => "01100010",12843 => "01111101",12844 => "00111100",12845 => "01001100",12846 => "10010101",12847 => "01001110",12848 => "01111001",12849 => "10111000",12850 => "01000000",12851 => "11000110",12852 => "10100111",12853 => "10010011",12854 => "01110111",12855 => "11100000",12856 => "11110001",12857 => "10010011",12858 => "11010010",12859 => "10000010",12860 => "10011110",12861 => "00000010",12862 => "11000111",12863 => "11101000",12864 => "11010000",12865 => "10001100",12866 => "01011111",12867 => "01010001",12868 => "01111100",12869 => "00111011",12870 => "01010101",12871 => "01010011",12872 => "00110001",12873 => "01111000",12874 => "01111010",12875 => "00110000",12876 => "01110100",12877 => "11101000",12878 => "10100100",12879 => "00000111",12880 => "11011100",12881 => "01101011",12882 => "10010110",12883 => "01111110",12884 => "11010101",12885 => "01010100",12886 => "10101001",12887 => "00110111",12888 => "11011101",12889 => "11000100",12890 => "11100010",12891 => "10100010",12892 => "11100110",12893 => "11100100",12894 => "10101010",12895 => "00111100",12896 => "01101100",12897 => "01101010",12898 => "01001111",12899 => "00010001",12900 => "11101111",12901 => "10011000",12902 => "01010001",12903 => "01100110",12904 => "11101101",12905 => "10100111",12906 => "10011001",12907 => "10110000",12908 => "00111101",12909 => "10100110",12910 => "10110001",12911 => "00111000",12912 => "01111000",12913 => "01101111",12914 => "00100001",12915 => "10110001",12916 => "01111010",12917 => "00100110",12918 => "11110000",12919 => "01111010",12920 => "10100000",12921 => "11100111",12922 => "10100000",12923 => "00110100",12924 => "00000000",12925 => "11110000",12926 => "01000110",12927 => "01111101",12928 => "11001101",12929 => "10111011",12930 => "01010011",12931 => "00001000",12932 => "11100001",12933 => "11101010",12934 => "01100100",12935 => "11011110",12936 => "10100010",12937 => "10011111",12938 => "01001110",12939 => "11010111",12940 => "01100010",12941 => "10100100",12942 => "00101001",12943 => "10011010",12944 => "01001110",12945 => "10110101",12946 => "00001111",12947 => "00111111",12948 => "10100101",12949 => "01101011",12950 => "01111011",12951 => "00100011",12952 => "10101000",12953 => "10011010",12954 => "11110101",12955 => "00000011",12956 => "10000111",12957 => "00111011",12958 => "00010101",12959 => "11000000",12960 => "11111110",12961 => "01010100",12962 => "01100001",12963 => "10110110",12964 => "11000011",12965 => "00000100",12966 => "01100000",12967 => "01000011",12968 => "00110101",12969 => "11100101",12970 => "10101001",12971 => "11010000",12972 => "00011000",12973 => "11011001",12974 => "00110101",12975 => "00010110",12976 => "00000100",12977 => "10011011",12978 => "00110111",12979 => "01101100",12980 => "00011010",12981 => "00111001",12982 => "10010100",12983 => "00011001",12984 => "10011110",12985 => "01111101",12986 => "01011111",12987 => "11000100",12988 => "00110001",12989 => "10010101",12990 => "10010111",12991 => "00111101",12992 => "11000011",12993 => "11010010",12994 => "10010010",12995 => "01000101",12996 => "00011110",12997 => "00101101",12998 => "00101111",12999 => "10010000",13000 => "01110011",13001 => "00110100",13002 => "11101000",13003 => "00000101",13004 => "11111000",13005 => "10010100",13006 => "10110111",13007 => "10101110",13008 => "00000000",13009 => "01110011",13010 => "11101001",13011 => "01111110",13012 => "01100010",13013 => "00000000",13014 => "10101110",13015 => "11111101",13016 => "11100010",13017 => "00100110",13018 => "11000010",13019 => "10110100",13020 => "11100000",13021 => "01010111",13022 => "10000111",13023 => "00011010",13024 => "11110111",13025 => "11010110",13026 => "00000110",13027 => "01000111",13028 => "10101110",13029 => "00111101",13030 => "11000111",13031 => "10001001",13032 => "10000100",13033 => "11110100",13034 => "00111101",13035 => "00001001",13036 => "10011110",13037 => "11010010",13038 => "00101001",13039 => "10110011",13040 => "00010000",13041 => "01010110",13042 => "11110110",13043 => "10101000",13044 => "11101000",13045 => "10010100",13046 => "00101000",13047 => "00001011",13048 => "11000011",13049 => "11000011",13050 => "00011111",13051 => "01101101",13052 => "10010110",13053 => "00010100",13054 => "00000011",13055 => "10001111",13056 => "11101100",13057 => "10111100",13058 => "10110100",13059 => "10101001",13060 => "10111111",13061 => "01000001",13062 => "10101110",13063 => "11001111",13064 => "01100110",13065 => "10001010",13066 => "11110011",13067 => "00001010",13068 => "01111011",13069 => "00001100",13070 => "01111100",13071 => "10111010",13072 => "11101000",13073 => "01100011",13074 => "01100001",13075 => "10010011",13076 => "00001010",13077 => "10100000",13078 => "10110100",13079 => "11111101",13080 => "10111001",13081 => "00001010",13082 => "10101101",13083 => "10111001",13084 => "11010110",13085 => "00110110",13086 => "11110010",13087 => "01110010",13088 => "00100100",13089 => "01101111",13090 => "10010111",13091 => "10101100",13092 => "11100010",13093 => "11100010",13094 => "11011101",13095 => "01101100",13096 => "01001010",13097 => "11011010",13098 => "10001101",13099 => "10111100",13100 => "01111100",13101 => "11011000",13102 => "10010011",13103 => "01001111",13104 => "01101001",13105 => "11011110",13106 => "10010110",13107 => "01001001",13108 => "00100010",13109 => "01111110",13110 => "10101000",13111 => "10000011",13112 => "01001000",13113 => "10100100",13114 => "00001101",13115 => "11111101",13116 => "10010001",13117 => "11101111",13118 => "00001000",13119 => "11100110",13120 => "00101101",13121 => "11101110",13122 => "10000011",13123 => "11011011",13124 => "11000100",13125 => "01100111",13126 => "11000101",13127 => "11011000",13128 => "00001111",13129 => "10011110",13130 => "01101000",13131 => "00010111",13132 => "10000000",13133 => "10001000",13134 => "10111011",13135 => "00101010",13136 => "10000110",13137 => "11101001",13138 => "01000100",13139 => "10001000",13140 => "10000111",13141 => "01011000",13142 => "10100100",13143 => "11000001",13144 => "11101100",13145 => "11000010",13146 => "10110110",13147 => "11100101",13148 => "11011101",13149 => "10011010",13150 => "10001111",13151 => "00101001",13152 => "01100010",13153 => "10011010",13154 => "10011001",13155 => "10100100",13156 => "00110010",13157 => "10110100",13158 => "01000011",13159 => "10111000",13160 => "00000011",13161 => "01000011",13162 => "11010000",13163 => "10001010",13164 => "11000010",13165 => "01111101",13166 => "01000011",13167 => "10011100",13168 => "00110100",13169 => "11101110",13170 => "11010101",13171 => "10010100",13172 => "10100110",13173 => "10110111",13174 => "01001001",13175 => "01101010",13176 => "01001110",13177 => "01001010",13178 => "01110010",13179 => "11100000",13180 => "11010000",13181 => "10001111",13182 => "11001001",13183 => "00010000",13184 => "11000001",13185 => "11110010",13186 => "01011111",13187 => "10011111",13188 => "00111101",13189 => "11110010",13190 => "10000101",13191 => "10001100",13192 => "01000000",13193 => "01110000",13194 => "00011001",13195 => "00100011",13196 => "10110101",13197 => "11101001",13198 => "01111001",13199 => "11010000",13200 => "00011000",13201 => "01101100",13202 => "10001000",13203 => "00011001",13204 => "01011110",13205 => "00110101",13206 => "01000010",13207 => "11101011",13208 => "11000100",13209 => "11100101",13210 => "01001111",13211 => "10111001",13212 => "01011101",13213 => "00000011",13214 => "11100010",13215 => "10101011",13216 => "10110100",13217 => "00111000",13218 => "01101110",13219 => "00010001",13220 => "11010111",13221 => "11111110",13222 => "01011010",13223 => "11111110",13224 => "10001100",13225 => "11000010",13226 => "01010010",13227 => "11010100",13228 => "11111111",13229 => "10010110",13230 => "01011000",13231 => "10100011",13232 => "10010011",13233 => "10100111",13234 => "00100010",13235 => "10000000",13236 => "00000111",13237 => "00110000",13238 => "11001010",13239 => "01001111",13240 => "00111011",13241 => "00100100",13242 => "11000100",13243 => "00000101",13244 => "01111111",13245 => "11001001",13246 => "10000001",13247 => "01110100",13248 => "01010100",13249 => "00010010",13250 => "00011010",13251 => "00101100",13252 => "10101111",13253 => "11111001",13254 => "01101010",13255 => "00011101",13256 => "10000001",13257 => "01000111",13258 => "10001011",13259 => "11111010",13260 => "10001100",13261 => "10000111",13262 => "11010110",13263 => "11001110",13264 => "01001001",13265 => "10011110",13266 => "00001111",13267 => "01111000",13268 => "01011111",13269 => "01011101",13270 => "11100011",13271 => "11001011",13272 => "01101111",13273 => "11101001",13274 => "01111000",13275 => "11000010",13276 => "10001110",13277 => "01010101",13278 => "11001001",13279 => "11000111",13280 => "01111001",13281 => "00111101",13282 => "10010101",13283 => "00110101",13284 => "11111110",13285 => "00100000",13286 => "00111100",13287 => "11101110",13288 => "00000000",13289 => "10000101",13290 => "01110111",13291 => "10011110",13292 => "11100100",13293 => "01101010",13294 => "01101101",13295 => "00110110",13296 => "00010001",13297 => "00110001",13298 => "11001110",13299 => "10101111",13300 => "10010000",13301 => "11110100",13302 => "00011011",13303 => "01101001",13304 => "01011001",13305 => "01010010",13306 => "00101101",13307 => "00000100",13308 => "11001001",13309 => "00001011",13310 => "01010110",13311 => "01010111",13312 => "01001010",13313 => "00101111",13314 => "11001100",13315 => "00000110",13316 => "11111001",13317 => "00100110",13318 => "10101100",13319 => "10101010",13320 => "01111010",13321 => "10111101",13322 => "11000100",13323 => "11110000",13324 => "11011001",13325 => "10101110",13326 => "11011110",13327 => "00110111",13328 => "00011000",13329 => "00000000",13330 => "10110100",13331 => "00010011",13332 => "11111100",13333 => "11110000",13334 => "10000101",13335 => "01101010",13336 => "01000001",13337 => "10000011",13338 => "00100110",13339 => "00011111",13340 => "00111111",13341 => "01010011",13342 => "00000100",13343 => "10110010",13344 => "11000111",13345 => "10001110",13346 => "01110001",13347 => "10111011",13348 => "01000011",13349 => "10001000",13350 => "00010101",13351 => "01001110",13352 => "00000111",13353 => "10010101",13354 => "11001010",13355 => "11101000",13356 => "00100000",13357 => "11101000",13358 => "01110000",13359 => "10101001",13360 => "11100001",13361 => "01001101",13362 => "01010010",13363 => "00100001",13364 => "00010100",13365 => "01001010",13366 => "00001111",13367 => "11110000",13368 => "01111110",13369 => "10110010",13370 => "00101101",13371 => "01101101",13372 => "00000100",13373 => "01100011",13374 => "11011000",13375 => "10100010",13376 => "00001001",13377 => "11011110",13378 => "10001111",13379 => "11001011",13380 => "00101110",13381 => "10111111",13382 => "00111000",13383 => "01101101",13384 => "00011011",13385 => "01011101",13386 => "01000101",13387 => "00010111",13388 => "10101101",13389 => "11000111",13390 => "10101011",13391 => "00010001",13392 => "01100000",13393 => "11001110",13394 => "10000000",13395 => "10110011",13396 => "01000101",13397 => "11001100",13398 => "11101001",13399 => "11101010",13400 => "11101010",13401 => "11011110",13402 => "01000100",13403 => "01101110",13404 => "10010100",13405 => "00100101",13406 => "10111101",13407 => "10110110",13408 => "00010101",13409 => "10000001",13410 => "01101011",13411 => "11111001",13412 => "10101010",13413 => "11010100",13414 => "01101010",13415 => "10111110",13416 => "01110010",13417 => "00111000",13418 => "11110001",13419 => "00011100",13420 => "11001011",13421 => "10101011",13422 => "00100001",13423 => "01010001",13424 => "10110010",13425 => "11010010",13426 => "11011110",13427 => "01010000",13428 => "00011101",13429 => "11100001",13430 => "00000000",13431 => "11001001",13432 => "10001011",13433 => "10100011",13434 => "10001100",13435 => "00001011",13436 => "01101110",13437 => "10111111",13438 => "10100100",13439 => "01110101",13440 => "01101100",13441 => "11111011",13442 => "10110110",13443 => "11001101",13444 => "00101010",13445 => "10001110",13446 => "01001000",13447 => "01101010",13448 => "11001000",13449 => "00000010",13450 => "10010010",13451 => "11000101",13452 => "01000000",13453 => "11000101",13454 => "10101101",13455 => "01000001",13456 => "11110110",13457 => "01001100",13458 => "00011110",13459 => "11001010",13460 => "00101001",13461 => "01111011",13462 => "11001001",13463 => "10000101",13464 => "01100000",13465 => "00101110",13466 => "00101000",13467 => "00110111",13468 => "00111111",13469 => "11100101",13470 => "11010111",13471 => "10000101",13472 => "00001011",13473 => "10011011",13474 => "01110110",13475 => "11110011",13476 => "10010011",13477 => "00111000",13478 => "00000110",13479 => "11110100",13480 => "00100011",13481 => "11000010",13482 => "00110011",13483 => "01111010",13484 => "00100100",13485 => "00010010",13486 => "10100111",13487 => "01110100",13488 => "10001110",13489 => "01001001",13490 => "10001001",13491 => "01111000",13492 => "11101001",13493 => "10010001",13494 => "01011011",13495 => "11100101",13496 => "11100010",13497 => "11011001",13498 => "01011101",13499 => "01011110",13500 => "11010010",13501 => "10110011",13502 => "10001111",13503 => "00001001",13504 => "10101000",13505 => "10010010",13506 => "10010010",13507 => "01101110",13508 => "11110110",13509 => "01101101",13510 => "01101010",13511 => "01000000",13512 => "10010001",13513 => "01010110",13514 => "11101001",13515 => "01000111",13516 => "01011100",13517 => "11010110",13518 => "01100100",13519 => "11010110",13520 => "11010000",13521 => "11110010",13522 => "00001011",13523 => "01000110",13524 => "00110101",13525 => "11011010",13526 => "00110110",13527 => "11001001",13528 => "10100101",13529 => "11101110",13530 => "01110010",13531 => "10010101",13532 => "11101010",13533 => "01000111",13534 => "00001110",13535 => "11111110",13536 => "00011111",13537 => "00110101",13538 => "11100001",13539 => "10010111",13540 => "11010000",13541 => "01111000",13542 => "10001000",13543 => "01001011",13544 => "10101010",13545 => "01100011",13546 => "10011011",13547 => "01101100",13548 => "00011100",13549 => "01111100",13550 => "00101011",13551 => "01100011",13552 => "01101011",13553 => "00010010",13554 => "10101101",13555 => "00000100",13556 => "01111011",13557 => "00000010",13558 => "11110001",13559 => "00110010",13560 => "10111011",13561 => "10000111",13562 => "11010101",13563 => "10011010",13564 => "00101010",13565 => "00000001",13566 => "01101101",13567 => "10111101",13568 => "00110111",13569 => "10101101",13570 => "01001010",13571 => "00000001",13572 => "10000001",13573 => "01000111",13574 => "10000001",13575 => "11011100",13576 => "10100001",13577 => "01000111",13578 => "11000011",13579 => "10001100",13580 => "11100010",13581 => "01000100",13582 => "00110111",13583 => "11100010",13584 => "11011110",13585 => "00100001",13586 => "01101010",13587 => "01111000",13588 => "11111111",13589 => "01010111",13590 => "10001001",13591 => "00101100",13592 => "01101010",13593 => "10101001",13594 => "11010001",13595 => "01011001",13596 => "10111110",13597 => "00011000",13598 => "00100101",13599 => "11110010",13600 => "01011100",13601 => "00111001",13602 => "01001011",13603 => "01010001",13604 => "00110110",13605 => "10011100",13606 => "01111000",13607 => "11111101",13608 => "10111111",13609 => "01110110",13610 => "00101100",13611 => "01100010",13612 => "00110010",13613 => "10100000",13614 => "00111110",13615 => "10111110",13616 => "11100111",13617 => "11010111",13618 => "01100110",13619 => "01000101",13620 => "10111000",13621 => "01111111",13622 => "11000000",13623 => "01111111",13624 => "11111001",13625 => "00110111",13626 => "10010010",13627 => "10100000",13628 => "11101101",13629 => "10010100",13630 => "10111010",13631 => "00011000",13632 => "00100000",13633 => "11100100",13634 => "10000111",13635 => "11011110",13636 => "10111111",13637 => "10010100",13638 => "11000011",13639 => "01010100",13640 => "11001011",13641 => "01100000",13642 => "10100111",13643 => "01011100",13644 => "01101111",13645 => "01111010",13646 => "11110111",13647 => "00110000",13648 => "01111101",13649 => "10110111",13650 => "01110111",13651 => "01100100",13652 => "00100001",13653 => "00111001",13654 => "10001101",13655 => "01000011",13656 => "00100011",13657 => "11000010",13658 => "01111100",13659 => "10011101",13660 => "10110011",13661 => "10001110",13662 => "10000110",13663 => "00110000",13664 => "11111000",13665 => "01001000",13666 => "10011101",13667 => "01001000",13668 => "10000111",13669 => "10110101",13670 => "11001100",13671 => "10100110",13672 => "10011111",13673 => "11100111",13674 => "00011001",13675 => "10101110",13676 => "11011000",13677 => "01000000",13678 => "00100010",13679 => "00101000",13680 => "10111011",13681 => "10111100",13682 => "01101111",13683 => "10110101",13684 => "11001010",13685 => "01001101",13686 => "10010010",13687 => "10011011",13688 => "11110100",13689 => "11110110",13690 => "11111010",13691 => "11101001",13692 => "00100100",13693 => "01011011",13694 => "01100110",13695 => "01011101",13696 => "00011100",13697 => "00011000",13698 => "00011101",13699 => "11111111",13700 => "00000001",13701 => "10010000",13702 => "11001110",13703 => "01011001",13704 => "11001000",13705 => "01001000",13706 => "10111101",13707 => "00111010",13708 => "10101100",13709 => "10100110",13710 => "10100011",13711 => "10100010",13712 => "00111110",13713 => "10111010",13714 => "01110010",13715 => "10010110",13716 => "10000010",13717 => "11001110",13718 => "01110100",13719 => "00100011",13720 => "00110101",13721 => "01101010",13722 => "01001110",13723 => "00011110",13724 => "01111000",13725 => "01010110",13726 => "10000100",13727 => "01100101",13728 => "01001011",13729 => "00000011",13730 => "10011001",13731 => "01100011",13732 => "00110110",13733 => "10011011",13734 => "00011111",13735 => "10110111",13736 => "11100101",13737 => "11000001",13738 => "11001001",13739 => "01011111",13740 => "01100000",13741 => "11011010",13742 => "01011010",13743 => "10001000",13744 => "11101010",13745 => "01100111",13746 => "01011010",13747 => "10000110",13748 => "11010011",13749 => "00010001",13750 => "10110000",13751 => "11110011",13752 => "01000101",13753 => "11110010",13754 => "10011111",13755 => "01111110",13756 => "01001101",13757 => "10101100",13758 => "10011010",13759 => "01101011",13760 => "01011010",13761 => "01000010",13762 => "10011001",13763 => "01110100",13764 => "10100011",13765 => "10101111",13766 => "01111111",13767 => "00101010",13768 => "10011111",13769 => "00000000",13770 => "10010101",13771 => "01011000",13772 => "01010111",13773 => "10000000",13774 => "11011001",13775 => "10100111",13776 => "11000001",13777 => "11110101",13778 => "01100110",13779 => "00101110",13780 => "11100110",13781 => "00100101",13782 => "11001100",13783 => "10110101",13784 => "10011110",13785 => "11001111",13786 => "01010001",13787 => "11011110",13788 => "11100110",13789 => "01010011",13790 => "10000010",13791 => "11010110",13792 => "11101010",13793 => "11000110",13794 => "01010000",13795 => "01111101",13796 => "01000101",13797 => "11110110",13798 => "10110101",13799 => "11110001",13800 => "10101011",13801 => "00011101",13802 => "01010101",13803 => "11111111",13804 => "00101100",13805 => "00110011",13806 => "10010010",13807 => "01101101",13808 => "11000110",13809 => "11010000",13810 => "11011001",13811 => "11111001",13812 => "10010111",13813 => "01001001",13814 => "01000001",13815 => "11010001",13816 => "10010000",13817 => "10001101",13818 => "10100010",13819 => "00111000",13820 => "01110101",13821 => "00101010",13822 => "01110001",13823 => "01010100",13824 => "10100111",13825 => "10001010",13826 => "01011010",13827 => "10000010",13828 => "00001100",13829 => "11101111",13830 => "10111110",13831 => "01101110",13832 => "10001010",13833 => "00000010",13834 => "00110010",13835 => "01011110",13836 => "11010011",13837 => "01000010",13838 => "01101001",13839 => "01010101",13840 => "00010111",13841 => "11011011",13842 => "11011100",13843 => "11111111",13844 => "01101011",13845 => "10011010",13846 => "10111010",13847 => "10110000",13848 => "00011111",13849 => "01111100",13850 => "01011111",13851 => "00010010",13852 => "10011110",13853 => "10110000",13854 => "10010100",13855 => "00101001",13856 => "01111010",13857 => "11011101",13858 => "00010001",13859 => "01101100",13860 => "00101100",13861 => "01100110",13862 => "01101011",13863 => "10000010",13864 => "11011001",13865 => "00110000",13866 => "00111111",13867 => "01111100",13868 => "01010101",13869 => "11000100",13870 => "01100000",13871 => "10000110",13872 => "01011101",13873 => "01011011",13874 => "01001110",13875 => "11001110",13876 => "01001101",13877 => "01100110",13878 => "11001001",13879 => "11001110",13880 => "10000110",13881 => "01101101",13882 => "10011000",13883 => "10001111",13884 => "10011111",13885 => "01110110",13886 => "01000101",13887 => "10010110",13888 => "11000110",13889 => "01110010",13890 => "00111101",13891 => "11100101",13892 => "00001111",13893 => "10111001",13894 => "11111101",13895 => "01011110",13896 => "01100011",13897 => "01001011",13898 => "00101000",13899 => "01000101",13900 => "00111010",13901 => "10101100",13902 => "00111110",13903 => "01110100",13904 => "10010111",13905 => "00000011",13906 => "00111110",13907 => "00111110",13908 => "10100111",13909 => "00111101",13910 => "00011001",13911 => "11001010",13912 => "11001011",13913 => "01111100",13914 => "11100111",13915 => "10111101",13916 => "01110010",13917 => "01101011",13918 => "10011010",13919 => "01101101",13920 => "00101000",13921 => "10001110",13922 => "00111010",13923 => "10111001",13924 => "00100011",13925 => "01000000",13926 => "11100000",13927 => "10000101",13928 => "00010110",13929 => "11001000",13930 => "00010110",13931 => "00000010",13932 => "00001011",13933 => "01011111",13934 => "10100010",13935 => "01011010",13936 => "11001110",13937 => "10100010",13938 => "00111100",13939 => "00011001",13940 => "10010001",13941 => "00001000",13942 => "00001101",13943 => "00110001",13944 => "10101001",13945 => "00011100",13946 => "10100100",13947 => "00000011",13948 => "11110010",13949 => "10011001",13950 => "10111110",13951 => "00000001",13952 => "11101100",13953 => "11110100",13954 => "00011111",13955 => "11010010",13956 => "11011000",13957 => "11110100",13958 => "00101101",13959 => "01110101",13960 => "11011101",13961 => "01011010",13962 => "11111001",13963 => "11000010",13964 => "01101111",13965 => "11110011",13966 => "00110100",13967 => "00111011",13968 => "01110011",13969 => "00000000",13970 => "11010000",13971 => "11100110",13972 => "11111010",13973 => "00010110",13974 => "11110011",13975 => "10100100",13976 => "10010000",13977 => "11111111",13978 => "00101101",13979 => "01010001",13980 => "10000110",13981 => "10010001",13982 => "01110100",13983 => "01010011",13984 => "11111111",13985 => "00000010",13986 => "01010010",13987 => "11111011",13988 => "01101001",13989 => "11000001",13990 => "11110010",13991 => "00000110",13992 => "01111001",13993 => "00101101",13994 => "10100110",13995 => "10100111",13996 => "11010100",13997 => "01110011",13998 => "10111100",13999 => "00000101",14000 => "01100111",14001 => "10110100",14002 => "00111101",14003 => "10100000",14004 => "11111110",14005 => "11101101",14006 => "10010010",14007 => "11101110",14008 => "00110000",14009 => "01000110",14010 => "01110111",14011 => "01110011",14012 => "01000111",14013 => "00000100",14014 => "00010100",14015 => "10101001",14016 => "01011100",14017 => "10100111",14018 => "11010101",14019 => "01110000",14020 => "00000100",14021 => "01011011",14022 => "01010100",14023 => "01100001",14024 => "11010111",14025 => "10110000",14026 => "10101001",14027 => "00101100",14028 => "10111100",14029 => "01010001",14030 => "00000001",14031 => "11000111",14032 => "11111000",14033 => "01111001",14034 => "00001111",14035 => "10010110",14036 => "11110010",14037 => "10110100",14038 => "11001011",14039 => "11101101",14040 => "00001100",14041 => "11000111",14042 => "11000110",14043 => "00011011",14044 => "10011111",14045 => "10100010",14046 => "00000111",14047 => "10000011",14048 => "01111111",14049 => "11000110",14050 => "00000010",14051 => "01101110",14052 => "00011011",14053 => "11110011",14054 => "11110100",14055 => "01000000",14056 => "00100000",14057 => "01011110",14058 => "11111000",14059 => "00110011",14060 => "10100110",14061 => "11010101",14062 => "01100111",14063 => "01100100",14064 => "00011010",14065 => "11111110",14066 => "11101011",14067 => "10000011",14068 => "00110101",14069 => "11101110",14070 => "10000000",14071 => "00110110",14072 => "10110101",14073 => "10010111",14074 => "00001101",14075 => "01010101",14076 => "10010110",14077 => "00001001",14078 => "01001010",14079 => "10110101",14080 => "00101111",14081 => "11111010",14082 => "11101010",14083 => "00110010",14084 => "00000001",14085 => "01011111",14086 => "10110001",14087 => "01001101",14088 => "01001000",14089 => "11111100",14090 => "00001111",14091 => "10010001",14092 => "01101101",14093 => "01100001",14094 => "00100001",14095 => "00000111",14096 => "11010111",14097 => "01100000",14098 => "01111001",14099 => "10101010",14100 => "11101101",14101 => "01011000",14102 => "01010111",14103 => "00101101",14104 => "11100110",14105 => "00010010",14106 => "00110100",14107 => "01101010",14108 => "10011000",14109 => "01101011",14110 => "10000000",14111 => "11000011",14112 => "11000101",14113 => "11101110",14114 => "01101000",14115 => "11111010",14116 => "11010110",14117 => "11010101",14118 => "00101111",14119 => "11011010",14120 => "00010010",14121 => "10100110",14122 => "01111110",14123 => "00100010",14124 => "10111010",14125 => "01111001",14126 => "00100000",14127 => "01000110",14128 => "11111110",14129 => "01101100",14130 => "11010101",14131 => "10000101",14132 => "11100001",14133 => "01000000",14134 => "11010001",14135 => "11011100",14136 => "01000110",14137 => "11000110",14138 => "01010100",14139 => "11001010",14140 => "00110111",14141 => "00101011",14142 => "10010101",14143 => "01100100",14144 => "01011000",14145 => "01011100",14146 => "11101001",14147 => "11001000",14148 => "01010111",14149 => "00000110",14150 => "00100101",14151 => "10100011",14152 => "00001000",14153 => "10000010",14154 => "10100000",14155 => "01110000",14156 => "10101100",14157 => "10111111",14158 => "00111001",14159 => "01010111",14160 => "01110111",14161 => "01101011",14162 => "00011010",14163 => "00001010",14164 => "00000001",14165 => "01001100",14166 => "01100100",14167 => "01001011",14168 => "01111011",14169 => "11011110",14170 => "00100001",14171 => "01100001",14172 => "10111110",14173 => "10010001",14174 => "00100100",14175 => "01010111",14176 => "00101001",14177 => "11101011",14178 => "10100001",14179 => "00010111",14180 => "01111001",14181 => "11000111",14182 => "00001100",14183 => "11100110",14184 => "00111101",14185 => "11110111",14186 => "00000010",14187 => "11100011",14188 => "01111110",14189 => "01010011",14190 => "00100010",14191 => "11111100",14192 => "01000010",14193 => "00110010",14194 => "11011111",14195 => "10000101",14196 => "01111101",14197 => "00010001",14198 => "10010000",14199 => "00110100",14200 => "00001011",14201 => "01001111",14202 => "10101011",14203 => "00010010",14204 => "01111000",14205 => "11111110",14206 => "00101110",14207 => "10000100",14208 => "10111000",14209 => "11111101",14210 => "10001000",14211 => "00101010",14212 => "00001001",14213 => "10100100",14214 => "11100011",14215 => "00011111",14216 => "11000100",14217 => "10101111",14218 => "11110110",14219 => "01011101",14220 => "00001001",14221 => "00111111",14222 => "10110101",14223 => "00011100",14224 => "01011011",14225 => "10110001",14226 => "11010011",14227 => "01011110",14228 => "10100111",14229 => "10011110",14230 => "01001111",14231 => "01001111",14232 => "01101111",14233 => "11010011",14234 => "10011101",14235 => "00010110",14236 => "00011011",14237 => "11101011",14238 => "00011101",14239 => "10111000",14240 => "11001010",14241 => "01101001",14242 => "11001000",14243 => "10010001",14244 => "10110010",14245 => "10010010",14246 => "00111010",14247 => "00101010",14248 => "01000010",14249 => "01101011",14250 => "10000000",14251 => "10001111",14252 => "10101110",14253 => "10111010",14254 => "00101011",14255 => "10011110",14256 => "10010001",14257 => "01111001",14258 => "11111100",14259 => "10001100",14260 => "11010011",14261 => "00110110",14262 => "10111111",14263 => "11111111",14264 => "01101111",14265 => "00110110",14266 => "10001110",14267 => "11110000",14268 => "00000011",14269 => "10100100",14270 => "10110000",14271 => "00010000",14272 => "01011011",14273 => "01100111",14274 => "01000000",14275 => "01101111",14276 => "01100101",14277 => "00100110",14278 => "01010010",14279 => "00001000",14280 => "11111010",14281 => "11111001",14282 => "00111111",14283 => "10010011",14284 => "01101010",14285 => "11001101",14286 => "00000110",14287 => "11100001",14288 => "00010010",14289 => "01110100",14290 => "10010101",14291 => "11000000",14292 => "01110010",14293 => "10100001",14294 => "11111011",14295 => "01110110",14296 => "10111101",14297 => "00010011",14298 => "10110001",14299 => "11011001",14300 => "11111000",14301 => "01000111",14302 => "10101111",14303 => "00001011",14304 => "10001001",14305 => "10111001",14306 => "10111001",14307 => "10111011",14308 => "11011010",14309 => "00101111",14310 => "01100000",14311 => "00111011",14312 => "01010011",14313 => "00001100",14314 => "01101000",14315 => "00011010",14316 => "01000010",14317 => "01010100",14318 => "00001010",14319 => "10000100",14320 => "01010101",14321 => "10111000",14322 => "00001101",14323 => "00010111",14324 => "11010111",14325 => "11111010",14326 => "00100101",14327 => "10011100",14328 => "10000110",14329 => "01101000",14330 => "01101100",14331 => "00101100",14332 => "00010100",14333 => "01111110",14334 => "11101011",14335 => "11001101",14336 => "11011000",14337 => "10111001",14338 => "10011101",14339 => "01111000",14340 => "10011010",14341 => "01110111",14342 => "00011000",14343 => "00010011",14344 => "11010110",14345 => "01000010",14346 => "01010010",14347 => "10111110",14348 => "00110011",14349 => "10001010",14350 => "00000100",14351 => "10100100",14352 => "01110110",14353 => "00111101",14354 => "00001100",14355 => "01101101",14356 => "01000001",14357 => "00110000",14358 => "00110010",14359 => "11100000",14360 => "10010011",14361 => "00000011",14362 => "01101110",14363 => "11110100",14364 => "00001110",14365 => "10110010",14366 => "00011101",14367 => "00101110",14368 => "01110110",14369 => "11110110",14370 => "10110001",14371 => "01111110",14372 => "11101101",14373 => "00001001",14374 => "11010111",14375 => "01010100",14376 => "11001010",14377 => "00111111",14378 => "10000010",14379 => "10000000",14380 => "01101000",14381 => "10100001",14382 => "00000111",14383 => "01111101",14384 => "11101000",14385 => "01011001",14386 => "10000110",14387 => "00110011",14388 => "00001010",14389 => "00011010",14390 => "10100100",14391 => "11000100",14392 => "01100010",14393 => "11010100",14394 => "10111100",14395 => "11000111",14396 => "01110000",14397 => "10000110",14398 => "00000000",14399 => "00001100",14400 => "01110101",14401 => "11100011",14402 => "01101011",14403 => "01001111",14404 => "11010000",14405 => "01110000",14406 => "10111000",14407 => "01011010",14408 => "01110100",14409 => "11001100",14410 => "11010111",14411 => "10011110",14412 => "01101101",14413 => "11111001",14414 => "01100101",14415 => "01101101",14416 => "00010010",14417 => "11111011",14418 => "10000111",14419 => "10010001",14420 => "01100000",14421 => "01001100",14422 => "10101010",14423 => "10111111",14424 => "01001010",14425 => "11000110",14426 => "10000100",14427 => "00101100",14428 => "10111101",14429 => "11000110",14430 => "11010110",14431 => "10110010",14432 => "01101110",14433 => "01100011",14434 => "10001100",14435 => "00100001",14436 => "01011010",14437 => "11111001",14438 => "01001001",14439 => "01010101",14440 => "01010111",14441 => "01011010",14442 => "10110011",14443 => "00001001",14444 => "11110101",14445 => "00111101",14446 => "10001001",14447 => "10001100",14448 => "01001010",14449 => "11110000",14450 => "00101110",14451 => "01010000",14452 => "11101001",14453 => "00011000",14454 => "00011100",14455 => "10100111",14456 => "00100100",14457 => "00001000",14458 => "01011100",14459 => "10101000",14460 => "10100101",14461 => "10110101",14462 => "11000011",14463 => "01111001",14464 => "10111110",14465 => "00000000",14466 => "10101011",14467 => "01001010",14468 => "11101001",14469 => "01100111",14470 => "11001011",14471 => "11010100",14472 => "10001100",14473 => "10100100",14474 => "10001100",14475 => "00110100",14476 => "01011101",14477 => "00101111",14478 => "00010110",14479 => "00011000",14480 => "10010000",14481 => "01100000",14482 => "10011010",14483 => "01111001",14484 => "10100011",14485 => "01111110",14486 => "01000000",14487 => "11001110",14488 => "01110000",14489 => "01010010",14490 => "11011100",14491 => "01110100",14492 => "10110001",14493 => "11000100",14494 => "00011011",14495 => "11110111",14496 => "11110010",14497 => "11110011",14498 => "11010011",14499 => "00110000",14500 => "11001110",14501 => "00110011",14502 => "11101011",14503 => "11111011",14504 => "10000111",14505 => "10101011",14506 => "00001100",14507 => "10101011",14508 => "10100111",14509 => "01000100",14510 => "10001110",14511 => "01010011",14512 => "11100101",14513 => "11011110",14514 => "01110011",14515 => "10010110",14516 => "01111110",14517 => "11000011",14518 => "10111011",14519 => "10010001",14520 => "00001101",14521 => "01101010",14522 => "00100101",14523 => "01101001",14524 => "10010111",14525 => "11111100",14526 => "10111101",14527 => "10111101",14528 => "11001101",14529 => "10100001",14530 => "10111100",14531 => "10110010",14532 => "01101100",14533 => "10100111",14534 => "00010001",14535 => "10110100",14536 => "01101101",14537 => "10011001",14538 => "01110100",14539 => "11010111",14540 => "00001111",14541 => "00010001",14542 => "10101001",14543 => "00111111",14544 => "00010010",14545 => "11110111",14546 => "11101111",14547 => "10001101",14548 => "11001001",14549 => "01010110",14550 => "10100100",14551 => "00000010",14552 => "10101110",14553 => "00100001",14554 => "00101111",14555 => "00011001",14556 => "01011111",14557 => "00110000",14558 => "11110001",14559 => "00101011",14560 => "11010010",14561 => "00010100",14562 => "00010010",14563 => "01100101",14564 => "10001110",14565 => "00011000",14566 => "00100101",14567 => "00111110",14568 => "10111000",14569 => "00101001",14570 => "10101010",14571 => "11010110",14572 => "01000010",14573 => "11001001",14574 => "10111110",14575 => "10001100",14576 => "01000010",14577 => "11011100",14578 => "11010001",14579 => "01110011",14580 => "10001100",14581 => "10001001",14582 => "10101010",14583 => "01000100",14584 => "01111000",14585 => "11100000",14586 => "11101010",14587 => "01110101",14588 => "01100110",14589 => "00111010",14590 => "00011001",14591 => "11111110",14592 => "11101000",14593 => "00001101",14594 => "00110110",14595 => "01010001",14596 => "01001010",14597 => "11000100",14598 => "10110100",14599 => "11110000",14600 => "11100011",14601 => "01111010",14602 => "10010000",14603 => "01111100",14604 => "01010111",14605 => "01001100",14606 => "11001001",14607 => "11111110",14608 => "00000100",14609 => "10010001",14610 => "11110101",14611 => "01100001",14612 => "10000011",14613 => "11001011",14614 => "11100110",14615 => "00100101",14616 => "01000101",14617 => "00111110",14618 => "11001011",14619 => "01011111",14620 => "10111001",14621 => "11000111",14622 => "11101001",14623 => "00001010",14624 => "11110100",14625 => "11011100",14626 => "11100111",14627 => "01111111",14628 => "00011110",14629 => "00011000",14630 => "10010111",14631 => "11101011",14632 => "10110101",14633 => "01010011",14634 => "10101011",14635 => "01010101",14636 => "00100101",14637 => "01001110",14638 => "00010000",14639 => "00000111",14640 => "01010101",14641 => "00001010",14642 => "10101110",14643 => "10001111",14644 => "10101110",14645 => "00010000",14646 => "11000001",14647 => "10110011",14648 => "11011111",14649 => "11111111",14650 => "11000011",14651 => "01111100",14652 => "10101000",14653 => "10110110",14654 => "11111110",14655 => "01110110",14656 => "10010000",14657 => "00000101",14658 => "00010010",14659 => "00100110",14660 => "11101001",14661 => "11101010",14662 => "00001100",14663 => "00000111",14664 => "00111110",14665 => "10111010",14666 => "10010111",14667 => "01101010",14668 => "01011010",14669 => "01000110",14670 => "00001000",14671 => "10101011",14672 => "00111101",14673 => "00111100",14674 => "01100001",14675 => "01010111",14676 => "10011001",14677 => "01101100",14678 => "00001001",14679 => "10010100",14680 => "01000000",14681 => "00000111",14682 => "11010101",14683 => "10101100",14684 => "00110111",14685 => "01100001",14686 => "11011111",14687 => "01111100",14688 => "00011011",14689 => "00110001",14690 => "00100010",14691 => "10001101",14692 => "11001010",14693 => "00101111",14694 => "00001111",14695 => "10000100",14696 => "10001100",14697 => "00001000",14698 => "01110100",14699 => "01011000",14700 => "10000111",14701 => "11001010",14702 => "00010010",14703 => "10101110",14704 => "01011011",14705 => "10010110",14706 => "00111001",14707 => "00110011",14708 => "00101110",14709 => "01010000",14710 => "01010010",14711 => "01010111",14712 => "00011100",14713 => "11110100",14714 => "11111110",14715 => "01101011",14716 => "10010101",14717 => "10100011",14718 => "00010011",14719 => "01110010",14720 => "10110000",14721 => "11010000",14722 => "10000100",14723 => "01011010",14724 => "00111101",14725 => "01010011",14726 => "01010001",14727 => "01010001",14728 => "01000101",14729 => "01100010",14730 => "00010101",14731 => "10011101",14732 => "10010111",14733 => "01111000",14734 => "01011101",14735 => "11101101",14736 => "10011001",14737 => "10100111",14738 => "01011011",14739 => "11101000",14740 => "10111100",14741 => "11011111",14742 => "10101110",14743 => "01011111",14744 => "10101001",14745 => "11100001",14746 => "11100011",14747 => "11111100",14748 => "11000000",14749 => "10100100",14750 => "11011011",14751 => "01101001",14752 => "00000010",14753 => "01111001",14754 => "11000100",14755 => "11111000",14756 => "00101001",14757 => "00111010",14758 => "01111111",14759 => "00100100",14760 => "00011100",14761 => "01001011",14762 => "00110110",14763 => "00100100",14764 => "00011110",14765 => "10001001",14766 => "01100110",14767 => "10100011",14768 => "11110011",14769 => "00010011",14770 => "00100011",14771 => "01101101",14772 => "11001001",14773 => "01101111",14774 => "00111111",14775 => "01011110",14776 => "10111111",14777 => "01100000",14778 => "10101111",14779 => "01111010",14780 => "01101100",14781 => "01101110",14782 => "01011001",14783 => "11110000",14784 => "01000011",14785 => "00001111",14786 => "00000000",14787 => "11001001",14788 => "10110001",14789 => "01000111",14790 => "00010110",14791 => "01100011",14792 => "00110101",14793 => "01010000",14794 => "01011111",14795 => "01110011",14796 => "11000011",14797 => "01011011",14798 => "10100111",14799 => "10111000",14800 => "01100101",14801 => "11110011",14802 => "11010011",14803 => "10111100",14804 => "10111010",14805 => "11111110",14806 => "10010110",14807 => "10101000",14808 => "01001100",14809 => "01000001",14810 => "00111010",14811 => "01010000",14812 => "00010001",14813 => "10100101",14814 => "11101000",14815 => "00100000",14816 => "00100000",14817 => "11110011",14818 => "01110011",14819 => "10011001",14820 => "11100000",14821 => "10000001",14822 => "10010010",14823 => "01001010",14824 => "11110001",14825 => "01111000",14826 => "00100011",14827 => "10101110",14828 => "10110011",14829 => "11110001",14830 => "11100001",14831 => "01000100",14832 => "11001000",14833 => "01101011",14834 => "01000011",14835 => "00100000",14836 => "11011001",14837 => "11101010",14838 => "10000001",14839 => "11100001",14840 => "10100000",14841 => "10000111",14842 => "01001100",14843 => "00111000",14844 => "00000101",14845 => "01010010",14846 => "00101111",14847 => "11110001",14848 => "10000000",14849 => "10001101",14850 => "00111010",14851 => "10011100",14852 => "01011011",14853 => "01110010",14854 => "01000110",14855 => "01001000",14856 => "01110001",14857 => "00011000",14858 => "11000000",14859 => "11001110",14860 => "10010110",14861 => "01100111",14862 => "11101001",14863 => "10110011",14864 => "11101111",14865 => "00001100",14866 => "11011011",14867 => "10001000",14868 => "11001000",14869 => "01001111",14870 => "11110111",14871 => "10110100",14872 => "00001100",14873 => "00011111",14874 => "00101111",14875 => "00100100",14876 => "01111110",14877 => "00100010",14878 => "10000000",14879 => "10111100",14880 => "11000101",14881 => "00010110",14882 => "10110011",14883 => "00111010",14884 => "01111001",14885 => "01010101",14886 => "01111110",14887 => "11101101",14888 => "11000110",14889 => "00101101",14890 => "10011010",14891 => "10010001",14892 => "10011010",14893 => "10100100",14894 => "11100001",14895 => "00100001",14896 => "10111001",14897 => "00000010",14898 => "11001010",14899 => "01101110",14900 => "11000001",14901 => "00011011",14902 => "11000101",14903 => "10011100",14904 => "10000000",14905 => "00101010",14906 => "01010000",14907 => "11000101",14908 => "00100011",14909 => "11010011",14910 => "11000010",14911 => "11111111",14912 => "01001110",14913 => "10101110",14914 => "00001010",14915 => "00010110",14916 => "10110000",14917 => "00000011",14918 => "11000011",14919 => "01010001",14920 => "00000101",14921 => "00001001",14922 => "11111001",14923 => "10011000",14924 => "10010001",14925 => "11010010",14926 => "00010100",14927 => "11110011",14928 => "11100100",14929 => "11111011",14930 => "00101010",14931 => "10001111",14932 => "00101100",14933 => "10111100",14934 => "00100110",14935 => "11100011",14936 => "10001110",14937 => "01110011",14938 => "01100011",14939 => "01101010",14940 => "00100000",14941 => "11001101",14942 => "11010100",14943 => "01000000",14944 => "00110001",14945 => "00011000",14946 => "01100001",14947 => "11111011",14948 => "01110101",14949 => "11111010",14950 => "00100110",14951 => "00000111",14952 => "10000001",14953 => "01100001",14954 => "01101000",14955 => "01011101",14956 => "00010010",14957 => "01101001",14958 => "11100110",14959 => "11001110",14960 => "01001110",14961 => "11110000",14962 => "11001011",14963 => "01001001",14964 => "00100101",14965 => "10000110",14966 => "11110000",14967 => "01011011",14968 => "01001000",14969 => "01111110",14970 => "11011011",14971 => "10111110",14972 => "10101110",14973 => "10011111",14974 => "00100110",14975 => "00110010",14976 => "10100011",14977 => "01000001",14978 => "11110111",14979 => "11100110",14980 => "11111100",14981 => "01011001",14982 => "11110101",14983 => "00000011",14984 => "01111011",14985 => "00100010",14986 => "00101001",14987 => "10010010",14988 => "01100111",14989 => "01000010",14990 => "01000111",14991 => "10010000",14992 => "01001100",14993 => "10000100",14994 => "10001101",14995 => "01011001",14996 => "11010001",14997 => "10000100",14998 => "00101010",14999 => "10000110",15000 => "00110101",15001 => "01100101",15002 => "00100100",15003 => "11000010",15004 => "00000101",15005 => "01101110",15006 => "11010101",15007 => "01111010",15008 => "11100101",15009 => "00111100",15010 => "11100000",15011 => "00100000",15012 => "11100000",15013 => "11000110",15014 => "01110010",15015 => "11100011",15016 => "01010010",15017 => "10001110",15018 => "00011110",15019 => "01011000",15020 => "00011111",15021 => "10001100",15022 => "01101100",15023 => "10110000",15024 => "00111110",15025 => "00100010",15026 => "11000100",15027 => "01000100",15028 => "01010000",15029 => "01111010",15030 => "01101001",15031 => "01011100",15032 => "01001011",15033 => "01000011",15034 => "11110011",15035 => "00010001",15036 => "01011010",15037 => "10111011",15038 => "10111001",15039 => "10011101",15040 => "01001111",15041 => "00010001",15042 => "11110101",15043 => "01000011",15044 => "00010100",15045 => "11100010",15046 => "11000111",15047 => "11000011",15048 => "01000011",15049 => "11111010",15050 => "11101111",15051 => "10111001",15052 => "01110101",15053 => "10100111",15054 => "10110100",15055 => "01100010",15056 => "00111010",15057 => "10111011",15058 => "11101000",15059 => "01111000",15060 => "00000010",15061 => "10001111",15062 => "00011010",15063 => "01001111",15064 => "10110100",15065 => "00010011",15066 => "10111010",15067 => "11100000",15068 => "01101011",15069 => "01001100",15070 => "10011010",15071 => "11011011",15072 => "01100110",15073 => "01101011",15074 => "01111011",15075 => "01110100",15076 => "10011001",15077 => "11001100",15078 => "00010000",15079 => "00010111",15080 => "10011101",15081 => "01100010",15082 => "01000111",15083 => "00010010",15084 => "11100110",15085 => "01000110",15086 => "00001011",15087 => "01111001",15088 => "10000001",15089 => "11010000",15090 => "10000111",15091 => "00011001",15092 => "10001101",15093 => "11110000",15094 => "10000000",15095 => "00000010",15096 => "10101001",15097 => "00101111",15098 => "11010101",15099 => "11001100",15100 => "01110010",15101 => "01110101",15102 => "10010111",15103 => "10001101",15104 => "00010000",15105 => "01100011",15106 => "11001001",15107 => "01011110",15108 => "11101100",15109 => "11000011",15110 => "00000110",15111 => "11111011",15112 => "00010001",15113 => "00110011",15114 => "00110000",15115 => "10011010",15116 => "01111101",15117 => "10010001",15118 => "11000100",15119 => "00011000",15120 => "01010111",15121 => "10101111",15122 => "00011011",15123 => "10100010",15124 => "01111100",15125 => "10011101",15126 => "11010101",15127 => "00000110",15128 => "10010101",15129 => "01110110",15130 => "11110101",15131 => "11111110",15132 => "01110011",15133 => "11000111",15134 => "10110111",15135 => "11111011",15136 => "10100001",15137 => "11000001",15138 => "00000101",15139 => "11110011",15140 => "00101001",15141 => "10001001",15142 => "11100101",15143 => "11100000",15144 => "10100000",15145 => "00011001",15146 => "00100000",15147 => "01011100",15148 => "11101100",15149 => "11001111",15150 => "00110010",15151 => "00010111",15152 => "01001010",15153 => "11011010",15154 => "11100111",15155 => "01011110",15156 => "00010110",15157 => "10001110",15158 => "01001001",15159 => "00111000",15160 => "11000101",15161 => "10101001",15162 => "10000111",15163 => "10100101",15164 => "01101100",15165 => "00010000",15166 => "00000111",15167 => "11011100",15168 => "00101101",15169 => "10010000",15170 => "00101000",15171 => "11110001",15172 => "01001000",15173 => "01101100",15174 => "01011001",15175 => "00101011",15176 => "00110000",15177 => "00110111",15178 => "01001100",15179 => "11000011",15180 => "00101111",15181 => "11110000",15182 => "10011101",15183 => "00000000",15184 => "01101000",15185 => "00010011",15186 => "11000101",15187 => "00101101",15188 => "01111110",15189 => "00001110",15190 => "11101000",15191 => "11110011",15192 => "10100111",15193 => "01101111",15194 => "11111011",15195 => "01100100",15196 => "11001111",15197 => "01001010",15198 => "00000011",15199 => "00000011",15200 => "00110101",15201 => "01001101",15202 => "10000110",15203 => "10101010",15204 => "11010000",15205 => "00111000",15206 => "11001111",15207 => "01100011",15208 => "01111010",15209 => "00000111",15210 => "11101001",15211 => "01100110",15212 => "01001010",15213 => "00000100",15214 => "01101001",15215 => "10010011",15216 => "01010001",15217 => "01000010",15218 => "00101000",15219 => "11011011",15220 => "00000101",15221 => "11100000",15222 => "01100110",15223 => "01110101",15224 => "10111101",15225 => "01111111",15226 => "00000001",15227 => "11100001",15228 => "11000110",15229 => "00100010",15230 => "00101010",15231 => "10010010",15232 => "01000110",15233 => "10001010",15234 => "00001101",15235 => "00110100",15236 => "11111111",15237 => "01000010",15238 => "11001110",15239 => "00010110",15240 => "01011101",15241 => "11011011",15242 => "01111110",15243 => "10000011",15244 => "00011011",15245 => "01010011",15246 => "00101111",15247 => "11010000",15248 => "11100001",15249 => "00010100",15250 => "10101011",15251 => "11110010",15252 => "10000110",15253 => "00110100",15254 => "00110000",15255 => "11000001",15256 => "10001101",15257 => "11110000",15258 => "01101111",15259 => "01011010",15260 => "01110101",15261 => "10111010",15262 => "00100101",15263 => "00001101",15264 => "01110110",15265 => "11001000",15266 => "01000100",15267 => "10000011",15268 => "00110111",15269 => "11111000",15270 => "10101111",15271 => "10000111",15272 => "11101000",15273 => "11001111",15274 => "10011101",15275 => "01010001",15276 => "01010011",15277 => "10110100",15278 => "01111001",15279 => "01011101",15280 => "10011010",15281 => "00011101",15282 => "01001110",15283 => "10110010",15284 => "10010010",15285 => "10111010",15286 => "00111100",15287 => "11111010",15288 => "11010101",15289 => "10001111",15290 => "11011111",15291 => "11110000",15292 => "10000000",15293 => "10111011",15294 => "11110010",15295 => "11100110",15296 => "10100101",15297 => "11111001",15298 => "01010010",15299 => "10100110",15300 => "01000100",15301 => "01011001",15302 => "00011101",15303 => "10100001",15304 => "11101101",15305 => "10010010",15306 => "11101101",15307 => "01000101",15308 => "00111000",15309 => "00110110",15310 => "10000110",15311 => "11111100",15312 => "01101110",15313 => "01011110",15314 => "00100001",15315 => "00001100",15316 => "10011111",15317 => "10001011",15318 => "11100110",15319 => "01110001",15320 => "11001111",15321 => "00011000",15322 => "10101000",15323 => "01101100",15324 => "00100100",15325 => "11110011",15326 => "01111100",15327 => "00000100",15328 => "00110011",15329 => "10000110",15330 => "10101100",15331 => "00011000",15332 => "10110100",15333 => "10110111",15334 => "01010110",15335 => "00011111",15336 => "00011100",15337 => "00100011",15338 => "00111000",15339 => "00110110",15340 => "01011000",15341 => "10001000",15342 => "11000000",15343 => "10101011",15344 => "01111100",15345 => "01011100",15346 => "10101111",15347 => "01110100",15348 => "11110011",15349 => "00111101",15350 => "00101010",15351 => "01101100",15352 => "00011011",15353 => "10110000",15354 => "11111010",15355 => "10101100",15356 => "10110001",15357 => "10011000",15358 => "10111111",15359 => "01010000",15360 => "01011101",15361 => "00010100",15362 => "01000110",15363 => "10110000",15364 => "10000000",15365 => "01111101",15366 => "11100101",15367 => "11010110",15368 => "11010111",15369 => "00001100",15370 => "00000010",15371 => "01100110",15372 => "10100010",15373 => "00010110",15374 => "00101111",15375 => "10100010",15376 => "10100110",15377 => "00100111",15378 => "10111010",15379 => "00011010",15380 => "11111011",15381 => "01000110",15382 => "01000011",15383 => "01111111",15384 => "01101111",15385 => "10111011",15386 => "10101010",15387 => "00011100",15388 => "10010101",15389 => "01000011",15390 => "01110111",15391 => "10001010",15392 => "00101100",15393 => "11111101",15394 => "00111001",15395 => "00001011",15396 => "00100111",15397 => "10101011",15398 => "11111101",15399 => "10010000",15400 => "00100110",15401 => "10101000",15402 => "01000101",15403 => "11000010",15404 => "11110111",15405 => "00010001",15406 => "00110101",15407 => "01000010",15408 => "10010011",15409 => "00110001",15410 => "01000111",15411 => "00000101",15412 => "01100100",15413 => "01000110",15414 => "01010101",15415 => "00010111",15416 => "11010110",15417 => "11110110",15418 => "01001101",15419 => "01101010",15420 => "11111000",15421 => "01000000",15422 => "00011001",15423 => "11101010",15424 => "00001111",15425 => "00001000",15426 => "01111111",15427 => "10000110",15428 => "10011101",15429 => "11101010",15430 => "01000111",15431 => "01100111",15432 => "11101000",15433 => "11101000",15434 => "11011100",15435 => "10101011",15436 => "10100110",15437 => "01101101",15438 => "10011011",15439 => "00110110",15440 => "00000000",15441 => "00110111",15442 => "11111101",15443 => "11110001",15444 => "10001011",15445 => "00010010",15446 => "00110110",15447 => "10001100",15448 => "01001111",15449 => "10110100",15450 => "10110001",15451 => "11011000",15452 => "11111111",15453 => "00101111",15454 => "00000100",15455 => "01000100",15456 => "11001110",15457 => "10101001",15458 => "11101011",15459 => "10110100",15460 => "00111100",15461 => "10101000",15462 => "01101010",15463 => "11100111",15464 => "00001111",15465 => "10010111",15466 => "11001001",15467 => "01001010",15468 => "11110011",15469 => "00100011",15470 => "01110111",15471 => "11001100",15472 => "01001111",15473 => "10110110",15474 => "11110000",15475 => "01110111",15476 => "11110110",15477 => "01010101",15478 => "00011010",15479 => "11001100",15480 => "00110001",15481 => "11100111",15482 => "00100111",15483 => "00010111",15484 => "11000010",15485 => "01010110",15486 => "00101110",15487 => "10000001",15488 => "00111001",15489 => "00001110",15490 => "01100111",15491 => "10111001",15492 => "11011011",15493 => "10010110",15494 => "11111000",15495 => "00011111",15496 => "01011000",15497 => "00011100",15498 => "01101111",15499 => "01100110",15500 => "10111111",15501 => "10000011",15502 => "10100100",15503 => "11001110",15504 => "01000111",15505 => "10011001",15506 => "11100001",15507 => "01011011",15508 => "00001101",15509 => "11000011",15510 => "10010001",15511 => "01010100",15512 => "00110011",15513 => "10111111",15514 => "10010001",15515 => "10100010",15516 => "11101110",15517 => "00001101",15518 => "00011001",15519 => "00111101",15520 => "10111100",15521 => "00001000",15522 => "11110110",15523 => "01000111",15524 => "11010011",15525 => "11010101",15526 => "10010110",15527 => "01000010",15528 => "00001000",15529 => "11111011",15530 => "00001110",15531 => "10001111",15532 => "10000101",15533 => "10100111",15534 => "11001101",15535 => "01010001",15536 => "11010110",15537 => "00101110",15538 => "00101000",15539 => "00001000",15540 => "00110100",15541 => "11111101",15542 => "00001100",15543 => "11111000",15544 => "10110101",15545 => "11010101",15546 => "01101011",15547 => "11010111",15548 => "10111001",15549 => "10011001",15550 => "01110111",15551 => "00101011",15552 => "11001001",15553 => "10100000",15554 => "00010000",15555 => "10000100",15556 => "10110010",15557 => "00011011",15558 => "01111101",15559 => "01000011",15560 => "01000000",15561 => "11010011",15562 => "01100000",15563 => "10000011",15564 => "01011110",15565 => "01100011",15566 => "11100100",15567 => "11100000",15568 => "01011000",15569 => "11000111",15570 => "01100001",15571 => "11101100",15572 => "01011110",15573 => "10011101",15574 => "11100100",15575 => "01110100",15576 => "11100011",15577 => "01110000",15578 => "00000001",15579 => "00010010",15580 => "00100011",15581 => "11100110",15582 => "00110011",15583 => "11100100",15584 => "01101101",15585 => "11000111",15586 => "10100011",15587 => "00111011",15588 => "10101110",15589 => "00001111",15590 => "01100010",15591 => "01100101",15592 => "00011110",15593 => "11111011",15594 => "10100000",15595 => "11110011",15596 => "00001000",15597 => "01001010",15598 => "00001110",15599 => "10010010",15600 => "00000101",15601 => "00110100",15602 => "00000011",15603 => "11101101",15604 => "11010001",15605 => "00000010",15606 => "11111110",15607 => "11100101",15608 => "10011100",15609 => "00010010",15610 => "00010111",15611 => "01111000",15612 => "10111111",15613 => "01100100",15614 => "00001100",15615 => "11001101",15616 => "00010111",15617 => "11111110",15618 => "00100100",15619 => "10101001",15620 => "00010010",15621 => "00000011",15622 => "01011011",15623 => "11110000",15624 => "10111101",15625 => "01011000",15626 => "10101111",15627 => "01111101",15628 => "01100100",15629 => "11111001",15630 => "01011010",15631 => "10011000",15632 => "00011011",15633 => "10110111",15634 => "10111110",15635 => "10110111",15636 => "01101100",15637 => "11101111",15638 => "11110001",15639 => "10010001",15640 => "01101111",15641 => "00101111",15642 => "10011000",15643 => "11111111",15644 => "10101111",15645 => "01110011",15646 => "00110010",15647 => "01011010",15648 => "00010100",15649 => "10111010",15650 => "11001111",15651 => "10001000",15652 => "11010010",15653 => "10001010",15654 => "10010111",15655 => "11110100",15656 => "01111110",15657 => "10001101",15658 => "00110101",15659 => "10001010",15660 => "11001110",15661 => "10111001",15662 => "01000110",15663 => "11100111",15664 => "01111111",15665 => "10001010",15666 => "10101110",15667 => "11010110",15668 => "01101011",15669 => "10010101",15670 => "11110110",15671 => "11110011",15672 => "11011001",15673 => "10110011",15674 => "01001011",15675 => "11110000",15676 => "10111001",15677 => "00100110",15678 => "10000100",15679 => "00011001",15680 => "00100100",15681 => "01110110",15682 => "10011001",15683 => "01100000",15684 => "10101111",15685 => "10101001",15686 => "01101001",15687 => "00111000",15688 => "00000010",15689 => "01010111",15690 => "00101001",15691 => "01111100",15692 => "10010100",15693 => "10110010",15694 => "01001110",15695 => "11110000",15696 => "00011101",15697 => "00011010",15698 => "11111010",15699 => "00010000",15700 => "10011100",15701 => "01001001",15702 => "11110101",15703 => "10101001",15704 => "11111111",15705 => "11110011",15706 => "00000000",15707 => "01001101",15708 => "01010000",15709 => "11001101",15710 => "10010101",15711 => "10111010",15712 => "01100000",15713 => "00101111",15714 => "10001000",15715 => "10111011",15716 => "01010010",15717 => "11100101",15718 => "10001011",15719 => "01110001",15720 => "10011011",15721 => "10001010",15722 => "00111010",15723 => "11100101",15724 => "11010111",15725 => "00110011",15726 => "10011100",15727 => "01111111",15728 => "10000001",15729 => "11111110",15730 => "01110000",15731 => "01001100",15732 => "10010010",15733 => "01110001",15734 => "01111111",15735 => "00001010",15736 => "11010100",15737 => "00011111",15738 => "10001110",15739 => "10100011",15740 => "10000111",15741 => "01010011",15742 => "10110011",15743 => "10000100",15744 => "01010001",15745 => "01001111",15746 => "00010111",15747 => "00001110",15748 => "10001010",15749 => "00110110",15750 => "11100010",15751 => "00101010",15752 => "00010000",15753 => "10100011",15754 => "01100110",15755 => "11111011",15756 => "00001101",15757 => "01000001",15758 => "11111000",15759 => "11000001",15760 => "01011001",15761 => "11100001",15762 => "10001111",15763 => "10111000",15764 => "11000010",15765 => "10110111",15766 => "00000111",15767 => "11100101",15768 => "01110010",15769 => "11110000",15770 => "01111111",15771 => "10110000",15772 => "11110000",15773 => "10010111",15774 => "01001111",15775 => "10101011",15776 => "11111101",15777 => "00010101",15778 => "11011001",15779 => "10101001",15780 => "01111010",15781 => "01101011",15782 => "00101000",15783 => "10101010",15784 => "00001010",15785 => "01011101",15786 => "00101110",15787 => "01011011",15788 => "10110000",15789 => "01101100",15790 => "01000001",15791 => "10010011",15792 => "01010000",15793 => "10010100",15794 => "10010111",15795 => "11100101",15796 => "10010011",15797 => "11100011",15798 => "11001001",15799 => "01111000",15800 => "11000001",15801 => "00010111",15802 => "01100010",15803 => "01110110",15804 => "00001110",15805 => "10100001",15806 => "11111001",15807 => "11001111",15808 => "01011100",15809 => "00010111",15810 => "01010011",15811 => "01110100",15812 => "11101001",15813 => "11111110",15814 => "00101011",15815 => "00010001",15816 => "10000111",15817 => "01001101",15818 => "10110010",15819 => "10101110",15820 => "11101000",15821 => "00001111",15822 => "10001110",15823 => "00011101",15824 => "11110111",15825 => "11011111",15826 => "10101110",15827 => "01101110",15828 => "01111001",15829 => "11000010",15830 => "11010111",15831 => "10100010",15832 => "11111111",15833 => "11100111",15834 => "00110111",15835 => "01101100",15836 => "00111001",15837 => "10111101",15838 => "00000101",15839 => "00110101",15840 => "10000000",15841 => "11110001",15842 => "11101001",15843 => "01110111",15844 => "10110001",15845 => "10101010",15846 => "10101100",15847 => "10101111",15848 => "11011111",15849 => "01110100",15850 => "10110100",15851 => "01100101",15852 => "10101111",15853 => "10001111",15854 => "01110110",15855 => "11010010",15856 => "01010010",15857 => "10001001",15858 => "00011000",15859 => "00001001",15860 => "10111110",15861 => "11001011",15862 => "00011101",15863 => "10001000",15864 => "10110110",15865 => "10000101",15866 => "00100011",15867 => "10001010",15868 => "10111100",15869 => "00011000",15870 => "10111100",15871 => "01100110",15872 => "00111001",15873 => "01011111",15874 => "10111011",15875 => "01101100",15876 => "11101110",15877 => "00010001",15878 => "11111100",15879 => "01001000",15880 => "10010110",15881 => "10101110",15882 => "01111101",15883 => "00000010",15884 => "10110100",15885 => "01100100",15886 => "10000111",15887 => "01001100",15888 => "01111100",15889 => "11100000",15890 => "01001001",15891 => "01101000",15892 => "00011110",15893 => "11011100",15894 => "00000011",15895 => "11100110",15896 => "00010100",15897 => "11111111",15898 => "00010101",15899 => "11000101",15900 => "00011100",15901 => "11100011",15902 => "10100000",15903 => "01011100",15904 => "00110111",15905 => "11000001",15906 => "10111101",15907 => "10100000",15908 => "01000010",15909 => "11101110",15910 => "11100000",15911 => "01011111",15912 => "00000011",15913 => "10110100",15914 => "01001010",15915 => "00110011",15916 => "01101111",15917 => "11011001",15918 => "11111101",15919 => "10000001",15920 => "00110001",15921 => "01001111",15922 => "11110101",15923 => "01011110",15924 => "10000110",15925 => "11101100",15926 => "11010011",15927 => "00100011",15928 => "00011111",15929 => "10110100",15930 => "01100000",15931 => "00011110",15932 => "11011110",15933 => "10100000",15934 => "01000011",15935 => "10100001",15936 => "01010011",15937 => "10010010",15938 => "00011010",15939 => "10111011",15940 => "11001110",15941 => "11101111",15942 => "01011100",15943 => "00100000",15944 => "10110010",15945 => "01101101",15946 => "10100001",15947 => "11100111",15948 => "11100111",15949 => "11010010",15950 => "01011111",15951 => "00110100",15952 => "11110000",15953 => "11011100",15954 => "10010010",15955 => "01011110",15956 => "00000010",15957 => "11100100",15958 => "10010001",15959 => "10100011",15960 => "00010011",15961 => "01100111",15962 => "01111011",15963 => "01101100",15964 => "10011010",15965 => "00101011",15966 => "01101100",15967 => "10011001",15968 => "00000010",15969 => "01011000",15970 => "00011111",15971 => "11010110",15972 => "10101000",15973 => "01001111",15974 => "00000100",15975 => "00000001",15976 => "10101001",15977 => "00100011",15978 => "01010101",15979 => "01000111",15980 => "11111111",15981 => "11110001",15982 => "11110111",15983 => "11000111",15984 => "00000100",15985 => "11100011",15986 => "00001100",15987 => "11010011",15988 => "00111111",15989 => "00011011",15990 => "11100010",15991 => "00001111",15992 => "00001001",15993 => "01011110",15994 => "01011011",15995 => "00011001",15996 => "00010010",15997 => "11001000",15998 => "00000010",15999 => "10111101",16000 => "10001101",16001 => "11111111",16002 => "11010011",16003 => "00110100",16004 => "11111111",16005 => "01101011",16006 => "10110111",16007 => "11000110",16008 => "01101111",16009 => "01110011",16010 => "11101011",16011 => "00011100",16012 => "01101100",16013 => "01100010",16014 => "00011010",16015 => "00010011",16016 => "10000100",16017 => "01011111",16018 => "01101111",16019 => "00110001",16020 => "01001001",16021 => "11001100",16022 => "01001001",16023 => "10110001",16024 => "10101101",16025 => "01101101",16026 => "00001010",16027 => "01111110",16028 => "01010011",16029 => "01100001",16030 => "00111000",16031 => "10101000",16032 => "10011001",16033 => "01100110",16034 => "10100111",16035 => "01010000",16036 => "00110100",16037 => "10000010",16038 => "10011001",16039 => "00000100",16040 => "11101100",16041 => "01111010",16042 => "10001101",16043 => "11010000",16044 => "10000100",16045 => "00100001",16046 => "01101110",16047 => "10000010",16048 => "00010010",16049 => "00110110",16050 => "01100110",16051 => "01001100",16052 => "10001101",16053 => "01111011",16054 => "10111110",16055 => "00100110",16056 => "11101011",16057 => "10101101",16058 => "11010100",16059 => "00011110",16060 => "11101010",16061 => "11110111",16062 => "01011001",16063 => "10000111",16064 => "01100111",16065 => "11001110",16066 => "01110000",16067 => "11000011",16068 => "10111110",16069 => "00001001",16070 => "11000111",16071 => "01110010",16072 => "11110010",16073 => "10000111",16074 => "00111001",16075 => "10110110",16076 => "11000101",16077 => "11000100",16078 => "11011111",16079 => "01100111",16080 => "01111000",16081 => "11000010",16082 => "10110001",16083 => "10011100",16084 => "10111101",16085 => "11100010",16086 => "00011100",16087 => "00111111",16088 => "10101001",16089 => "10101110",16090 => "01000110",16091 => "11000110",16092 => "10110010",16093 => "01110111",16094 => "01000110",16095 => "01010010",16096 => "01101101",16097 => "10110001",16098 => "00111011",16099 => "01000010",16100 => "01111011",16101 => "00000011",16102 => "01111111",16103 => "11100111",16104 => "11100111",16105 => "00001100",16106 => "00010101",16107 => "01101100",16108 => "11111111",16109 => "11011100",16110 => "11010111",16111 => "00011001",16112 => "11010100",16113 => "01111100",16114 => "11011101",16115 => "00111111",16116 => "10010101",16117 => "11110100",16118 => "00110000",16119 => "11011010",16120 => "00000011",16121 => "01101100",16122 => "00001110",16123 => "00000011",16124 => "01110000",16125 => "01000001",16126 => "10101000",16127 => "11111111",16128 => "01101001",16129 => "01100110",16130 => "01001101",16131 => "11100001",16132 => "01001101",16133 => "01111000",16134 => "00011001",16135 => "11101010",16136 => "00000000",16137 => "01100100",16138 => "01011000",16139 => "01110011",16140 => "00000110",16141 => "11011110",16142 => "01011011",16143 => "01000111",16144 => "10010000",16145 => "11001001",16146 => "00100100",16147 => "01111010",16148 => "00100010",16149 => "10100011",16150 => "00100011",16151 => "11111110",16152 => "11111111",16153 => "10000100",16154 => "10001010",16155 => "00111111",16156 => "01101011",16157 => "01110000",16158 => "00000101",16159 => "11101100",16160 => "01000010",16161 => "00110100",16162 => "11010000",16163 => "11001000",16164 => "10110011",16165 => "10000001",16166 => "10011000",16167 => "11111101",16168 => "01000101",16169 => "00110101",16170 => "11101111",16171 => "10011110",16172 => "10110010",16173 => "00101100",16174 => "11101111",16175 => "00101001",16176 => "01101010",16177 => "01101001",16178 => "10100001",16179 => "00010000",16180 => "10110010",16181 => "11111000",16182 => "10110011",16183 => "11001101",16184 => "11001001",16185 => "10001010",16186 => "00101011",16187 => "01100110",16188 => "11000011",16189 => "00011011",16190 => "00011011",16191 => "10111001",16192 => "11001010",16193 => "11011110",16194 => "11000110",16195 => "01010001",16196 => "01101110",16197 => "11011110",16198 => "10010010",16199 => "11010100",16200 => "00110110",16201 => "01011011",16202 => "10011010",16203 => "01101110",16204 => "11011110",16205 => "00100101",16206 => "00101111",16207 => "00000101",16208 => "11001011",16209 => "00111100",16210 => "01100010",16211 => "11100000",16212 => "11010101",16213 => "00000011",16214 => "01011010",16215 => "11001100",16216 => "00100011",16217 => "11011010",16218 => "00100011",16219 => "11110010",16220 => "01011101",16221 => "00110001",16222 => "11111000",16223 => "11110001",16224 => "00001101",16225 => "10100000",16226 => "11001100",16227 => "11110010",16228 => "00100110",16229 => "11001011",16230 => "00001101",16231 => "01001101",16232 => "11011010",16233 => "01100111",16234 => "11110000",16235 => "01001010",16236 => "10011101",16237 => "00000010",16238 => "10111100",16239 => "10011011",16240 => "11000100",16241 => "11100000",16242 => "00011100",16243 => "11000010",16244 => "00011010",16245 => "10110111",16246 => "11110111",16247 => "11111101",16248 => "11111000",16249 => "10010101",16250 => "11010101",16251 => "01110011",16252 => "11010110",16253 => "00010111",16254 => "10010011",16255 => "01011101",16256 => "00111000",16257 => "00101111",16258 => "01110011",16259 => "10011011",16260 => "10010010",16261 => "11000101",16262 => "00110011",16263 => "11001001",16264 => "00000000",16265 => "10101101",16266 => "11100001",16267 => "01000110",16268 => "01101011",16269 => "00000110",16270 => "01000111",16271 => "00011000",16272 => "10010001",16273 => "01000000",16274 => "00111101",16275 => "10111111",16276 => "10010010",16277 => "01100101",16278 => "11111100",16279 => "11010110",16280 => "10110001",16281 => "10010101",16282 => "11000011",16283 => "11000101",16284 => "01011010",16285 => "01101110",16286 => "11110010",16287 => "01101001",16288 => "00000010",16289 => "01100001",16290 => "11101101",16291 => "11101100",16292 => "11101011",16293 => "11011011",16294 => "11100001",16295 => "01110011",16296 => "10100100",16297 => "10001101",16298 => "11011000",16299 => "00011000",16300 => "10111111",16301 => "10110100",16302 => "00000011",16303 => "11000001",16304 => "01001101",16305 => "10001100",16306 => "10001111",16307 => "11010110",16308 => "11100000",16309 => "00101011",16310 => "10000111",16311 => "11000001",16312 => "10111011",16313 => "01101101",16314 => "10000101",16315 => "11000000",16316 => "00010101",16317 => "01101000",16318 => "01010011",16319 => "01110100",16320 => "00000100",16321 => "10101011",16322 => "00111000",16323 => "11001101",16324 => "00100100",16325 => "00110001",16326 => "01111010",16327 => "10100010",16328 => "00001011",16329 => "00111111",16330 => "11011001",16331 => "11101111",16332 => "00101000",16333 => "00011110",16334 => "01010110",16335 => "00100110",16336 => "01111000",16337 => "11110010",16338 => "11101111",16339 => "01000010",16340 => "00100001",16341 => "10111010",16342 => "00110010",16343 => "11101010",16344 => "01010010",16345 => "01111100",16346 => "01111000",16347 => "00111001",16348 => "10000001",16349 => "10000001",16350 => "01000001",16351 => "10010111",16352 => "00010000",16353 => "11101100",16354 => "11101110",16355 => "10110010",16356 => "01111110",16357 => "10000001",16358 => "01000111",16359 => "00001110",16360 => "00001100",16361 => "00011101",16362 => "00101111",16363 => "01011000",16364 => "00011001",16365 => "00110000",16366 => "01000100",16367 => "10011000",16368 => "01001001",16369 => "00011011",16370 => "11010110",16371 => "01010011",16372 => "01100111",16373 => "00000011",16374 => "10111101",16375 => "11011000",16376 => "01001010",16377 => "11010000",16378 => "01100000",16379 => "10011010",16380 => "01110110",16381 => "00101100",16382 => "01111011",16383 => "00110001",16384 => "10010010",16385 => "01101000",16386 => "00111010",16387 => "00000000",16388 => "01111111",16389 => "10101001",16390 => "10011111",16391 => "00000101",16392 => "01011001",16393 => "11101111",16394 => "10000001",16395 => "00111111",16396 => "10101001",16397 => "10011001",16398 => "11101010",16399 => "11010011",16400 => "10011101",16401 => "00010111",16402 => "01011010",16403 => "00000000",16404 => "11011111",16405 => "10010001",16406 => "11111111",16407 => "11111000",16408 => "00000110",16409 => "00100100",16410 => "10100000",16411 => "00101111",16412 => "01001111",16413 => "10010000",16414 => "00100011",16415 => "11001000",16416 => "10110100",16417 => "00010110",16418 => "11100100",16419 => "11101011",16420 => "00010010",16421 => "10011011",16422 => "11101111",16423 => "01001101",16424 => "00100111",16425 => "00110110",16426 => "00001001",16427 => "10010101",16428 => "01111010",16429 => "10101001",16430 => "11110110",16431 => "10100100",16432 => "10101110",16433 => "11011001",16434 => "00001010",16435 => "01001111",16436 => "00001100",16437 => "11001110",16438 => "11010111",16439 => "00100111",16440 => "00010001",16441 => "01011100",16442 => "10010010",16443 => "01011011",16444 => "01101000",16445 => "11101000",16446 => "10110100",16447 => "01101001",16448 => "00100000",16449 => "01101011",16450 => "11110100",16451 => "01000000",16452 => "11011100",16453 => "00010000",16454 => "10110101",16455 => "00100011",16456 => "11011000",16457 => "01000001",16458 => "01101101",16459 => "01111011",16460 => "00100100",16461 => "10100101",16462 => "10111110",16463 => "01000110",16464 => "01000001",16465 => "11011111",16466 => "10101010",16467 => "10100100",16468 => "10000000",16469 => "01111001",16470 => "11000110",16471 => "11000111",16472 => "00000000",16473 => "10111011",16474 => "11101100",16475 => "10000000",16476 => "00111001",16477 => "11001011",16478 => "11111001",16479 => "11110011",16480 => "00111100",16481 => "11001101",16482 => "11000001",16483 => "00111011",16484 => "01110011",16485 => "11111101",16486 => "11010110",16487 => "10100000",16488 => "11111101",16489 => "10100101",16490 => "00111011",16491 => "01000010",16492 => "00011110",16493 => "11010110",16494 => "01000000",16495 => "10100110",16496 => "00001010",16497 => "10110101",16498 => "01110001",16499 => "11110111",16500 => "00011111",16501 => "01101110",16502 => "00001011",16503 => "00011101",16504 => "01011100",16505 => "10000101",16506 => "01101101",16507 => "00000111",16508 => "00110111",16509 => "11001111",16510 => "01100100",16511 => "10010111",16512 => "11110010",16513 => "01010111",16514 => "00101000",16515 => "00010101",16516 => "00011011",16517 => "00111111",16518 => "00000111",16519 => "00111011",16520 => "00001010",16521 => "00101001",16522 => "11110000",16523 => "11011100",16524 => "00010011",16525 => "11000010",16526 => "00100011",16527 => "01000011",16528 => "00011110",16529 => "11010001",16530 => "01000011",16531 => "01111010",16532 => "10011000",16533 => "01101011",16534 => "01000010",16535 => "01010111",16536 => "10100100",16537 => "11110000",16538 => "00010011",16539 => "11001001",16540 => "11011111",16541 => "10010000",16542 => "01011010",16543 => "10110110",16544 => "01000110",16545 => "00100100",16546 => "11011111",16547 => "10111111",16548 => "11111010",16549 => "01100100",16550 => "11100000",16551 => "01110010",16552 => "00000110",16553 => "00000010",16554 => "10011101",16555 => "01010000",16556 => "01101111",16557 => "00100010",16558 => "00111011",16559 => "11011000",16560 => "10011100",16561 => "00000000",16562 => "11100000",16563 => "01001011",16564 => "10000110",16565 => "00100000",16566 => "10100010",16567 => "00011101",16568 => "11010001",16569 => "11000110",16570 => "11011101",16571 => "11100100",16572 => "11010000",16573 => "10111000",16574 => "11000110",16575 => "11111111",16576 => "01000100",16577 => "01011010",16578 => "01011010",16579 => "01000010",16580 => "10001001",16581 => "01101000",16582 => "10100101",16583 => "11101001",16584 => "01111100",16585 => "10011110",16586 => "10101101",16587 => "01000011",16588 => "11000111",16589 => "01011010",16590 => "00111111",16591 => "11111110",16592 => "11101011",16593 => "11010000",16594 => "01011011",16595 => "10101010",16596 => "01100101",16597 => "01010011",16598 => "10011110",16599 => "11100010",16600 => "01111010",16601 => "11101001",16602 => "10100110",16603 => "01111100",16604 => "11001110",16605 => "00100100",16606 => "11101111",16607 => "10000101",16608 => "00100010",16609 => "00110101",16610 => "10010011",16611 => "01000100",16612 => "10100110",16613 => "11101000",16614 => "00101000",16615 => "00000010",16616 => "10100111",16617 => "01111001",16618 => "10101110",16619 => "00010100",16620 => "00010010",16621 => "01111010",16622 => "00111111",16623 => "10100101",16624 => "00110110",16625 => "10000110",16626 => "01110110",16627 => "11100011",16628 => "11000110",16629 => "00111011",16630 => "11101001",16631 => "10100110",16632 => "00111000",16633 => "01000111",16634 => "00011111",16635 => "11000110",16636 => "01100001",16637 => "00000001",16638 => "10000000",16639 => "01101110",16640 => "00000001",16641 => "10111010",16642 => "10110100",16643 => "00001000",16644 => "11011000",16645 => "00000011",16646 => "10001111",16647 => "11110011",16648 => "11011000",16649 => "10110001",16650 => "11111000",16651 => "00110001",16652 => "01110111",16653 => "00110100",16654 => "11101001",16655 => "01000111",16656 => "00110001",16657 => "00111011",16658 => "01111100",16659 => "00100011",16660 => "11111110",16661 => "10110001",16662 => "10011111",16663 => "00011010",16664 => "01011110",16665 => "00010111",16666 => "01101111",16667 => "01010000",16668 => "11100010",16669 => "00111001",16670 => "11010110",16671 => "01111010",16672 => "00100011",16673 => "00010000",16674 => "00001011",16675 => "10101010",16676 => "10001111",16677 => "00100111",16678 => "00100111",16679 => "10011110",16680 => "11100111",16681 => "10001100",16682 => "00001010",16683 => "10011010",16684 => "11001011",16685 => "10000100",16686 => "00110010",16687 => "00000110",16688 => "01010101",16689 => "10001110",16690 => "01101111",16691 => "01110110",16692 => "11111010",16693 => "11000100",16694 => "11111100",16695 => "10001011",16696 => "11111011",16697 => "01000100",16698 => "10101101",16699 => "11010011",16700 => "10101110",16701 => "10101111",16702 => "00010000",16703 => "11100111",16704 => "11100101",16705 => "01101111",16706 => "00111001",16707 => "10110100",16708 => "11111000",16709 => "01110101",16710 => "10010101",16711 => "10010011",16712 => "11011001",16713 => "11110001",16714 => "10011110",16715 => "11011000",16716 => "11111111",16717 => "10001100",16718 => "01001111",16719 => "10001110",16720 => "10011010",16721 => "10011001",16722 => "00101100",16723 => "01101001",16724 => "11110001",16725 => "10000001",16726 => "01111101",16727 => "01000011",16728 => "10001110",16729 => "11110010",16730 => "11100101",16731 => "01110101",16732 => "01010101",16733 => "00100101",16734 => "00000001",16735 => "11100010",16736 => "10010001",16737 => "01111100",16738 => "00100001",16739 => "01110100",16740 => "11011100",16741 => "10100111",16742 => "11101100",16743 => "10100110",16744 => "01111001",16745 => "10011001",16746 => "11111101",16747 => "01111000",16748 => "01011010",16749 => "00000110",16750 => "01001100",16751 => "00000110",16752 => "11110001",16753 => "00101101",16754 => "10100010",16755 => "01110000",16756 => "01100101",16757 => "01011011",16758 => "01100001",16759 => "00001001",16760 => "11000101",16761 => "11110010",16762 => "10101100",16763 => "00000110",16764 => "01001101",16765 => "01111000",16766 => "11011101",16767 => "00010001",16768 => "10001101",16769 => "10111000",16770 => "00110111",16771 => "01110000",16772 => "11011001",16773 => "11101100",16774 => "11000010",16775 => "01001001",16776 => "01110001",16777 => "11110001",16778 => "10101110",16779 => "00100010",16780 => "01011101",16781 => "10101001",16782 => "01100011",16783 => "01011111",16784 => "01011001",16785 => "10001011",16786 => "01010011",16787 => "01110001",16788 => "11000001",16789 => "01100011",16790 => "01100110",16791 => "11111110",16792 => "00111010",16793 => "00110101",16794 => "00011110",16795 => "10111100",16796 => "11101110",16797 => "10100010",16798 => "00000101",16799 => "11010001",16800 => "00111100",16801 => "10100011",16802 => "10000000",16803 => "10000111",16804 => "11010001",16805 => "00101011",16806 => "00110000",16807 => "00101000",16808 => "10100010",16809 => "11100000",16810 => "00111110",16811 => "01011001",16812 => "00111110",16813 => "01100010",16814 => "01011101",16815 => "01111111",16816 => "01010000",16817 => "01110001",16818 => "11100000",16819 => "00110100",16820 => "11111001",16821 => "11010101",16822 => "01010011",16823 => "11010111",16824 => "11100001",16825 => "00000100",16826 => "11110101",16827 => "11001011",16828 => "10110101",16829 => "01001001",16830 => "00000110",16831 => "10000001",16832 => "00011101",16833 => "10000101",16834 => "10101001",16835 => "00101001",16836 => "00101110",16837 => "00110110",16838 => "11011000",16839 => "01100100",16840 => "10010011",16841 => "01111001",16842 => "10011111",16843 => "00110000",16844 => "01110010",16845 => "10110000",16846 => "00111010",16847 => "00110100",16848 => "01010000",16849 => "01001000",16850 => "00111100",16851 => "10001000",16852 => "11000011",16853 => "00110101",16854 => "00000110",16855 => "11001000",16856 => "01111011",16857 => "11000011",16858 => "00011100",16859 => "10110100",16860 => "11001001",16861 => "00000111",16862 => "01001001",16863 => "11011111",16864 => "11001110",16865 => "10001011",16866 => "11101110",16867 => "01011111",16868 => "10111111",16869 => "00010001",16870 => "10010001",16871 => "01100010",16872 => "01000111",16873 => "10011100",16874 => "00001011",16875 => "01101001",16876 => "10010100",16877 => "11000000",16878 => "00100011",16879 => "00010000",16880 => "00101110",16881 => "11011010",16882 => "11110010",16883 => "11001000",16884 => "01000100",16885 => "10011010",16886 => "11110111",16887 => "00001000",16888 => "10000000",16889 => "00000011",16890 => "00001111",16891 => "10000001",16892 => "01001011",16893 => "10001111",16894 => "10000001",16895 => "01101000",16896 => "11010010",16897 => "10001101",16898 => "01110110",16899 => "01110010",16900 => "01111100",16901 => "01100010",16902 => "00001100",16903 => "10011011",16904 => "00110000",16905 => "00010111",16906 => "01011111",16907 => "10100110",16908 => "01101100",16909 => "00110011",16910 => "00000110",16911 => "10111010",16912 => "11110000",16913 => "00001101",16914 => "01010100",16915 => "11110111",16916 => "10100011",16917 => "10100110",16918 => "11100110",16919 => "10111000",16920 => "01111100",16921 => "11110110",16922 => "10000100",16923 => "00110001",16924 => "11001010",16925 => "01110001",16926 => "10001010",16927 => "00001101",16928 => "01101100",16929 => "01010001",16930 => "01111001",16931 => "11000001",16932 => "00100100",16933 => "11110111",16934 => "10111011",16935 => "10101001",16936 => "00000000",16937 => "10000001",16938 => "00001110",16939 => "10101010",16940 => "10101110",16941 => "11101100",16942 => "00101010",16943 => "11100011",16944 => "01000000",16945 => "10010100",16946 => "11101011",16947 => "00110001",16948 => "00111111",16949 => "00011001",16950 => "10100011",16951 => "10010101",16952 => "10001010",16953 => "00000110",16954 => "10111010",16955 => "01000000",16956 => "00011110",16957 => "11011010",16958 => "01110111",16959 => "11000010",16960 => "11110111",16961 => "10011101",16962 => "01100110",16963 => "11010011",16964 => "00101011",16965 => "00011010",16966 => "10001001",16967 => "10111111",16968 => "01110101",16969 => "10011011",16970 => "11000111",16971 => "10100010",16972 => "00111010",16973 => "00000000",16974 => "11100111",16975 => "10100101",16976 => "01011110",16977 => "10011101",16978 => "00010000",16979 => "01101100",16980 => "01100010",16981 => "00000100",16982 => "11101101",16983 => "01110011",16984 => "10101110",16985 => "00010100",16986 => "11011111",16987 => "00100111",16988 => "11011000",16989 => "11011011",16990 => "10100100",16991 => "11000011",16992 => "10110100",16993 => "10111000",16994 => "10100010",16995 => "11001001",16996 => "01101110",16997 => "00111101",16998 => "10100101",16999 => "01000101",17000 => "00000011",17001 => "10110100",17002 => "10010000",17003 => "00001010",17004 => "11101100",17005 => "01111000",17006 => "10000100",17007 => "00011110",17008 => "01100010",17009 => "01000101",17010 => "01000011",17011 => "01111001",17012 => "10001000",17013 => "01000110",17014 => "00100111",17015 => "11011010",17016 => "11010100",17017 => "11101001",17018 => "11111100",17019 => "10001100",17020 => "11110100",17021 => "10110001",17022 => "00100101",17023 => "01010001",17024 => "10110011",17025 => "00111011",17026 => "10010110",17027 => "01100111",17028 => "00010110",17029 => "11100010",17030 => "11000101",17031 => "11010110",17032 => "10010100",17033 => "11010100",17034 => "01010011",17035 => "10001101",17036 => "01000101",17037 => "10101100",17038 => "11000101",17039 => "00100011",17040 => "01111100",17041 => "01110101",17042 => "11001100",17043 => "10100111",17044 => "00100000",17045 => "10010101",17046 => "00011001",17047 => "01100111",17048 => "01011010",17049 => "11010110",17050 => "00111100",17051 => "10111111",17052 => "11000100",17053 => "01111001",17054 => "00110111",17055 => "00000101",17056 => "10001100",17057 => "00111100",17058 => "10010110",17059 => "01110011",17060 => "11101101",17061 => "01011110",17062 => "10111010",17063 => "01111011",17064 => "11010010",17065 => "00010000",17066 => "00111010",17067 => "11101000",17068 => "01000011",17069 => "01011110",17070 => "00111100",17071 => "10000110",17072 => "10010010",17073 => "01101000",17074 => "10011111",17075 => "11000110",17076 => "11111100",17077 => "10100010",17078 => "01001100",17079 => "01100111",17080 => "00110011",17081 => "11000010",17082 => "10001000",17083 => "10100011",17084 => "10111000",17085 => "01111111",17086 => "00100000",17087 => "10010100",17088 => "01000010",17089 => "01001111",17090 => "00000110",17091 => "10111100",17092 => "10011011",17093 => "00001000",17094 => "00101001",17095 => "11110110",17096 => "00011111",17097 => "00110101",17098 => "10001011",17099 => "01100011",17100 => "01110010",17101 => "00110111",17102 => "10100001",17103 => "01011100",17104 => "10110101",17105 => "00010010",17106 => "11110111",17107 => "11011110",17108 => "00011110",17109 => "01011001",17110 => "11101100",17111 => "10010110",17112 => "01111100",17113 => "11100110",17114 => "10000001",17115 => "10111110",17116 => "10101001",17117 => "01110000",17118 => "01100000",17119 => "11011010",17120 => "01100010",17121 => "10110100",17122 => "01011111",17123 => "00000010",17124 => "01000011",17125 => "00011001",17126 => "11101110",17127 => "00100010",17128 => "01010011",17129 => "01011101",17130 => "10000110",17131 => "10000110",17132 => "11101100",17133 => "01101100",17134 => "11011110",17135 => "11101110",17136 => "01000111",17137 => "10100101",17138 => "00010100",17139 => "11011110",17140 => "10010110",17141 => "00001000",17142 => "01101111",17143 => "11010000",17144 => "01011110",17145 => "11111000",17146 => "01001110",17147 => "11100010",17148 => "00110111",17149 => "01001010",17150 => "11100101",17151 => "00010111",17152 => "00011111",17153 => "11100101",17154 => "01011011",17155 => "11101010",17156 => "10010111",17157 => "01110100",17158 => "11000010",17159 => "10100110",17160 => "01000110",17161 => "10000111",17162 => "10110010",17163 => "11010101",17164 => "11100011",17165 => "00010010",17166 => "00100011",17167 => "11100101",17168 => "01110101",17169 => "00000111",17170 => "00000011",17171 => "11010001",17172 => "11111001",17173 => "00110010",17174 => "11111001",17175 => "10011000",17176 => "01111110",17177 => "10101100",17178 => "00100010",17179 => "01100010",17180 => "10101001",17181 => "01011111",17182 => "11010110",17183 => "00011111",17184 => "01111010",17185 => "00000000",17186 => "11010010",17187 => "00000111",17188 => "11101110",17189 => "01100011",17190 => "01111111",17191 => "11111001",17192 => "01111111",17193 => "11011101",17194 => "01111101",17195 => "01101011",17196 => "10001110",17197 => "01011100",17198 => "11011100",17199 => "11111101",17200 => "00111101",17201 => "00011000",17202 => "00011010",17203 => "10110110",17204 => "01010101",17205 => "01110000",17206 => "01011000",17207 => "01010101",17208 => "01001001",17209 => "00101101",17210 => "01011001",17211 => "11010111",17212 => "01101000",17213 => "01100010",17214 => "01101110",17215 => "11011110",17216 => "01001100",17217 => "01100111",17218 => "00010000",17219 => "11101111",17220 => "01010001",17221 => "10110110",17222 => "01100000",17223 => "10110011",17224 => "01001010",17225 => "00100100",17226 => "11101011",17227 => "01010100",17228 => "10011111",17229 => "00101000",17230 => "01001110",17231 => "10001011",17232 => "10100000",17233 => "11000000",17234 => "10101011",17235 => "10111111",17236 => "10010110",17237 => "01110000",17238 => "10011000",17239 => "00101100",17240 => "11010111",17241 => "10011100",17242 => "10110101",17243 => "10011101",17244 => "01111110",17245 => "10101000",17246 => "10110010",17247 => "11011000",17248 => "10110111",17249 => "11001010",17250 => "10010010",17251 => "11011000",17252 => "10101100",17253 => "10110110",17254 => "11101000",17255 => "00111011",17256 => "01011000",17257 => "10010010",17258 => "00000001",17259 => "01011100",17260 => "11010010",17261 => "01100001",17262 => "01011111",17263 => "00110010",17264 => "00000110",17265 => "10011101",17266 => "11011111",17267 => "01011100",17268 => "10000000",17269 => "10101101",17270 => "00110001",17271 => "00110011",17272 => "11100011",17273 => "01111000",17274 => "11011110",17275 => "11110111",17276 => "00100000",17277 => "00101101",17278 => "10101111",17279 => "11011010",17280 => "10100111",17281 => "11110101",17282 => "01000101",17283 => "01110110",17284 => "10001000",17285 => "10100111",17286 => "00010010",17287 => "00000110",17288 => "01110111",17289 => "01010011",17290 => "11111101",17291 => "10011101",17292 => "01001101",17293 => "11110111",17294 => "11110101",17295 => "01010111",17296 => "10100111",17297 => "10110000",17298 => "11110111",17299 => "01000001",17300 => "01000001",17301 => "11100010",17302 => "10001101",17303 => "00000101",17304 => "10101100",17305 => "00000101",17306 => "01001110",17307 => "11010100",17308 => "01001000",17309 => "10101010",17310 => "11111111",17311 => "00100010",17312 => "01000110",17313 => "00000011",17314 => "10010100",17315 => "10100100",17316 => "11011001",17317 => "00111101",17318 => "01110110",17319 => "01010010",17320 => "00111010",17321 => "11101000",17322 => "11000100",17323 => "00100010",17324 => "01111111",17325 => "00110100",17326 => "01001000",17327 => "00000001",17328 => "10010100",17329 => "00001111",17330 => "00101010",17331 => "11010101",17332 => "10111100",17333 => "01010001",17334 => "11101011",17335 => "01000111",17336 => "11011101",17337 => "00011001",17338 => "00111001",17339 => "00000010",17340 => "01110111",17341 => "10101011",17342 => "10010100",17343 => "10000001",17344 => "10000100",17345 => "11110111",17346 => "00001010",17347 => "00000111",17348 => "11011001",17349 => "11000110",17350 => "11000101",17351 => "10010100",17352 => "01110001",17353 => "01010100",17354 => "11001110",17355 => "00001101",17356 => "00100001",17357 => "01011100",17358 => "00110010",17359 => "00001100",17360 => "01100000",17361 => "01101011",17362 => "01110100",17363 => "10110000",17364 => "10110011",17365 => "01110100",17366 => "01010110",17367 => "01111000",17368 => "00110101",17369 => "01110010",17370 => "11001011",17371 => "00011111",17372 => "11010101",17373 => "11000001",17374 => "10100110",17375 => "01110100",17376 => "00001110",17377 => "10100010",17378 => "10010001",17379 => "00011110",17380 => "00001110",17381 => "00001100",17382 => "11110000",17383 => "11100001",17384 => "10111000",17385 => "10100101",17386 => "00010101",17387 => "01001001",17388 => "00001100",17389 => "11101101",17390 => "00101100",17391 => "01001000",17392 => "01111010",17393 => "10101111",17394 => "00011101",17395 => "00101000",17396 => "01001110",17397 => "10001100",17398 => "00000111",17399 => "11101001",17400 => "01010010",17401 => "00111011",17402 => "11010111",17403 => "01111011",17404 => "00111001",17405 => "10001011",17406 => "11100001",17407 => "11010000",17408 => "00010010",17409 => "01101011",17410 => "01100100",17411 => "00110001",17412 => "11000000",17413 => "10000001",17414 => "00001101",17415 => "00100001",17416 => "00001000",17417 => "01010100",17418 => "11011000",17419 => "00111001",17420 => "00101101",17421 => "10011101",17422 => "10101110",17423 => "10001100",17424 => "10001110",17425 => "11100000",17426 => "10111001",17427 => "10110001",17428 => "10110001",17429 => "11010001",17430 => "11000111",17431 => "10000001",17432 => "11010001",17433 => "00100000",17434 => "01011010",17435 => "10111000",17436 => "11011001",17437 => "10010011",17438 => "00010010",17439 => "00000101",17440 => "00010011",17441 => "10000110",17442 => "10111010",17443 => "00101000",17444 => "01111010",17445 => "11100000",17446 => "10000110",17447 => "10101100",17448 => "11100111",17449 => "00011011",17450 => "10111101",17451 => "00001000",17452 => "10100110",17453 => "01110001",17454 => "10001111",17455 => "00110111",17456 => "11100110",17457 => "10101100",17458 => "01010000",17459 => "10110000",17460 => "01011101",17461 => "10001100",17462 => "11000001",17463 => "01011001",17464 => "10111001",17465 => "10101010",17466 => "00100001",17467 => "00011001",17468 => "00101111",17469 => "10111001",17470 => "01110010",17471 => "11000100",17472 => "01000010",17473 => "00101011",17474 => "00100110",17475 => "01100010",17476 => "10101001",17477 => "10011011",17478 => "11001010",17479 => "00011001",17480 => "01100011",17481 => "00010001",17482 => "10110100",17483 => "10110010",17484 => "01101001",17485 => "01111000",17486 => "10010110",17487 => "10101100",17488 => "00101100",17489 => "00000110",17490 => "11101100",17491 => "00011000",17492 => "00101110",17493 => "00100000",17494 => "11001100",17495 => "10010110",17496 => "00001110",17497 => "11010100",17498 => "10110001",17499 => "10101000",17500 => "10111011",17501 => "01100101",17502 => "01000101",17503 => "00100101",17504 => "11000001",17505 => "11010011",17506 => "11011101",17507 => "11001111",17508 => "10001111",17509 => "11000010",17510 => "11000100",17511 => "11001110",17512 => "10011011",17513 => "00001001",17514 => "11100100",17515 => "01100001",17516 => "10000111",17517 => "00001000",17518 => "11110111",17519 => "01001110",17520 => "01110000",17521 => "00110000",17522 => "11000000",17523 => "10101011",17524 => "00000110",17525 => "11100010",17526 => "01110101",17527 => "01111011",17528 => "10110100",17529 => "11101100",17530 => "10011110",17531 => "10100011",17532 => "10110111",17533 => "11001001",17534 => "01100110",17535 => "00000100",17536 => "00111010",17537 => "10001110",17538 => "00011010",17539 => "00001011",17540 => "10010111",17541 => "01101100",17542 => "00100001",17543 => "00011000",17544 => "10110100",17545 => "01111011",17546 => "11110100",17547 => "01100001",17548 => "01001101",17549 => "11000010",17550 => "01011010",17551 => "11010110",17552 => "01000001",17553 => "01010001",17554 => "11001101",17555 => "00100000",17556 => "01000001",17557 => "11001110",17558 => "00101010",17559 => "10100100",17560 => "00001100",17561 => "01100101",17562 => "11110000",17563 => "01110010",17564 => "11000101",17565 => "11010001",17566 => "00100100",17567 => "01010001",17568 => "00010110",17569 => "00100010",17570 => "00100111",17571 => "01001101",17572 => "01110111",17573 => "01001011",17574 => "01001111",17575 => "00110100",17576 => "01111001",17577 => "11110100",17578 => "01101101",17579 => "01011010",17580 => "10110110",17581 => "11100011",17582 => "01010010",17583 => "01101001",17584 => "00010111",17585 => "10110110",17586 => "11001101",17587 => "01010100",17588 => "10011010",17589 => "00000111",17590 => "01101111",17591 => "11101100",17592 => "10001101",17593 => "01100001",17594 => "01101101",17595 => "01111010",17596 => "10111111",17597 => "01111000",17598 => "00011111",17599 => "01101011",17600 => "00111100",17601 => "01100001",17602 => "00100111",17603 => "00001010",17604 => "01111001",17605 => "11111010",17606 => "10010000",17607 => "01010100",17608 => "00111010",17609 => "01010000",17610 => "11011010",17611 => "10011101",17612 => "01110010",17613 => "01110111",17614 => "00100001",17615 => "10101000",17616 => "01000000",17617 => "10100111",17618 => "11101101",17619 => "01000001",17620 => "11011011",17621 => "11101100",17622 => "00100100",17623 => "11001011",17624 => "11011011",17625 => "11101001",17626 => "11011010",17627 => "11000101",17628 => "10111010",17629 => "11001110",17630 => "10011111",17631 => "11111111",17632 => "11010111",17633 => "00111100",17634 => "10011001",17635 => "01111110",17636 => "00111001",17637 => "11010101",17638 => "00010000",17639 => "10111010",17640 => "10001111",17641 => "00111000",17642 => "10000010",17643 => "01100111",17644 => "10000000",17645 => "00110011",17646 => "11010010",17647 => "10011010",17648 => "11110000",17649 => "11001100",17650 => "01011010",17651 => "00101011",17652 => "01111101",17653 => "00100000",17654 => "01101000",17655 => "01001011",17656 => "01110010",17657 => "11101010",17658 => "11101111",17659 => "10011101",17660 => "00011000",17661 => "00111101",17662 => "11100011",17663 => "00110001",17664 => "00010101",17665 => "01110100",17666 => "10010010",17667 => "10100011",17668 => "00011000",17669 => "11111111",17670 => "10011001",17671 => "10110100",17672 => "01000001",17673 => "11111111",17674 => "10111000",17675 => "11010110",17676 => "11001111",17677 => "10011100",17678 => "11000001",17679 => "10011111",17680 => "11000101",17681 => "10000111",17682 => "00100111",17683 => "01111010",17684 => "00110011",17685 => "01011110",17686 => "01110000",17687 => "01000010",17688 => "00001101",17689 => "10100001",17690 => "01000010",17691 => "01100111",17692 => "00110001",17693 => "11010001",17694 => "00110000",17695 => "11100011",17696 => "10001101",17697 => "00111000",17698 => "10010100",17699 => "10100111",17700 => "10101111",17701 => "00111000",17702 => "10101101",17703 => "11111101",17704 => "01001000",17705 => "01101101",17706 => "11111100",17707 => "11101110",17708 => "00000001",17709 => "01010001",17710 => "10001111",17711 => "00100001",17712 => "01101111",17713 => "00011011",17714 => "10101101",17715 => "01101111",17716 => "10111100",17717 => "11111101",17718 => "10100010",17719 => "01000111",17720 => "10111100",17721 => "00001000",17722 => "01010111",17723 => "00011110",17724 => "00000010",17725 => "11011001",17726 => "00110111",17727 => "11011011",17728 => "00111010",17729 => "10010000",17730 => "10110000",17731 => "10000100",17732 => "00100010",17733 => "01000110",17734 => "11000100",17735 => "10100001",17736 => "00101110",17737 => "01111100",17738 => "01010100",17739 => "11110101",17740 => "10001010",17741 => "00110100",17742 => "10101000",17743 => "10001110",17744 => "10010001",17745 => "00110101",17746 => "11111010",17747 => "01000001",17748 => "01110010",17749 => "10111000",17750 => "11101011",17751 => "11001000",17752 => "10110111",17753 => "11110000",17754 => "00111001",17755 => "01110100",17756 => "01001111",17757 => "01001010",17758 => "00001101",17759 => "10010101",17760 => "10010101",17761 => "01000001",17762 => "00010011",17763 => "11111011",17764 => "00000100",17765 => "01101100",17766 => "11100111",17767 => "10010100",17768 => "00001010",17769 => "00010101",17770 => "11010111",17771 => "10101111",17772 => "01011011",17773 => "01100111",17774 => "01000001",17775 => "01100110",17776 => "10000000",17777 => "01001001",17778 => "11001010",17779 => "11010101",17780 => "11001000",17781 => "10111000",17782 => "01110101",17783 => "10011110",17784 => "11000110",17785 => "01000111",17786 => "11100001",17787 => "11110001",17788 => "00111110",17789 => "01011011",17790 => "11010001",17791 => "01010010",17792 => "00101110",17793 => "10101011",17794 => "10100000",17795 => "01011000",17796 => "00001000",17797 => "11001010",17798 => "10000000",17799 => "11100110",17800 => "10100101",17801 => "00111101",17802 => "00001000",17803 => "10111010",17804 => "00011101",17805 => "11010111",17806 => "10111110",17807 => "11101001",17808 => "00001010",17809 => "01001010",17810 => "01110011",17811 => "10001001",17812 => "01011000",17813 => "00110001",17814 => "11101000",17815 => "10000001",17816 => "11010000",17817 => "11100110",17818 => "01111100",17819 => "01001111",17820 => "00110100",17821 => "11110011",17822 => "01101101",17823 => "11001100",17824 => "11100011",17825 => "10010111",17826 => "00101001",17827 => "01010101",17828 => "01110111",17829 => "10001011",17830 => "01101011",17831 => "00001000",17832 => "11111011",17833 => "00000011",17834 => "00111110",17835 => "10001100",17836 => "01010010",17837 => "00010101",17838 => "00111100",17839 => "11100011",17840 => "01101110",17841 => "00101110",17842 => "01000111",17843 => "10000101",17844 => "00000010",17845 => "01110111",17846 => "00000001",17847 => "11100100",17848 => "01101001",17849 => "01000111",17850 => "00000111",17851 => "11101011",17852 => "00001110",17853 => "01010100",17854 => "10010101",17855 => "01111110",17856 => "11111001",17857 => "11101010",17858 => "00000111",17859 => "00000111",17860 => "00001111",17861 => "01111100",17862 => "01011001",17863 => "01110111",17864 => "01100000",17865 => "10100100",17866 => "10101011",17867 => "01010101",17868 => "11111000",17869 => "11010110",17870 => "01001110",17871 => "11101111",17872 => "11011001",17873 => "01001001",17874 => "10110111",17875 => "11101011",17876 => "11001100",17877 => "00100000",17878 => "01101100",17879 => "01010010",17880 => "10100011",17881 => "01001101",17882 => "00110011",17883 => "00011111",17884 => "10001000",17885 => "01101000",17886 => "10011011",17887 => "00010111",17888 => "10101010",17889 => "10111110",17890 => "00101110",17891 => "10000100",17892 => "01011111",17893 => "00001011",17894 => "00000101",17895 => "01011100",17896 => "11101100",17897 => "11111111",17898 => "10001100",17899 => "01000000",17900 => "01111100",17901 => "00111011",17902 => "11001000",17903 => "00001110",17904 => "00110000",17905 => "00010001",17906 => "00101000",17907 => "00000001",17908 => "10011010",17909 => "00101010",17910 => "11101000",17911 => "10000000",17912 => "01011110",17913 => "11110000",17914 => "01010001",17915 => "10011001",17916 => "11010100",17917 => "10011001",17918 => "01100011",17919 => "11010000",17920 => "01011011",17921 => "00010100",17922 => "01110100",17923 => "11010000",17924 => "00001001",17925 => "00000111",17926 => "01010100",17927 => "00110000",17928 => "00010100",17929 => "10111100",17930 => "00001110",17931 => "01110100",17932 => "00111110",17933 => "10000111",17934 => "11110100",17935 => "00100101",17936 => "10100001",17937 => "00001001",17938 => "10100000",17939 => "11111010",17940 => "00000110",17941 => "11001001",17942 => "01100110",17943 => "00111010",17944 => "11101110",17945 => "00001001",17946 => "01010101",17947 => "11100011",17948 => "10001000",17949 => "11001100",17950 => "11111001",17951 => "11101010",17952 => "10000110",17953 => "11110101",17954 => "10000101",17955 => "00001000",17956 => "01010011",17957 => "01111001",17958 => "11000100",17959 => "00001101",17960 => "00101000",17961 => "00111101",17962 => "00100000",17963 => "00111100",17964 => "10101110",17965 => "10011011",17966 => "00010110",17967 => "00010110",17968 => "11111111",17969 => "10100110",17970 => "00010100",17971 => "11111001",17972 => "00011011",17973 => "10010101",17974 => "01100001",17975 => "00010101",17976 => "11001000",17977 => "10110010",17978 => "11011010",17979 => "11100001",17980 => "01110111",17981 => "01000010",17982 => "11100110",17983 => "00010001",17984 => "00101110",17985 => "01110101",17986 => "10100010",17987 => "01000110",17988 => "00001010",17989 => "01001110",17990 => "11100011",17991 => "01010111",17992 => "11011000",17993 => "11111000",17994 => "00111111",17995 => "00011100",17996 => "10010001",17997 => "01000000",17998 => "11111000",17999 => "01101100",18000 => "01111111",18001 => "00111000",18002 => "00010100",18003 => "11101101",18004 => "00011011",18005 => "01010101",18006 => "11000111",18007 => "01000101",18008 => "11111010",18009 => "01000110",18010 => "10111000",18011 => "00010001",18012 => "00110011",18013 => "10010010",18014 => "00010101",18015 => "00011111",18016 => "00000010",18017 => "10010000",18018 => "11111001",18019 => "11010001",18020 => "11001100",18021 => "11010001",18022 => "11000100",18023 => "11001001",18024 => "01110010",18025 => "10101111",18026 => "00010111",18027 => "11111011",18028 => "01011111",18029 => "00000001",18030 => "00011110",18031 => "10101000",18032 => "01000100",18033 => "10101110",18034 => "10110000",18035 => "10100011",18036 => "10010011",18037 => "00101011",18038 => "11011000",18039 => "01011001",18040 => "10110111",18041 => "10000000",18042 => "00110000",18043 => "00010011",18044 => "11010011",18045 => "01110101",18046 => "01011110",18047 => "01011000",18048 => "10001111",18049 => "11011100",18050 => "11011111",18051 => "00110101",18052 => "10100010",18053 => "01000000",18054 => "01010110",18055 => "11100111",18056 => "01100101",18057 => "00110111",18058 => "00101011",18059 => "00011000",18060 => "00000011",18061 => "10000000",18062 => "00101101",18063 => "10011011",18064 => "00000101",18065 => "00100111",18066 => "01000011",18067 => "01011001",18068 => "10000110",18069 => "00011010",18070 => "10011000",18071 => "00000111",18072 => "01010011",18073 => "01001110",18074 => "11001000",18075 => "11111101",18076 => "00000011",18077 => "01111000",18078 => "10111011",18079 => "01100111",18080 => "11111010",18081 => "01100000",18082 => "11011110",18083 => "01011010",18084 => "00001010",18085 => "00011110",18086 => "10101100",18087 => "10110011",18088 => "11111001",18089 => "01101000",18090 => "11011000",18091 => "11001011",18092 => "11000101",18093 => "00010110",18094 => "01110001",18095 => "11110000",18096 => "01000110",18097 => "01001000",18098 => "00010101",18099 => "11100111",18100 => "00000010",18101 => "01111100",18102 => "00111111",18103 => "01001000",18104 => "01111001",18105 => "00111000",18106 => "11001110",18107 => "00100001",18108 => "00101111",18109 => "10110011",18110 => "10110010",18111 => "00111101",18112 => "11010111",18113 => "10110010",18114 => "10000101",18115 => "10001100",18116 => "01000011",18117 => "00100100",18118 => "01101111",18119 => "11011000",18120 => "11101101",18121 => "01110111",18122 => "10010001",18123 => "11100000",18124 => "10011100",18125 => "01110000",18126 => "01000001",18127 => "11110110",18128 => "01100101",18129 => "01011010",18130 => "01100001",18131 => "01001010",18132 => "01010101",18133 => "11001011",18134 => "00101011",18135 => "00011000",18136 => "00110100",18137 => "01101010",18138 => "00111011",18139 => "00001001",18140 => "00101110",18141 => "00011110",18142 => "01100001",18143 => "11100000",18144 => "01000001",18145 => "10001001",18146 => "10110110",18147 => "01010000",18148 => "11100100",18149 => "11101110",18150 => "00100110",18151 => "01011110",18152 => "00010100",18153 => "11111011",18154 => "01111101",18155 => "10001100",18156 => "01110111",18157 => "11001001",18158 => "11110001",18159 => "00011100",18160 => "00110110",18161 => "11101011",18162 => "01010111",18163 => "01010110",18164 => "00101001",18165 => "01110000",18166 => "11010110",18167 => "10101011",18168 => "10000111",18169 => "11000110",18170 => "01111101",18171 => "10001001",18172 => "10100110",18173 => "01110010",18174 => "01000100",18175 => "11010110",18176 => "01011100",18177 => "11001101",18178 => "00111111",18179 => "00111111",18180 => "01111011",18181 => "00000011",18182 => "11111000",18183 => "01100000",18184 => "01100000",18185 => "01100101",18186 => "11000100",18187 => "01110010",18188 => "01101010",18189 => "11010100",18190 => "10001011",18191 => "11011011",18192 => "10100000",18193 => "10101111",18194 => "10010000",18195 => "01010101",18196 => "01010101",18197 => "11001010",18198 => "10000010",18199 => "00110101",18200 => "11001101",18201 => "01111101",18202 => "00110001",18203 => "00001111",18204 => "01011011",18205 => "00101111",18206 => "01101100",18207 => "00010000",18208 => "11011111",18209 => "00110111",18210 => "11100010",18211 => "01010111",18212 => "11111011",18213 => "11110111",18214 => "10101110",18215 => "01001001",18216 => "10010011",18217 => "00101110",18218 => "10100010",18219 => "10000010",18220 => "00011100",18221 => "10100010",18222 => "00001110",18223 => "01110100",18224 => "01000101",18225 => "00001111",18226 => "11110010",18227 => "11000100",18228 => "01010100",18229 => "10010011",18230 => "10010111",18231 => "10001010",18232 => "11101111",18233 => "10111100",18234 => "11010110",18235 => "11000011",18236 => "00100011",18237 => "00000101",18238 => "01111100",18239 => "11100000",18240 => "01110011",18241 => "01011001",18242 => "11010101",18243 => "00111111",18244 => "00110100",18245 => "10110010",18246 => "00100101",18247 => "10110100",18248 => "01100111",18249 => "00100101",18250 => "00111000",18251 => "10110000",18252 => "10001110",18253 => "00010101",18254 => "11100101",18255 => "00000000",18256 => "00101111",18257 => "11000011",18258 => "00101101",18259 => "01010101",18260 => "11001111",18261 => "10101110",18262 => "00001010",18263 => "01110111",18264 => "00000010",18265 => "00011100",18266 => "11001100",18267 => "00111101",18268 => "00001111",18269 => "11000111",18270 => "11000000",18271 => "00100101",18272 => "10111111",18273 => "01011011",18274 => "00111000",18275 => "00000101",18276 => "00111101",18277 => "00001101",18278 => "11010110",18279 => "10011010",18280 => "11000100",18281 => "00111011",18282 => "10010101",18283 => "11110110",18284 => "00011010",18285 => "10100110",18286 => "11110110",18287 => "10101010",18288 => "10110111",18289 => "00110010",18290 => "11010100",18291 => "10100101",18292 => "01010101",18293 => "11111110",18294 => "10001000",18295 => "10010000",18296 => "01111001",18297 => "01011111",18298 => "11100001",18299 => "10110011",18300 => "00101011",18301 => "00001101",18302 => "01101011",18303 => "00010111",18304 => "10111011",18305 => "00110100",18306 => "10100001",18307 => "10010001",18308 => "00010100",18309 => "01101111",18310 => "00010011",18311 => "10000001",18312 => "01001011",18313 => "10101010",18314 => "00001011",18315 => "11000111",18316 => "10001001",18317 => "00011001",18318 => "10111011",18319 => "11110101",18320 => "00110011",18321 => "00110000",18322 => "11110110",18323 => "01000100",18324 => "10000000",18325 => "00001111",18326 => "11001111",18327 => "10010100",18328 => "01001100",18329 => "11100011",18330 => "10000000",18331 => "01101111",18332 => "01000001",18333 => "10011011",18334 => "10001110",18335 => "01110010",18336 => "00101111",18337 => "00010001",18338 => "01100011",18339 => "00011100",18340 => "00111111",18341 => "01111101",18342 => "10010000",18343 => "00110111",18344 => "11111100",18345 => "00010100",18346 => "11111101",18347 => "00110110",18348 => "00101001",18349 => "11110110",18350 => "01111100",18351 => "10010001",18352 => "10000111",18353 => "01010000",18354 => "01100011",18355 => "01011011",18356 => "11011101",18357 => "01100010",18358 => "00100110",18359 => "11100011",18360 => "11011100",18361 => "11111000",18362 => "10000100",18363 => "01011010",18364 => "01010000",18365 => "01000110",18366 => "01001101",18367 => "00101000",18368 => "00100000",18369 => "01001001",18370 => "10010101",18371 => "10110010",18372 => "01000001",18373 => "10001101",18374 => "01011001",18375 => "01111010",18376 => "10100001",18377 => "10101000",18378 => "00100011",18379 => "10110101",18380 => "00110001",18381 => "01101001",18382 => "01011101",18383 => "10000011",18384 => "11001010",18385 => "10011000",18386 => "00100111",18387 => "01100000",18388 => "10101001",18389 => "11110100",18390 => "01101110",18391 => "01101011",18392 => "11110011",18393 => "11011111",18394 => "10000100",18395 => "00011000",18396 => "11100110",18397 => "10000010",18398 => "10010101",18399 => "01110011",18400 => "11111110",18401 => "10010101",18402 => "10111001",18403 => "01111110",18404 => "11101110",18405 => "01100011",18406 => "00001010",18407 => "00110111",18408 => "11000011",18409 => "10101111",18410 => "01000000",18411 => "11000111",18412 => "11101010",18413 => "00101000",18414 => "00011000",18415 => "00101000",18416 => "10011110",18417 => "00000111",18418 => "10100100",18419 => "10001011",18420 => "11111110",18421 => "10111100",18422 => "00011010",18423 => "00000010",18424 => "01101101",18425 => "10110101",18426 => "10001001",18427 => "11110111",18428 => "10001111",18429 => "11100111",18430 => "11101100",18431 => "10110011",18432 => "01101011",18433 => "01011000",18434 => "10000010",18435 => "11100100",18436 => "11101001",18437 => "10100000",18438 => "11110011",18439 => "01111101",18440 => "00010111",18441 => "00000100",18442 => "11010101",18443 => "11010111",18444 => "10000111",18445 => "00011011",18446 => "00000011",18447 => "10101000",18448 => "00110001",18449 => "11101110",18450 => "11000010",18451 => "11110011",18452 => "01010110",18453 => "00110110",18454 => "01100111",18455 => "01101101",18456 => "01011100",18457 => "10111101",18458 => "00111001",18459 => "10101100",18460 => "11010110",18461 => "00110110",18462 => "11100100",18463 => "10110011",18464 => "00100010",18465 => "00010001",18466 => "10001000",18467 => "00011011",18468 => "00100110",18469 => "11111000",18470 => "11001100",18471 => "11111001",18472 => "11010110",18473 => "00111000",18474 => "10011000",18475 => "10111101",18476 => "10100011",18477 => "00110000",18478 => "01000011",18479 => "00101011",18480 => "00011001",18481 => "00101011",18482 => "11110001",18483 => "01110001",18484 => "11100100",18485 => "10111100",18486 => "10011101",18487 => "10111000",18488 => "01100000",18489 => "11100111",18490 => "10000110",18491 => "11001100",18492 => "10010011",18493 => "10000001",18494 => "01101011",18495 => "01111000",18496 => "10001100",18497 => "11001111",18498 => "01001110",18499 => "01110001",18500 => "10110100",18501 => "00111010",18502 => "01000100",18503 => "11001111",18504 => "10000001",18505 => "10000101",18506 => "00110110",18507 => "11110110",18508 => "11011010",18509 => "11100000",18510 => "01101110",18511 => "11001001",18512 => "00100011",18513 => "00000100",18514 => "10000010",18515 => "11110010",18516 => "01010111",18517 => "00111001",18518 => "11101101",18519 => "10011100",18520 => "10111111",18521 => "10001111",18522 => "01110011",18523 => "11001001",18524 => "01011101",18525 => "10000010",18526 => "01010101",18527 => "11010111",18528 => "01011101",18529 => "11100100",18530 => "01100110",18531 => "10101010",18532 => "00100011",18533 => "10111111",18534 => "10101111",18535 => "11000010",18536 => "10100100",18537 => "00110101",18538 => "10100011",18539 => "11101000",18540 => "00011101",18541 => "10010101",18542 => "11101000",18543 => "11000000",18544 => "10010011",18545 => "10100011",18546 => "01000111",18547 => "10011100",18548 => "00000001",18549 => "00000111",18550 => "00111100",18551 => "01110111",18552 => "01101000",18553 => "11010111",18554 => "01111000",18555 => "11101111",18556 => "10111101",18557 => "01101010",18558 => "00101001",18559 => "10000100",18560 => "00001010",18561 => "00010111",18562 => "11110110",18563 => "11011100",18564 => "00001101",18565 => "11010110",18566 => "00000101",18567 => "00010110",18568 => "00010111",18569 => "01011000",18570 => "11100011",18571 => "10101100",18572 => "00010001",18573 => "10101000",18574 => "01111101",18575 => "01100011",18576 => "01010000",18577 => "00110011",18578 => "10100101",18579 => "00101001",18580 => "01110101",18581 => "11011010",18582 => "11001110",18583 => "01100100",18584 => "01010000",18585 => "00000101",18586 => "01010011",18587 => "11011101",18588 => "10100000",18589 => "00110100",18590 => "01000000",18591 => "00100001",18592 => "01100010",18593 => "10111000",18594 => "11100111",18595 => "11111000",18596 => "01111111",18597 => "11001000",18598 => "10101111",18599 => "11001100",18600 => "00010010",18601 => "10110010",18602 => "11001001",18603 => "00110001",18604 => "11001001",18605 => "11101001",18606 => "11001101",18607 => "01000000",18608 => "00000101",18609 => "01111010",18610 => "11001100",18611 => "10111110",18612 => "11100001",18613 => "00010110",18614 => "11000111",18615 => "00110001",18616 => "11000000",18617 => "11000111",18618 => "10101111",18619 => "00010011",18620 => "11100010",18621 => "01010111",18622 => "00101111",18623 => "00010101",18624 => "10010010",18625 => "11111011",18626 => "10111111",18627 => "00001101",18628 => "01001000",18629 => "00010011",18630 => "01011110",18631 => "01001110",18632 => "10100000",18633 => "00010101",18634 => "00111110",18635 => "00101001",18636 => "00110111",18637 => "01010001",18638 => "00011111",18639 => "00110110",18640 => "10110001",18641 => "10000001",18642 => "10111101",18643 => "10001100",18644 => "10010101",18645 => "11110010",18646 => "11110111",18647 => "10110101",18648 => "10111001",18649 => "10001100",18650 => "00110001",18651 => "01011111",18652 => "10000001",18653 => "10010001",18654 => "01000000",18655 => "10101000",18656 => "11100010",18657 => "10111011",18658 => "01110100",18659 => "00101010",18660 => "00001011",18661 => "00011000",18662 => "00001100",18663 => "01101100",18664 => "01001111",18665 => "01000001",18666 => "10101010",18667 => "10001111",18668 => "10000100",18669 => "10100000",18670 => "01111011",18671 => "00011010",18672 => "11110110",18673 => "10100001",18674 => "11000101",18675 => "01010100",18676 => "10000101",18677 => "01000101",18678 => "01010110",18679 => "10101100",18680 => "01001110",18681 => "11100011",18682 => "10001011",18683 => "10001001",18684 => "10010001",18685 => "00111000",18686 => "00010001",18687 => "10110000",18688 => "01010010",18689 => "00111010",18690 => "00110100",18691 => "11101000",18692 => "11100010",18693 => "00001011",18694 => "11000011",18695 => "01111000",18696 => "10101100",18697 => "00100011",18698 => "00010010",18699 => "10100011",18700 => "00100000",18701 => "00110100",18702 => "10011001",18703 => "11000000",18704 => "11010011",18705 => "01110100",18706 => "01110110",18707 => "01000000",18708 => "10101010",18709 => "01000011",18710 => "00000000",18711 => "10100101",18712 => "00101101",18713 => "01001110",18714 => "11000001",18715 => "01111011",18716 => "10001100",18717 => "01011011",18718 => "10110100",18719 => "01111010",18720 => "01010100",18721 => "01100011",18722 => "11110010",18723 => "10100000",18724 => "10010101",18725 => "01101011",18726 => "10111101",18727 => "10101110",18728 => "11110100",18729 => "01010000",18730 => "01101001",18731 => "11011100",18732 => "01101100",18733 => "11101011",18734 => "11100101",18735 => "00011011",18736 => "11101010",18737 => "11000001",18738 => "01011110",18739 => "11100101",18740 => "01001000",18741 => "01011101",18742 => "01011010",18743 => "11000101",18744 => "00100110",18745 => "01011010",18746 => "01110101",18747 => "11101110",18748 => "10110011",18749 => "10010101",18750 => "00110111",18751 => "10000110",18752 => "00000101",18753 => "00111001",18754 => "00111110",18755 => "11001010",18756 => "11000000",18757 => "00000001",18758 => "10001111",18759 => "01101010",18760 => "10101111",18761 => "10011001",18762 => "00011100",18763 => "01000010",18764 => "01111011",18765 => "11011101",18766 => "01010110",18767 => "01001101",18768 => "01100001",18769 => "00001000",18770 => "00101110",18771 => "11101111",18772 => "01011001",18773 => "11000110",18774 => "10011000",18775 => "11011100",18776 => "10110101",18777 => "11100011",18778 => "10011111",18779 => "00001011",18780 => "00111100",18781 => "00100100",18782 => "11010011",18783 => "11000101",18784 => "01001011",18785 => "11100001",18786 => "00001000",18787 => "01000100",18788 => "10000010",18789 => "01010000",18790 => "01111001",18791 => "11110110",18792 => "00001001",18793 => "10011110",18794 => "10000110",18795 => "00011101",18796 => "10100011",18797 => "10011011",18798 => "11101001",18799 => "10110110",18800 => "00111100",18801 => "11011001",18802 => "00100101",18803 => "01110001",18804 => "10010111",18805 => "00001001",18806 => "10110110",18807 => "10010001",18808 => "11110001",18809 => "11111000",18810 => "11111110",18811 => "00100110",18812 => "01100110",18813 => "10110111",18814 => "00111010",18815 => "00110011",18816 => "11100011",18817 => "00001101",18818 => "10101001",18819 => "10000000",18820 => "00110000",18821 => "10110001",18822 => "00110010",18823 => "01111000",18824 => "10001101",18825 => "01011000",18826 => "00011010",18827 => "01101001",18828 => "01101001",18829 => "11111100",18830 => "11100000",18831 => "11000110",18832 => "11110001",18833 => "01001010",18834 => "10010000",18835 => "10001101",18836 => "10011101",18837 => "10011111",18838 => "01100000",18839 => "00011101",18840 => "01100010",18841 => "01001001",18842 => "11111000",18843 => "00110111",18844 => "10111101",18845 => "10001011",18846 => "10000111",18847 => "01011010",18848 => "10001000",18849 => "10100111",18850 => "00111111",18851 => "00110001",18852 => "10110111",18853 => "10010101",18854 => "11010001",18855 => "10000101",18856 => "01011110",18857 => "11101100",18858 => "11001011",18859 => "10010110",18860 => "01100011",18861 => "00000100",18862 => "01010011",18863 => "00101111",18864 => "11000000",18865 => "00111010",18866 => "01000100",18867 => "11001110",18868 => "00010100",18869 => "00100000",18870 => "10111011",18871 => "00000011",18872 => "00110001",18873 => "11011011",18874 => "10110011",18875 => "00111010",18876 => "00010100",18877 => "00000011",18878 => "11110010",18879 => "10000011",18880 => "01101111",18881 => "11111100",18882 => "00001111",18883 => "00101001",18884 => "01101111",18885 => "01000010",18886 => "11000001",18887 => "01101100",18888 => "11101000",18889 => "10110001",18890 => "11110101",18891 => "01001101",18892 => "01111110",18893 => "10111001",18894 => "00111000",18895 => "10011001",18896 => "10100100",18897 => "00110010",18898 => "00101011",18899 => "01101111",18900 => "01001110",18901 => "11000100",18902 => "11100001",18903 => "01011001",18904 => "01101010",18905 => "01110100",18906 => "01101100",18907 => "11111111",18908 => "00100110",18909 => "11010011",18910 => "01000110",18911 => "00000101",18912 => "11000101",18913 => "00110011",18914 => "11101100",18915 => "10100111",18916 => "01111001",18917 => "11001010",18918 => "10000101",18919 => "10000111",18920 => "00000100",18921 => "10100110",18922 => "01011010",18923 => "01101111",18924 => "01000011",18925 => "11100010",18926 => "01111000",18927 => "00010110",18928 => "00111000",18929 => "01011010",18930 => "00010000",18931 => "11100111",18932 => "11010001",18933 => "01011110",18934 => "10110100",18935 => "01001101",18936 => "10110110",18937 => "01101110",18938 => "10100010",18939 => "11001000",18940 => "10111001",18941 => "01011110",18942 => "11000011",18943 => "11100101",18944 => "11000110",18945 => "11111111",18946 => "11110101",18947 => "10101000",18948 => "00111100",18949 => "01000111",18950 => "10110100",18951 => "00111111",18952 => "10001101",18953 => "10010000",18954 => "10011110",18955 => "01000101",18956 => "00110001",18957 => "00100011",18958 => "01010000",18959 => "01100000",18960 => "10110000",18961 => "10111100",18962 => "10011010",18963 => "10010000",18964 => "01011110",18965 => "00110001",18966 => "11010101",18967 => "01111011",18968 => "10111111",18969 => "11001110",18970 => "01111011",18971 => "10111010",18972 => "10101011",18973 => "11001111",18974 => "01111010",18975 => "11011110",18976 => "10001011",18977 => "01100111",18978 => "01010010",18979 => "01011011",18980 => "10111010",18981 => "01101011",18982 => "00011110",18983 => "11001011",18984 => "10011010",18985 => "01000110",18986 => "00010010",18987 => "11100111",18988 => "10101111",18989 => "11001101",18990 => "11100110",18991 => "00100110",18992 => "11110111",18993 => "00111100",18994 => "10011110",18995 => "11111011",18996 => "00101100",18997 => "01110110",18998 => "11001010",18999 => "01011010",19000 => "11110100",19001 => "01010011",19002 => "01111110",19003 => "11110000",19004 => "10000000",19005 => "10100001",19006 => "00100100",19007 => "11111001",19008 => "01100111",19009 => "10011010",19010 => "10111001",19011 => "00111101",19012 => "10101000",19013 => "10110001",19014 => "00101011",19015 => "01010010",19016 => "00101011",19017 => "11100000",19018 => "01000010",19019 => "00010010",19020 => "00000010",19021 => "01011101",19022 => "10001110",19023 => "11110001",19024 => "00010010",19025 => "10101001",19026 => "11100011",19027 => "00011000",19028 => "01010100",19029 => "11001111",19030 => "10101100",19031 => "00101110",19032 => "10001011",19033 => "11101101",19034 => "11111000",19035 => "01000000",19036 => "01010001",19037 => "10000001",19038 => "11010110",19039 => "01000001",19040 => "00001001",19041 => "10111011",19042 => "11001101",19043 => "01100100",19044 => "00011000",19045 => "10000111",19046 => "10001000",19047 => "11011001",19048 => "00010110",19049 => "00111100",19050 => "10001000",19051 => "10111001",19052 => "00010000",19053 => "11111011",19054 => "01011000",19055 => "11010100",19056 => "10000100",19057 => "10110011",19058 => "01100110",19059 => "00111000",19060 => "10100101",19061 => "11010000",19062 => "01000010",19063 => "01011011",19064 => "01111010",19065 => "11000000",19066 => "10011001",19067 => "01101110",19068 => "00101000",19069 => "00000100",19070 => "01000011",19071 => "01110000",19072 => "10111111",19073 => "11001101",19074 => "01011010",19075 => "01000110",19076 => "11110010",19077 => "10010110",19078 => "10101100",19079 => "10110001",19080 => "10110100",19081 => "11001111",19082 => "10110100",19083 => "01110100",19084 => "00111101",19085 => "11011011",19086 => "00100000",19087 => "01001011",19088 => "00110000",19089 => "11001111",19090 => "10100110",19091 => "00111111",19092 => "11011000",19093 => "10111110",19094 => "10100110",19095 => "10111001",19096 => "11101001",19097 => "11000001",19098 => "11101011",19099 => "01010000",19100 => "00001010",19101 => "00011110",19102 => "00110000",19103 => "10001110",19104 => "01100011",19105 => "11000010",19106 => "01001101",19107 => "00100000",19108 => "01101001",19109 => "00011011",19110 => "00111110",19111 => "11101010",19112 => "01011100",19113 => "00111101",19114 => "11100000",19115 => "11111000",19116 => "10110110",19117 => "01010101",19118 => "00101110",19119 => "11110101",19120 => "00101010",19121 => "11111111",19122 => "10111010",19123 => "00011010",19124 => "11001010",19125 => "01000011",19126 => "10000001",19127 => "00010111",19128 => "10001101",19129 => "00011011",19130 => "00111111",19131 => "00000010",19132 => "10110101",19133 => "10101000",19134 => "11011101",19135 => "00111011",19136 => "01100101",19137 => "11100100",19138 => "00010000",19139 => "10001011",19140 => "00010100",19141 => "00001110",19142 => "00011100",19143 => "10001000",19144 => "01111111",19145 => "00001000",19146 => "01101101",19147 => "10000100",19148 => "00110110",19149 => "10001111",19150 => "11001000",19151 => "01101010",19152 => "00010001",19153 => "11010000",19154 => "11011111",19155 => "11101001",19156 => "11010111",19157 => "11011100",19158 => "11011011",19159 => "01101010",19160 => "01101011",19161 => "01111110",19162 => "01110100",19163 => "01110110",19164 => "11000000",19165 => "11001001",19166 => "01001101",19167 => "10111001",19168 => "01000110",19169 => "00110101",19170 => "10110100",19171 => "01110100",19172 => "11100101",19173 => "00000000",19174 => "10001011",19175 => "10011111",19176 => "01111111",19177 => "01101100",19178 => "10001110",19179 => "00101000",19180 => "10110011",19181 => "10101000",19182 => "01111101",19183 => "11100000",19184 => "00110100",19185 => "11100010",19186 => "01011111",19187 => "11110010",19188 => "00101101",19189 => "10011000",19190 => "10001111",19191 => "10001111",19192 => "01100101",19193 => "01110110",19194 => "01001011",19195 => "01000110",19196 => "10000100",19197 => "10110110",19198 => "10001101",19199 => "01000100",19200 => "00011100",19201 => "11000001",19202 => "11010011",19203 => "11100100",19204 => "00011000",19205 => "01100000",19206 => "00010011",19207 => "00100101",19208 => "01010111",19209 => "01010000",19210 => "11111110",19211 => "10100110",19212 => "11101110",19213 => "10100010",19214 => "11111100",19215 => "11110111",19216 => "11111111",19217 => "11110011",19218 => "01111100",19219 => "11011011",19220 => "10100101",19221 => "00011001",19222 => "00101101",19223 => "11010000",19224 => "01001011",19225 => "00010001",19226 => "00011001",19227 => "10000110",19228 => "10001110",19229 => "01100010",19230 => "10010001",19231 => "11100111",19232 => "11010111",19233 => "11011010",19234 => "01001000",19235 => "11100101",19236 => "00110010",19237 => "00110101",19238 => "01010101",19239 => "10101101",19240 => "00101110",19241 => "01110001",19242 => "11001000",19243 => "00011101",19244 => "01101111",19245 => "10001111",19246 => "11010100",19247 => "11101100",19248 => "01010100",19249 => "01100010",19250 => "11111111",19251 => "01001010",19252 => "01010100",19253 => "01011010",19254 => "11010110",19255 => "00110100",19256 => "00111001",19257 => "01101011",19258 => "00101100",19259 => "01010110",19260 => "01101110",19261 => "00101111",19262 => "10000001",19263 => "01000000",19264 => "00100100",19265 => "11011110",19266 => "10111110",19267 => "10111100",19268 => "10011100",19269 => "01000110",19270 => "00101100",19271 => "10111000",19272 => "00000001",19273 => "11010000",19274 => "00010010",19275 => "01001000",19276 => "01101111",19277 => "01110001",19278 => "01000110",19279 => "11100001",19280 => "01100000",19281 => "10010101",19282 => "01111110",19283 => "00000101",19284 => "11010000",19285 => "00110110",19286 => "11000101",19287 => "00100110",19288 => "11011001",19289 => "01011000",19290 => "01000111",19291 => "10000011",19292 => "10011111",19293 => "10110111",19294 => "01111001",19295 => "00111001",19296 => "00110101",19297 => "01000010",19298 => "00111001",19299 => "10110100",19300 => "10010101",19301 => "01101001",19302 => "00111110",19303 => "10111011",19304 => "00000000",19305 => "11001110",19306 => "10100001",19307 => "11110101",19308 => "01001000",19309 => "10101110",19310 => "11001011",19311 => "10010100",19312 => "01000001",19313 => "01000000",19314 => "00101001",19315 => "10100011",19316 => "11100010",19317 => "11110000",19318 => "10000110",19319 => "10000110",19320 => "00101110",19321 => "00001111",19322 => "11100001",19323 => "10100110",19324 => "00011011",19325 => "11110000",19326 => "01001111",19327 => "11111111",19328 => "00111001",19329 => "01111001",19330 => "10100100",19331 => "01110001",19332 => "00010000",19333 => "11001111",19334 => "10110000",19335 => "11011000",19336 => "00010011",19337 => "00110100",19338 => "00011000",19339 => "01001101",19340 => "01111101",19341 => "11111100",19342 => "00010010",19343 => "00100000",19344 => "00010010",19345 => "00000101",19346 => "10001100",19347 => "00101101",19348 => "11110100",19349 => "01111101",19350 => "10101110",19351 => "01011101",19352 => "10100001",19353 => "01110011",19354 => "00001011",19355 => "11011110",19356 => "00110101",19357 => "11010111",19358 => "10010001",19359 => "01100000",19360 => "00111101",19361 => "10000110",19362 => "01110001",19363 => "01011101",19364 => "01111101",19365 => "11111101",19366 => "01101000",19367 => "10001101",19368 => "01011011",19369 => "10011101",19370 => "10011110",19371 => "10010011",19372 => "11000010",19373 => "00000011",19374 => "11100001",19375 => "10011100",19376 => "10100000",19377 => "11000000",19378 => "11100110",19379 => "00010001",19380 => "11010101",19381 => "01001000",19382 => "01000000",19383 => "01011011",19384 => "10011001",19385 => "00100111",19386 => "00101001",19387 => "00011100",19388 => "11111001",19389 => "11010010",19390 => "00011000",19391 => "11110101",19392 => "00000100",19393 => "01110011",19394 => "10100001",19395 => "01101010",19396 => "10001011",19397 => "10111001",19398 => "01111110",19399 => "00101011",19400 => "01010010",19401 => "11111000",19402 => "00110110",19403 => "11011110",19404 => "01010001",19405 => "10001011",19406 => "00110101",19407 => "00100111",19408 => "11001000",19409 => "10001000",19410 => "00010100",19411 => "00011101",19412 => "11010000",19413 => "01000001",19414 => "10001000",19415 => "10001000",19416 => "01000010",19417 => "11000011",19418 => "01001100",19419 => "11001011",19420 => "11101011",19421 => "01101001",19422 => "10100101",19423 => "10010110",19424 => "01000110",19425 => "01100011",19426 => "00101011",19427 => "11111110",19428 => "11001110",19429 => "11001011",19430 => "01000000",19431 => "11011011",19432 => "00010001",19433 => "10000111",19434 => "01111110",19435 => "10010010",19436 => "00000101",19437 => "01110010",19438 => "01010110",19439 => "01100101",19440 => "00010011",19441 => "10000010",19442 => "10010001",19443 => "11010010",19444 => "01010001",19445 => "11100000",19446 => "00110011",19447 => "01010101",19448 => "00111110",19449 => "00110011",19450 => "01001011",19451 => "00010001",19452 => "00101001",19453 => "10100001",19454 => "10111101",19455 => "00110000",19456 => "00000110",19457 => "00111000",19458 => "10011011",19459 => "01001100",19460 => "11001110",19461 => "10010001",19462 => "00001001",19463 => "10010110",19464 => "00100111",19465 => "10010111",19466 => "00000101",19467 => "00011111",19468 => "10111000",19469 => "11001011",19470 => "01001001",19471 => "01101110",19472 => "00000110",19473 => "10000001",19474 => "11111001",19475 => "01000000",19476 => "00111011",19477 => "00001010",19478 => "01110000",19479 => "11000101",19480 => "10001110",19481 => "01000100",19482 => "11011010",19483 => "11100100",19484 => "11101000",19485 => "11010001",19486 => "11110100",19487 => "00100000",19488 => "11010111",19489 => "00111011",19490 => "01100111",19491 => "11000000",19492 => "10011011",19493 => "01101001",19494 => "10011001",19495 => "01110010",19496 => "01001011",19497 => "01010000",19498 => "01001111",19499 => "00111100",19500 => "10001000",19501 => "10010111",19502 => "10001000",19503 => "10101001",19504 => "01010100",19505 => "01110111",19506 => "10011111",19507 => "11111001",19508 => "11110111",19509 => "10000100",19510 => "00111101",19511 => "01010010",19512 => "01010101",19513 => "01001100",19514 => "00101100",19515 => "11000011",19516 => "11011111",19517 => "11110001",19518 => "01101001",19519 => "00001000",19520 => "01101101",19521 => "00010010",19522 => "10000000",19523 => "11110011",19524 => "10100100",19525 => "11010000",19526 => "10010100",19527 => "10010100",19528 => "11111101",19529 => "00111001",19530 => "10011001",19531 => "00001110",19532 => "11110111",19533 => "10111111",19534 => "00010100",19535 => "01110100",19536 => "00011101",19537 => "01101010",19538 => "10111111",19539 => "11011011",19540 => "01101000",19541 => "01011110",19542 => "00001000",19543 => "10101000",19544 => "00011011",19545 => "11101011",19546 => "10111110",19547 => "11011010",19548 => "11101010",19549 => "10010111",19550 => "11000100",19551 => "10100011",19552 => "10010011",19553 => "10001110",19554 => "01001001",19555 => "11001011",19556 => "00100001",19557 => "10000101",19558 => "00110101",19559 => "10000111",19560 => "01110000",19561 => "10011100",19562 => "01101110",19563 => "11100011",19564 => "01001101",19565 => "01101111",19566 => "01001000",19567 => "01100011",19568 => "10110011",19569 => "01101000",19570 => "01111100",19571 => "11101100",19572 => "00001000",19573 => "01000101",19574 => "00100100",19575 => "11110001",19576 => "01010111",19577 => "10011011",19578 => "01100010",19579 => "01011101",19580 => "00000111",19581 => "10011101",19582 => "01101100",19583 => "10110111",19584 => "00000101",19585 => "10111010",19586 => "01001011",19587 => "11000111",19588 => "10000111",19589 => "11100101",19590 => "10010110",19591 => "10110001",19592 => "00100100",19593 => "11100011",19594 => "11100011",19595 => "10001100",19596 => "00100010",19597 => "10001100",19598 => "11110011",19599 => "10101111",19600 => "11011000",19601 => "00000110",19602 => "11011000",19603 => "11011010",19604 => "00011001",19605 => "10000010",19606 => "10111111",19607 => "00001111",19608 => "11001101",19609 => "11001011",19610 => "10001011",19611 => "01010101",19612 => "11011100",19613 => "00111000",19614 => "11001110",19615 => "11100000",19616 => "10011111",19617 => "00001110",19618 => "11000100",19619 => "11001111",19620 => "11010010",19621 => "10001000",19622 => "01110000",19623 => "10100001",19624 => "00101110",19625 => "11010101",19626 => "10000000",19627 => "01101110",19628 => "11110101",19629 => "01000010",19630 => "01101001",19631 => "00110001",19632 => "10011101",19633 => "10001100",19634 => "00011111",19635 => "11110101",19636 => "01101011",19637 => "11010010",19638 => "01001111",19639 => "10100010",19640 => "00111011",19641 => "01011110",19642 => "00101111",19643 => "00010100",19644 => "11011001",19645 => "01001011",19646 => "01100111",19647 => "10101000",19648 => "11011110",19649 => "00101001",19650 => "00110101",19651 => "10100000",19652 => "10101011",19653 => "00100011",19654 => "10000101",19655 => "11011111",19656 => "01111001",19657 => "10101001",19658 => "11111000",19659 => "11001010",19660 => "00011111",19661 => "10011111",19662 => "10000001",19663 => "00110001",19664 => "11111011",19665 => "11110011",19666 => "10000001",19667 => "10000100",19668 => "10100110",19669 => "01111110",19670 => "00011000",19671 => "00100110",19672 => "00010000",19673 => "01011110",19674 => "01111000",19675 => "11111001",19676 => "00101110",19677 => "01110010",19678 => "01011100",19679 => "01000011",19680 => "01001011",19681 => "00011001",19682 => "01010010",19683 => "10001100",19684 => "00110101",19685 => "10000101",19686 => "01110010",19687 => "11101110",19688 => "10100001",19689 => "01110110",19690 => "11010111",19691 => "01010001",19692 => "01110110",19693 => "10010000",19694 => "01101010",19695 => "01110000",19696 => "10001111",19697 => "00001010",19698 => "10000010",19699 => "00111110",19700 => "11100001",19701 => "00100101",19702 => "11101111",19703 => "00111110",19704 => "11000110",19705 => "11100111",19706 => "01000111",19707 => "00100000",19708 => "10101010",19709 => "10100100",19710 => "01011100",19711 => "11110101",19712 => "00011111",19713 => "01100110",19714 => "11111010",19715 => "01100110",19716 => "01111011",19717 => "00000001",19718 => "01010101",19719 => "11011110",19720 => "10000110",19721 => "11110111",19722 => "10111000",19723 => "11000100",19724 => "00011110",19725 => "11010000",19726 => "11010110",19727 => "01110000",19728 => "10100011",19729 => "10011011",19730 => "11000111",19731 => "00001101",19732 => "10100001",19733 => "00001111",19734 => "10010100",19735 => "10000011",19736 => "01001000",19737 => "01000000",19738 => "10000010",19739 => "10101101",19740 => "11011100",19741 => "00010101",19742 => "10101110",19743 => "10110011",19744 => "00101111",19745 => "10110001",19746 => "01101111",19747 => "11110011",19748 => "01010100",19749 => "11110101",19750 => "11010000",19751 => "01100101",19752 => "01101100",19753 => "10100100",19754 => "00011011",19755 => "00110000",19756 => "01011001",19757 => "11001111",19758 => "01100010",19759 => "10110100",19760 => "01011001",19761 => "00011101",19762 => "00010000",19763 => "10111100",19764 => "10111111",19765 => "01111110",19766 => "10110010",19767 => "01110101",19768 => "00100110",19769 => "11101111",19770 => "11001001",19771 => "10010110",19772 => "01000000",19773 => "01101111",19774 => "00000101",19775 => "00110010",19776 => "01001000",19777 => "00111100",19778 => "11010101",19779 => "01100100",19780 => "10111000",19781 => "11100010",19782 => "11001000",19783 => "00011001",19784 => "01110000",19785 => "11110000",19786 => "10011000",19787 => "00101100",19788 => "01010101",19789 => "00111000",19790 => "11010100",19791 => "10111000",19792 => "11100010",19793 => "00101110",19794 => "10001111",19795 => "10110110",19796 => "00001100",19797 => "11001011",19798 => "11111010",19799 => "01000000",19800 => "00001110",19801 => "01000100",19802 => "01011110",19803 => "10010101",19804 => "10011100",19805 => "10111000",19806 => "00110100",19807 => "11011011",19808 => "11001011",19809 => "11000101",19810 => "01001001",19811 => "10001100",19812 => "11101011",19813 => "11111100",19814 => "10000110",19815 => "00101101",19816 => "00000100",19817 => "11010010",19818 => "10101101",19819 => "11010100",19820 => "10000111",19821 => "01001001",19822 => "10111000",19823 => "00110000",19824 => "00011110",19825 => "10011110",19826 => "00110111",19827 => "00001110",19828 => "11011010",19829 => "10101001",19830 => "00111110",19831 => "11100110",19832 => "10111010",19833 => "01011011",19834 => "00111011",19835 => "01010100",19836 => "01000001",19837 => "10100101",19838 => "11011010",19839 => "00010100",19840 => "11111110",19841 => "11011100",19842 => "11101101",19843 => "01011000",19844 => "10100010",19845 => "11110001",19846 => "01110000",19847 => "00111010",19848 => "00000011",19849 => "10111111",19850 => "00010000",19851 => "01010111",19852 => "10111001",19853 => "01001111",19854 => "00011011",19855 => "10111011",19856 => "01000011",19857 => "01010011",19858 => "11011101",19859 => "01101010",19860 => "00000000",19861 => "01101101",19862 => "00100110",19863 => "10011010",19864 => "10101110",19865 => "10010100",19866 => "10001010",19867 => "10100100",19868 => "01100000",19869 => "10101101",19870 => "01110110",19871 => "01110010",19872 => "00111111",19873 => "10010001",19874 => "10000000",19875 => "10001010",19876 => "01011100",19877 => "00010100",19878 => "10101101",19879 => "00100001",19880 => "10010011",19881 => "01001010",19882 => "10000011",19883 => "00011101",19884 => "10101011",19885 => "10010111",19886 => "01010101",19887 => "00011010",19888 => "10001010",19889 => "01000101",19890 => "11111101",19891 => "00101100",19892 => "01111000",19893 => "11011110",19894 => "11001111",19895 => "00011011",19896 => "11101011",19897 => "11001001",19898 => "01000001",19899 => "10011010",19900 => "00100110",19901 => "00100000",19902 => "01100100",19903 => "11100101",19904 => "01010111",19905 => "10010101",19906 => "00010110",19907 => "00001000",19908 => "10111111",19909 => "00100000",19910 => "01111010",19911 => "00101100",19912 => "01000101",19913 => "10001110",19914 => "10001100",19915 => "10000000",19916 => "00111010",19917 => "00101100",19918 => "10101100",19919 => "11100110",19920 => "10100011",19921 => "11111011",19922 => "00100100",19923 => "11011110",19924 => "11000111",19925 => "11101111",19926 => "11001110",19927 => "01111110",19928 => "01010110",19929 => "11011101",19930 => "11101000",19931 => "10010000",19932 => "01100101",19933 => "00011000",19934 => "00000100",19935 => "10100010",19936 => "00000111",19937 => "10111111",19938 => "10010100",19939 => "00010010",19940 => "00010101",19941 => "00001111",19942 => "11010110",19943 => "01100011",19944 => "11111111",19945 => "00110111",19946 => "00100010",19947 => "10010111",19948 => "01010001",19949 => "01011011",19950 => "00100101",19951 => "01111010",19952 => "11010010",19953 => "11010111",19954 => "11100110",19955 => "10101111",19956 => "10001110",19957 => "10110001",19958 => "11000100",19959 => "10001111",19960 => "01010000",19961 => "00000110",19962 => "00110000",19963 => "00001011",19964 => "00011001",19965 => "00010111",19966 => "10001001",19967 => "01001000",19968 => "10000001",19969 => "00111010",19970 => "11100001",19971 => "01011100",19972 => "01111111",19973 => "01010011",19974 => "10111000",19975 => "01101001",19976 => "10010100",19977 => "01010001",19978 => "00010111",19979 => "01001010",19980 => "11000111",19981 => "01001111",19982 => "10110000",19983 => "10111011",19984 => "00100001",19985 => "10011101",19986 => "01100111",19987 => "00110111",19988 => "00110011",19989 => "10000101",19990 => "01101010",19991 => "11110000",19992 => "11000111",19993 => "01010111",19994 => "01010101",19995 => "10010000",19996 => "00000100",19997 => "01000100",19998 => "00001000",19999 => "10101110",20000 => "00001101",20001 => "11110101",20002 => "10111000",20003 => "10110001",20004 => "00101111",20005 => "01000101",20006 => "00110111",20007 => "00111111",20008 => "11111110",20009 => "01111011",20010 => "11000010",20011 => "10111001",20012 => "01110110",20013 => "01010100",20014 => "01001111",20015 => "10001100",20016 => "00011001",20017 => "11111110",20018 => "00111010",20019 => "01010100",20020 => "00101011",20021 => "01110011",20022 => "10010000",20023 => "10101010",20024 => "00101010",20025 => "01111011",20026 => "11001100",20027 => "10000000",20028 => "01101111",20029 => "00000101",20030 => "11111100",20031 => "00101101",20032 => "00101001",20033 => "10010100",20034 => "11010100",20035 => "00110010",20036 => "00000001",20037 => "01101011",20038 => "01110100",20039 => "00001000",20040 => "11011001",20041 => "01110011",20042 => "10111001",20043 => "11000011",20044 => "11111100",20045 => "10110000",20046 => "01110010",20047 => "10110011",20048 => "11000010",20049 => "00110001",20050 => "01110011",20051 => "10001101",20052 => "11100010",20053 => "10000001",20054 => "00010101",20055 => "11001000",20056 => "10110101",20057 => "00011000",20058 => "11011100",20059 => "01101000",20060 => "11110000",20061 => "00000001",20062 => "10100001",20063 => "00001101",20064 => "11010000",20065 => "00011111",20066 => "10101000",20067 => "00000111",20068 => "11110000",20069 => "01100011",20070 => "10001111",20071 => "11001100",20072 => "10010110",20073 => "01011111",20074 => "01111010",20075 => "11101100",20076 => "00111100",20077 => "00110011",20078 => "01110000",20079 => "01000100",20080 => "11101110",20081 => "01100010",20082 => "11010100",20083 => "01000000",20084 => "00111001",20085 => "00000001",20086 => "00011110",20087 => "01001110",20088 => "11101010",20089 => "00111100",20090 => "00101101",20091 => "10010000",20092 => "00001000",20093 => "10010111",20094 => "11100011",20095 => "01001110",20096 => "10011000",20097 => "11111101",20098 => "00000000",20099 => "00011100",20100 => "11111110",20101 => "10111010",20102 => "01010111",20103 => "00110101",20104 => "10111011",20105 => "00110100",20106 => "10010111",20107 => "11001101",20108 => "00001100",20109 => "11101101",20110 => "11001010",20111 => "10110111",20112 => "01001110",20113 => "00101111",20114 => "01111010",20115 => "00000101",20116 => "10001001",20117 => "11101010",20118 => "11010011",20119 => "11110010",20120 => "01101001",20121 => "10011001",20122 => "00101100",20123 => "01101101",20124 => "10010011",20125 => "00100111",20126 => "00101111",20127 => "00101010",20128 => "11010010",20129 => "10011011",20130 => "01111100",20131 => "00011100",20132 => "00100001",20133 => "01101001",20134 => "10000001",20135 => "10000011",20136 => "11011111",20137 => "00000011",20138 => "11110110",20139 => "01100101",20140 => "11100111",20141 => "00110101",20142 => "00011101",20143 => "01001001",20144 => "00100001",20145 => "01100100",20146 => "01010001",20147 => "10100100",20148 => "01011111",20149 => "01100011",20150 => "11010111",20151 => "00100110",20152 => "00101110",20153 => "00101101",20154 => "01100100",20155 => "10101010",20156 => "00111110",20157 => "10110000",20158 => "10110000",20159 => "11110010",20160 => "01001000",20161 => "10010101",20162 => "11011001",20163 => "11110000",20164 => "11000110",20165 => "00100100",20166 => "00111010",20167 => "10010001",20168 => "00001011",20169 => "10001001",20170 => "00110011",20171 => "11001000",20172 => "11101111",20173 => "01111000",20174 => "00011010",20175 => "00100111",20176 => "11110100",20177 => "01010000",20178 => "01100111",20179 => "10010110",20180 => "01011100",20181 => "11001000",20182 => "11000101",20183 => "00011100",20184 => "11101111",20185 => "01011010",20186 => "11110001",20187 => "00100011",20188 => "10001000",20189 => "00111000",20190 => "11101011",20191 => "11001111",20192 => "11100000",20193 => "11111101",20194 => "00100000",20195 => "01110110",20196 => "11001011",20197 => "10101111",20198 => "01011010",20199 => "00011000",20200 => "10100110",20201 => "01110111",20202 => "01111101",20203 => "11110001",20204 => "01001110",20205 => "11101011",20206 => "10100110",20207 => "11111011",20208 => "00100001",20209 => "00001100",20210 => "10011110",20211 => "00100011",20212 => "10011101",20213 => "01011001",20214 => "10010100",20215 => "11110001",20216 => "01010000",20217 => "00100111",20218 => "01001011",20219 => "11110010",20220 => "10010000",20221 => "11100000",20222 => "10001011",20223 => "00010001",20224 => "01011000",20225 => "01110001",20226 => "11001110",20227 => "00101110",20228 => "01011011",20229 => "10110110",20230 => "10100001",20231 => "10011010",20232 => "00100111",20233 => "01010110",20234 => "01001010",20235 => "10011010",20236 => "00110000",20237 => "00001101",20238 => "11000101",20239 => "01001100",20240 => "11001101",20241 => "01001001",20242 => "11010010",20243 => "01111100",20244 => "01111000",20245 => "10010001",20246 => "01101111",20247 => "01001011",20248 => "01000011",20249 => "11111101",20250 => "01000110",20251 => "11101100",20252 => "10010001",20253 => "10111100",20254 => "01001011",20255 => "00011010",20256 => "01000011",20257 => "01110110",20258 => "01010000",20259 => "11001000",20260 => "10100111",20261 => "10100000",20262 => "00110110",20263 => "00010011",20264 => "11010110",20265 => "11111010",20266 => "00010011",20267 => "11001010",20268 => "11100011",20269 => "10111010",20270 => "00101111",20271 => "11001110",20272 => "11100100",20273 => "01010000",20274 => "00110110",20275 => "10011011",20276 => "10110101",20277 => "01110111",20278 => "10011001",20279 => "11100011",20280 => "10001010",20281 => "00111111",20282 => "01111101",20283 => "11110001",20284 => "10100110",20285 => "11101110",20286 => "00010111",20287 => "10000101",20288 => "10000000",20289 => "11011101",20290 => "00100101",20291 => "01010011",20292 => "01001000",20293 => "00011010",20294 => "11011111",20295 => "00101000",20296 => "01111010",20297 => "10111011",20298 => "01110100",20299 => "10110000",20300 => "11010110",20301 => "00110110",20302 => "00101011",20303 => "11101101",20304 => "11100011",20305 => "11100110",20306 => "00110100",20307 => "10111111",20308 => "10001100",20309 => "01111101",20310 => "11100110",20311 => "01001000",20312 => "11001111",20313 => "00010110",20314 => "10100001",20315 => "00000011",20316 => "01000110",20317 => "11001101",20318 => "00111000",20319 => "11100100",20320 => "11111001",20321 => "00000110",20322 => "10000011",20323 => "11101010",20324 => "11110110",20325 => "10001010",20326 => "01100010",20327 => "00011011",20328 => "11011100",20329 => "11110111",20330 => "11011101",20331 => "01000011",20332 => "11110001",20333 => "01111010",20334 => "10110101",20335 => "10001110",20336 => "01011100",20337 => "11110010",20338 => "11111010",20339 => "01100010",20340 => "11110111",20341 => "00110100",20342 => "11010101",20343 => "11110110",20344 => "10111011",20345 => "11110001",20346 => "11010101",20347 => "00011010",20348 => "10111011",20349 => "00101100",20350 => "01010011",20351 => "11001011",20352 => "10011111",20353 => "01110100",20354 => "10001110",20355 => "01101010",20356 => "01111011",20357 => "10111000",20358 => "00000110",20359 => "01111000",20360 => "00101101",20361 => "01101101",20362 => "10101101",20363 => "00011101",20364 => "11101001",20365 => "10010101",20366 => "01001001",20367 => "01100010",20368 => "00011100",20369 => "11101011",20370 => "11011010",20371 => "00011110",20372 => "01111010",20373 => "10011011",20374 => "01001001",20375 => "00011100",20376 => "00111011",20377 => "01010111",20378 => "11001011",20379 => "11110011",20380 => "10110010",20381 => "10101100",20382 => "01010000",20383 => "11100101",20384 => "10110001",20385 => "11101011",20386 => "11111111",20387 => "00111011",20388 => "11001100",20389 => "10111010",20390 => "11110111",20391 => "00010001",20392 => "01111101",20393 => "00010001",20394 => "11010000",20395 => "10111011",20396 => "11001111",20397 => "01101001",20398 => "11011000",20399 => "10110001",20400 => "11100110",20401 => "10001100",20402 => "01010110",20403 => "01101111",20404 => "11010100",20405 => "00100000",20406 => "00101100",20407 => "10111010",20408 => "10100101",20409 => "10100100",20410 => "00110100",20411 => "10000000",20412 => "00001010",20413 => "00111100",20414 => "11100010",20415 => "11010101",20416 => "11000101",20417 => "10100100",20418 => "00110101",20419 => "11000100",20420 => "11110001",20421 => "10101011",20422 => "01001001",20423 => "11111011",20424 => "01100000",20425 => "01100111",20426 => "01100101",20427 => "00101110",20428 => "11001010",20429 => "11110010",20430 => "10101100",20431 => "10001101",20432 => "10111001",20433 => "01011110",20434 => "11110000",20435 => "00110101",20436 => "00010000",20437 => "10110000",20438 => "11101010",20439 => "00111100",20440 => "10000110",20441 => "00010111",20442 => "11101100",20443 => "00101010",20444 => "10001001",20445 => "10000000",20446 => "01111001",20447 => "10110111",20448 => "11100001",20449 => "00011011",20450 => "01011000",20451 => "10001110",20452 => "00110111",20453 => "01000111",20454 => "01111111",20455 => "00011010",20456 => "10001010",20457 => "01010001",20458 => "11010000",20459 => "00001111",20460 => "00011011",20461 => "00100100",20462 => "01000010",20463 => "00010110",20464 => "10000101",20465 => "00000000",20466 => "11011100",20467 => "01011111",20468 => "00110011",20469 => "00111110",20470 => "00101101",20471 => "00111001",20472 => "10000110",20473 => "01111011",20474 => "10010010",20475 => "01010110",20476 => "10001001",20477 => "01010001",20478 => "01110011",20479 => "11011011",20480 => "01101111",20481 => "00000111",20482 => "01111111",20483 => "00000101",20484 => "01110010",20485 => "10100101",20486 => "10110000",20487 => "01011000",20488 => "11010001",20489 => "00010101",20490 => "00010010",20491 => "01001001",20492 => "11001011",20493 => "10011000",20494 => "00000010",20495 => "01001101",20496 => "10111111",20497 => "01100001",20498 => "01001010",20499 => "01010111",20500 => "01101100",20501 => "10000011",20502 => "00001111",20503 => "00111111",20504 => "00101100",20505 => "00101111",20506 => "11001100",20507 => "01011001",20508 => "11010010",20509 => "11100110",20510 => "10011000",20511 => "10000001",20512 => "01111101",20513 => "10101101",20514 => "10111110",20515 => "10000001",20516 => "00100001",20517 => "00111111",20518 => "11111000",20519 => "11010110",20520 => "11111110",20521 => "00011001",20522 => "00110011",20523 => "11100001",20524 => "00011011",20525 => "00011010",20526 => "11111001",20527 => "10000011",20528 => "01001000",20529 => "00111110",20530 => "10100010",20531 => "00110010",20532 => "01000010",20533 => "11110010",20534 => "00001111",20535 => "11101010",20536 => "11101000",20537 => "10001000",20538 => "00111011",20539 => "01111001",20540 => "11110001",20541 => "01000011",20542 => "11111001",20543 => "11110110",20544 => "00000100",20545 => "00110000",20546 => "01001010",20547 => "00011110",20548 => "01001011",20549 => "00000011",20550 => "00001011",20551 => "10011101",20552 => "11010100",20553 => "00011100",20554 => "00010100",20555 => "01010111",20556 => "10100110",20557 => "01111010",20558 => "10111111",20559 => "11100011",20560 => "00011000",20561 => "10110100",20562 => "01110111",20563 => "11101001",20564 => "10100100",20565 => "10101001",20566 => "11000111",20567 => "10000100",20568 => "10010110",20569 => "01110001",20570 => "01000100",20571 => "01000100",20572 => "00111101",20573 => "00011000",20574 => "01011010",20575 => "10110110",20576 => "11010000",20577 => "01100000",20578 => "01010100",20579 => "01100010",20580 => "00101001",20581 => "10011110",20582 => "10000111",20583 => "11000000",20584 => "00000100",20585 => "10001111",20586 => "01011100",20587 => "01100101",20588 => "01111100",20589 => "11011010",20590 => "11011111",20591 => "11000001",20592 => "10000010",20593 => "10110010",20594 => "00101101",20595 => "00001101",20596 => "00101110",20597 => "00111000",20598 => "11001100",20599 => "00010011",20600 => "00101111",20601 => "01000111",20602 => "01011010",20603 => "01010010",20604 => "10111000",20605 => "11100001",20606 => "11001010",20607 => "00100110",20608 => "11011111",20609 => "00110010",20610 => "11100100",20611 => "00011000",20612 => "11001100",20613 => "00110001",20614 => "01110101",20615 => "01110110",20616 => "00001100",20617 => "10101111",20618 => "11110001",20619 => "10110011",20620 => "10000001",20621 => "10100100",20622 => "10011111",20623 => "11011100",20624 => "01001110",20625 => "11010110",20626 => "00110110",20627 => "10101001",20628 => "10001100",20629 => "00111110",20630 => "01000100",20631 => "11111101",20632 => "00100010",20633 => "01010111",20634 => "10011100",20635 => "11001101",20636 => "00001101",20637 => "10000000",20638 => "00110110",20639 => "11100010",20640 => "00100100",20641 => "01101000",20642 => "01011111",20643 => "10000001",20644 => "11110110",20645 => "10101010",20646 => "00011010",20647 => "00000111",20648 => "11011001",20649 => "10011110",20650 => "00001010",20651 => "11100001",20652 => "01110011",20653 => "00000011",20654 => "10000011",20655 => "10100111",20656 => "11011010",20657 => "11100111",20658 => "10101111",20659 => "11000010",20660 => "00011100",20661 => "10000110",20662 => "11000001",20663 => "10000111",20664 => "11001111",20665 => "00110101",20666 => "01101001",20667 => "11000100",20668 => "11111001",20669 => "10001100",20670 => "11110101",20671 => "10100011",20672 => "11001100",20673 => "01001000",20674 => "01100111",20675 => "10101111",20676 => "00110000",20677 => "00101100",20678 => "00111001",20679 => "10010100",20680 => "00100000",20681 => "01110001",20682 => "10101011",20683 => "00000011",20684 => "00010111",20685 => "01010010",20686 => "00101011",20687 => "01011111",20688 => "01100011",20689 => "10010011",20690 => "00010001",20691 => "11000111",20692 => "01010110",20693 => "10111010",20694 => "01001111",20695 => "00001110",20696 => "11100100",20697 => "01101000",20698 => "10010010",20699 => "10101010",20700 => "01001110",20701 => "11011101",20702 => "11110011",20703 => "00100010",20704 => "01100011",20705 => "10111011",20706 => "10100011",20707 => "10111101",20708 => "01011000",20709 => "01001000",20710 => "10010011",20711 => "11101101",20712 => "10010101",20713 => "10111111",20714 => "01100110",20715 => "01000000",20716 => "10000101",20717 => "01110010",20718 => "00010010",20719 => "10110101",20720 => "10111110",20721 => "11010110",20722 => "00010111",20723 => "00110010",20724 => "00110101",20725 => "00011111",20726 => "01100000",20727 => "10111011",20728 => "01100110",20729 => "01000010",20730 => "01101110",20731 => "10110101",20732 => "10100110",20733 => "00011011",20734 => "00111100",20735 => "01110011",20736 => "00010111",20737 => "00011100",20738 => "00111000",20739 => "11011111",20740 => "11101111",20741 => "00000100",20742 => "10000010",20743 => "11101101",20744 => "11010000",20745 => "11100011",20746 => "11010011",20747 => "11010101",20748 => "00000011",20749 => "01101010",20750 => "11001111",20751 => "00101111",20752 => "00010010",20753 => "00110001",20754 => "00001011",20755 => "11111011",20756 => "11000111",20757 => "01111110",20758 => "11111110",20759 => "11110001",20760 => "00000100",20761 => "00101010",20762 => "01000100",20763 => "10101100",20764 => "01101101",20765 => "10111110",20766 => "01010101",20767 => "10100100",20768 => "00100011",20769 => "00111111",20770 => "00110101",20771 => "00110111",20772 => "00100010",20773 => "01000011",20774 => "11001010",20775 => "11110101",20776 => "11100001",20777 => "11001110",20778 => "01011101",20779 => "11110010",20780 => "00001001",20781 => "10011001",20782 => "10000111",20783 => "01000000",20784 => "01010001",20785 => "10100111",20786 => "10110100",20787 => "01110110",20788 => "11011000",20789 => "11101010",20790 => "10110110",20791 => "11100000",20792 => "00001011",20793 => "11101001",20794 => "00110110",20795 => "11000101",20796 => "11100010",20797 => "01111110",20798 => "01001001",20799 => "11101011",20800 => "01000101",20801 => "11101111",20802 => "01010011",20803 => "00101000",20804 => "10110001",20805 => "10101011",20806 => "10111000",20807 => "01000110",20808 => "00010100",20809 => "10100101",20810 => "00111011",20811 => "00101111",20812 => "10110011",20813 => "10110111",20814 => "10110000",20815 => "01001100",20816 => "11101111",20817 => "11100111",20818 => "10101110",20819 => "00110011",20820 => "00010111",20821 => "00110000",20822 => "11001011",20823 => "10010101",20824 => "11111110",20825 => "01101110",20826 => "01101000",20827 => "10000110",20828 => "01111011",20829 => "10001101",20830 => "11100010",20831 => "00001000",20832 => "00011010",20833 => "10000100",20834 => "10101001",20835 => "00110010",20836 => "10111111",20837 => "01000011",20838 => "11111111",20839 => "01011000",20840 => "00010100",20841 => "01010010",20842 => "00111111",20843 => "00010111",20844 => "01101111",20845 => "00110010",20846 => "10100010",20847 => "00000111",20848 => "01111000",20849 => "00010110",20850 => "01101010",20851 => "01001011",20852 => "00001001",20853 => "00111110",20854 => "01101101",20855 => "10101011",20856 => "10111000",20857 => "00111111",20858 => "01010010",20859 => "10110001",20860 => "01110100",20861 => "10011101",20862 => "01010011",20863 => "01001011",20864 => "01000111",20865 => "11000001",20866 => "11001010",20867 => "11100011",20868 => "10110000",20869 => "11110111",20870 => "10000110",20871 => "11001010",20872 => "01000100",20873 => "01000101",20874 => "11111011",20875 => "11111001",20876 => "11110111",20877 => "10111101",20878 => "10000100",20879 => "10000101",20880 => "01111101",20881 => "10100111",20882 => "00110011",20883 => "00011001",20884 => "10101011",20885 => "11100110",20886 => "11010001",20887 => "01010110",20888 => "11110111",20889 => "01110111",20890 => "10010000",20891 => "11000100",20892 => "01011010",20893 => "10000001",20894 => "10010101",20895 => "10101001",20896 => "00110110",20897 => "11111100",20898 => "11110001",20899 => "11010110",20900 => "10111110",20901 => "00010100",20902 => "00010111",20903 => "01010101",20904 => "01001101",20905 => "11101011",20906 => "00111101",20907 => "10101000",20908 => "01111010",20909 => "10111101",20910 => "01010001",20911 => "01100111",20912 => "00110110",20913 => "01100000",20914 => "00101111",20915 => "11111001",20916 => "10001000",20917 => "10010010",20918 => "11000010",20919 => "10011100",20920 => "11111111",20921 => "01110010",20922 => "10100111",20923 => "11000101",20924 => "00011010",20925 => "11110011",20926 => "00011001",20927 => "00001000",20928 => "11010010",20929 => "00010011",20930 => "01000111",20931 => "01001110",20932 => "11101100",20933 => "00001110",20934 => "10001101",20935 => "00000010",20936 => "11100010",20937 => "00101110",20938 => "00100101",20939 => "00000001",20940 => "11100010",20941 => "00101100",20942 => "01001100",20943 => "01010101",20944 => "11011100",20945 => "10011001",20946 => "10110110",20947 => "01101010",20948 => "10000101",20949 => "11011111",20950 => "00001011",20951 => "10110010",20952 => "10011100",20953 => "01000100",20954 => "10110010",20955 => "00010000",20956 => "10110100",20957 => "10101010",20958 => "10010101",20959 => "10001010",20960 => "11001010",20961 => "01100000",20962 => "11110111",20963 => "00100011",20964 => "10110010",20965 => "00001001",20966 => "11111011",20967 => "11010110",20968 => "01101010",20969 => "00000010",20970 => "10110101",20971 => "01111110",20972 => "11000100",20973 => "11110111",20974 => "10010111",20975 => "00001001",20976 => "11000111",20977 => "10000111",20978 => "11100000",20979 => "01100000",20980 => "01111110",20981 => "00100011",20982 => "00010111",20983 => "10001011",20984 => "01110000",20985 => "10100010",20986 => "10101011",20987 => "11011000",20988 => "01100100",20989 => "00000000",20990 => "00010001",20991 => "11100001",20992 => "00111010",20993 => "00000010",20994 => "00010101",20995 => "10001001",20996 => "01110000",20997 => "01110010",20998 => "10101111",20999 => "01100101",21000 => "01010011",21001 => "11001001",21002 => "01101101",21003 => "11101101",21004 => "11110011",21005 => "10000111",21006 => "01001110",21007 => "00000101",21008 => "11110100",21009 => "11111010",21010 => "10000011",21011 => "00111110",21012 => "00001011",21013 => "01100001",21014 => "01100110",21015 => "10000111",21016 => "11010101",21017 => "11010100",21018 => "00010100",21019 => "10010001",21020 => "10011011",21021 => "11110010",21022 => "01000000",21023 => "01001010",21024 => "11000000",21025 => "00101100",21026 => "01001100",21027 => "00000111",21028 => "10111111",21029 => "01111000",21030 => "11101010",21031 => "01010001",21032 => "11111110",21033 => "10011001",21034 => "01110001",21035 => "00001000",21036 => "01110011",21037 => "00001101",21038 => "10001100",21039 => "10111010",21040 => "11110001",21041 => "01101110",21042 => "10111010",21043 => "01011011",21044 => "01110100",21045 => "11001011",21046 => "01100110",21047 => "01101010",21048 => "11110000",21049 => "10101001",21050 => "00010000",21051 => "10101110",21052 => "11100100",21053 => "10001001",21054 => "00011100",21055 => "10111011",21056 => "11111011",21057 => "10001111",21058 => "01101100",21059 => "11101110",21060 => "10010101",21061 => "11000011",21062 => "01101010",21063 => "11111101",21064 => "10010000",21065 => "00101101",21066 => "00010001",21067 => "00000100",21068 => "11100100",21069 => "00001110",21070 => "00111000",21071 => "11000100",21072 => "10111000",21073 => "01101110",21074 => "11010110",21075 => "01011100",21076 => "11001110",21077 => "11110110",21078 => "10110001",21079 => "00000111",21080 => "01000100",21081 => "01110010",21082 => "10000101",21083 => "01111110",21084 => "10011011",21085 => "01100000",21086 => "00101011",21087 => "11010110",21088 => "10000110",21089 => "01101101",21090 => "11110101",21091 => "10010010",21092 => "00000111",21093 => "11000110",21094 => "01000110",21095 => "10011001",21096 => "01110000",21097 => "00100010",21098 => "10100101",21099 => "00101010",21100 => "01101010",21101 => "00101101",21102 => "01110001",21103 => "01110000",21104 => "00011001",21105 => "01101010",21106 => "01110101",21107 => "00000101",21108 => "01111011",21109 => "11111101",21110 => "10100001",21111 => "10111011",21112 => "01011101",21113 => "01101100",21114 => "01001110",21115 => "11111000",21116 => "11110111",21117 => "10001001",21118 => "01000100",21119 => "00000110",21120 => "00010110",21121 => "11010110",21122 => "10010100",21123 => "11110011",21124 => "01111000",21125 => "10011111",21126 => "01000101",21127 => "01011101",21128 => "01110101",21129 => "11110110",21130 => "10101100",21131 => "00100100",21132 => "00000010",21133 => "11101010",21134 => "10011010",21135 => "10100011",21136 => "10011111",21137 => "10000011",21138 => "10010100",21139 => "11110000",21140 => "11111100",21141 => "10010011",21142 => "10101110",21143 => "01101010",21144 => "10100010",21145 => "01101000",21146 => "00001101",21147 => "11111111",21148 => "11100100",21149 => "10010100",21150 => "11101001",21151 => "00110001",21152 => "00101000",21153 => "01110110",21154 => "01101001",21155 => "00011001",21156 => "11100010",21157 => "11100100",21158 => "01101101",21159 => "11011100",21160 => "00000010",21161 => "00111010",21162 => "01100010",21163 => "11100100",21164 => "10001111",21165 => "10011100",21166 => "01000110",21167 => "01110010",21168 => "10110000",21169 => "01011110",21170 => "01111110",21171 => "01001001",21172 => "11101001",21173 => "11101111",21174 => "01001101",21175 => "10110111",21176 => "10111010",21177 => "01110101",21178 => "10001100",21179 => "01001111",21180 => "00100001",21181 => "10011100",21182 => "01011001",21183 => "10011000",21184 => "11011111",21185 => "11111011",21186 => "01110010",21187 => "01000110",21188 => "00100011",21189 => "11100001",21190 => "10100111",21191 => "00110110",21192 => "01000000",21193 => "11100010",21194 => "10000100",21195 => "01010110",21196 => "00100001",21197 => "11100101",21198 => "10110010",21199 => "00000001",21200 => "00010100",21201 => "11001110",21202 => "01101111",21203 => "00100111",21204 => "01110001",21205 => "01101111",21206 => "01011000",21207 => "10011001",21208 => "10111100",21209 => "01011000",21210 => "11110011",21211 => "00001010",21212 => "00110111",21213 => "10011110",21214 => "10111101",21215 => "10011011",21216 => "00100001",21217 => "01010010",21218 => "11000010",21219 => "11001100",21220 => "01110000",21221 => "00001110",21222 => "00110110",21223 => "11010011",21224 => "10100001",21225 => "11001000",21226 => "11100001",21227 => "11001011",21228 => "01111011",21229 => "11011111",21230 => "11111010",21231 => "01101101",21232 => "01111001",21233 => "11010011",21234 => "01011100",21235 => "00101010",21236 => "00001111",21237 => "01111110",21238 => "10111110",21239 => "11000111",21240 => "10111000",21241 => "00000100",21242 => "10000010",21243 => "10000011",21244 => "00000101",21245 => "01010101",21246 => "01011001",21247 => "11110100",21248 => "11100101",21249 => "11011111",21250 => "10001110",21251 => "00010100",21252 => "00100001",21253 => "01101000",21254 => "00110110",21255 => "00100100",21256 => "10010100",21257 => "01100000",21258 => "10111000",21259 => "10010100",21260 => "10111111",21261 => "10010010",21262 => "01001100",21263 => "11010011",21264 => "10001100",21265 => "00001000",21266 => "01111100",21267 => "01111000",21268 => "11101100",21269 => "11011110",21270 => "10100110",21271 => "11010100",21272 => "00101010",21273 => "11001000",21274 => "10100001",21275 => "00101111",21276 => "01000101",21277 => "01000100",21278 => "11111101",21279 => "10111100",21280 => "00010101",21281 => "00011001",21282 => "11110000",21283 => "11101000",21284 => "11101100",21285 => "11001010",21286 => "00100110",21287 => "11111101",21288 => "11010011",21289 => "00101010",21290 => "11011010",21291 => "01011011",21292 => "01110101",21293 => "01110101",21294 => "11110111",21295 => "00000101",21296 => "01101011",21297 => "10000011",21298 => "10101011",21299 => "01000101",21300 => "11011110",21301 => "10101010",21302 => "00100101",21303 => "10010001",21304 => "01110111",21305 => "11010011",21306 => "10011000",21307 => "11010110",21308 => "10011110",21309 => "01100010",21310 => "10111001",21311 => "10111100",21312 => "01000011",21313 => "11101111",21314 => "10010111",21315 => "10101010",21316 => "01100001",21317 => "01110001",21318 => "00101000",21319 => "00110111",21320 => "11000110",21321 => "00100000",21322 => "11011110",21323 => "00110001",21324 => "01011001",21325 => "11011100",21326 => "00010100",21327 => "01101011",21328 => "01110110",21329 => "11100100",21330 => "00001111",21331 => "11001110",21332 => "10011010",21333 => "00110110",21334 => "00110011",21335 => "10101001",21336 => "00000101",21337 => "01001101",21338 => "10101001",21339 => "01001101",21340 => "10100001",21341 => "11001101",21342 => "01100010",21343 => "11010100",21344 => "00111010",21345 => "01001110",21346 => "10001100",21347 => "10010110",21348 => "01100000",21349 => "10000110",21350 => "01011000",21351 => "01111101",21352 => "10000011",21353 => "11101110",21354 => "00000001",21355 => "00110010",21356 => "00010111",21357 => "00100000",21358 => "11011100",21359 => "11001101",21360 => "00011110",21361 => "11111010",21362 => "01111100",21363 => "01010011",21364 => "11011001",21365 => "11011110",21366 => "11100111",21367 => "11101101",21368 => "10011101",21369 => "11110111",21370 => "00010101",21371 => "00101111",21372 => "01101001",21373 => "00000110",21374 => "01000101",21375 => "11001101",21376 => "01111101",21377 => "11000000",21378 => "00111110",21379 => "10001010",21380 => "00010100",21381 => "00000011",21382 => "11101110",21383 => "01010001",21384 => "00001011",21385 => "01111100",21386 => "00100011",21387 => "11011001",21388 => "00111000",21389 => "00011001",21390 => "11001111",21391 => "01011110",21392 => "10100100",21393 => "01000110",21394 => "01011000",21395 => "01011011",21396 => "00111011",21397 => "01001101",21398 => "11101111",21399 => "00100000",21400 => "00100100",21401 => "11001101",21402 => "01110100",21403 => "00100010",21404 => "11100010",21405 => "10111011",21406 => "11101011",21407 => "11100011",21408 => "10100110",21409 => "01001000",21410 => "00011011",21411 => "11110000",21412 => "00110011",21413 => "10100111",21414 => "00011100",21415 => "11010100",21416 => "11101011",21417 => "00011110",21418 => "00101100",21419 => "00001001",21420 => "10101011",21421 => "01110011",21422 => "01010000",21423 => "11010100",21424 => "11000111",21425 => "00011011",21426 => "11001100",21427 => "01101101",21428 => "00011101",21429 => "11101000",21430 => "10111011",21431 => "10000011",21432 => "00010110",21433 => "11010110",21434 => "00010000",21435 => "00011001",21436 => "11110000",21437 => "10111001",21438 => "01111010",21439 => "00110010",21440 => "10011001",21441 => "10110011",21442 => "00000111",21443 => "11010101",21444 => "11001001",21445 => "00000000",21446 => "10110000",21447 => "11001111",21448 => "01100010",21449 => "10100000",21450 => "10010100",21451 => "11100100",21452 => "01001101",21453 => "01110000",21454 => "00100111",21455 => "01100111",21456 => "10011110",21457 => "11000000",21458 => "01001011",21459 => "00110010",21460 => "10111100",21461 => "01110100",21462 => "01011011",21463 => "11010110",21464 => "01010111",21465 => "00100000",21466 => "00110001",21467 => "01011011",21468 => "01011110",21469 => "11111001",21470 => "01000101",21471 => "00101011",21472 => "00000001",21473 => "01111001",21474 => "10001110",21475 => "10111001",21476 => "10011001",21477 => "11000010",21478 => "10100101",21479 => "11010110",21480 => "00110101",21481 => "00010110",21482 => "01000000",21483 => "01011111",21484 => "00110000",21485 => "01010010",21486 => "01100100",21487 => "10001100",21488 => "10101100",21489 => "00101001",21490 => "00011111",21491 => "01000011",21492 => "11111101",21493 => "00111110",21494 => "00001110",21495 => "11111010",21496 => "11100000",21497 => "00111011",21498 => "01100111",21499 => "10010000",21500 => "11010110",21501 => "11000101",21502 => "01011110",21503 => "11001111",21504 => "10110001",21505 => "10100011",21506 => "11010010",21507 => "01101011",21508 => "01101011",21509 => "01100110",21510 => "00100100",21511 => "10010101",21512 => "11110101",21513 => "11100011",21514 => "11101001",21515 => "11001011",21516 => "10010111",21517 => "01001101",21518 => "00000000",21519 => "00100110",21520 => "11001100",21521 => "11101011",21522 => "01100010",21523 => "11110010",21524 => "11110011",21525 => "00001001",21526 => "11100111",21527 => "00011101",21528 => "10111101",21529 => "11001101",21530 => "00001110",21531 => "01011110",21532 => "11000110",21533 => "11011010",21534 => "11000110",21535 => "00010101",21536 => "10010010",21537 => "01000000",21538 => "10001011",21539 => "00011111",21540 => "11001101",21541 => "10110001",21542 => "00001010",21543 => "11111010",21544 => "00011100",21545 => "11001001",21546 => "01110010",21547 => "10011000",21548 => "11100100",21549 => "01001000",21550 => "11111110",21551 => "10101110",21552 => "00010010",21553 => "10001010",21554 => "10100101",21555 => "11000010",21556 => "00011111",21557 => "00110101",21558 => "10011010",21559 => "00001110",21560 => "00111111",21561 => "01000000",21562 => "10011101",21563 => "00111000",21564 => "00101011",21565 => "01000000",21566 => "11100100",21567 => "01001010",21568 => "01110000",21569 => "11100010",21570 => "00100011",21571 => "11001110",21572 => "00011001",21573 => "00100001",21574 => "00111110",21575 => "11111001",21576 => "10010111",21577 => "01110110",21578 => "00011010",21579 => "00101111",21580 => "10010011",21581 => "00001000",21582 => "00110111",21583 => "10111000",21584 => "00111001",21585 => "11001010",21586 => "00001000",21587 => "10011010",21588 => "11111100",21589 => "01100100",21590 => "00101011",21591 => "01010100",21592 => "01001111",21593 => "11011111",21594 => "01010110",21595 => "11000100",21596 => "10101000",21597 => "10010111",21598 => "01100111",21599 => "00100111",21600 => "10000011",21601 => "01110100",21602 => "10001100",21603 => "10001100",21604 => "11101101",21605 => "01001110",21606 => "00010111",21607 => "00010111",21608 => "00001001",21609 => "00010000",21610 => "11001101",21611 => "11111010",21612 => "00110000",21613 => "01101100",21614 => "11000111",21615 => "10101100",21616 => "01000101",21617 => "11100110",21618 => "00101001",21619 => "01000010",21620 => "11001100",21621 => "10100100",21622 => "11111111",21623 => "11011011",21624 => "11010110",21625 => "00001010",21626 => "10110000",21627 => "10011011",21628 => "10101101",21629 => "00000100",21630 => "00100111",21631 => "10100010",21632 => "01000101",21633 => "10011001",21634 => "00110100",21635 => "01010010",21636 => "10001001",21637 => "00010001",21638 => "00111010",21639 => "01000111",21640 => "00011001",21641 => "00011000",21642 => "01001100",21643 => "00000110",21644 => "10001110",21645 => "11100001",21646 => "01011111",21647 => "11000001",21648 => "01110001",21649 => "11010111",21650 => "00100111",21651 => "01001011",21652 => "01100100",21653 => "10101000",21654 => "11100010",21655 => "00000111",21656 => "00010101",21657 => "11001000",21658 => "11011100",21659 => "01100100",21660 => "10011000",21661 => "10101110",21662 => "00110111",21663 => "10010110",21664 => "00001011",21665 => "10001011",21666 => "01001000",21667 => "10111100",21668 => "00110110",21669 => "10101100",21670 => "10100110",21671 => "01110110",21672 => "00010011",21673 => "01010001",21674 => "00011010",21675 => "00001000",21676 => "01010101",21677 => "00110110",21678 => "00100111",21679 => "01110100",21680 => "11111011",21681 => "10010100",21682 => "11000110",21683 => "11111111",21684 => "01011010",21685 => "00100101",21686 => "00001101",21687 => "10001001",21688 => "11001111",21689 => "10110000",21690 => "11111111",21691 => "11001010",21692 => "01110001",21693 => "01101000",21694 => "01110000",21695 => "01100000",21696 => "01011111",21697 => "00100010",21698 => "11010110",21699 => "11000011",21700 => "11101010",21701 => "10000011",21702 => "01000110",21703 => "01001010",21704 => "10111101",21705 => "00111011",21706 => "01001000",21707 => "01010110",21708 => "00100100",21709 => "10010111",21710 => "00001001",21711 => "11010101",21712 => "00111011",21713 => "00100011",21714 => "01111001",21715 => "01110011",21716 => "10101100",21717 => "01110010",21718 => "00101011",21719 => "00001111",21720 => "01011110",21721 => "11100010",21722 => "01011101",21723 => "01000110",21724 => "11000001",21725 => "11010011",21726 => "01011101",21727 => "00000110",21728 => "10011100",21729 => "10111000",21730 => "10111000",21731 => "11100100",21732 => "01100000",21733 => "10000101",21734 => "11110101",21735 => "00101111",21736 => "00011001",21737 => "00101100",21738 => "00100100",21739 => "00110100",21740 => "00111111",21741 => "01111101",21742 => "11010110",21743 => "10011101",21744 => "01010000",21745 => "10111000",21746 => "11111110",21747 => "11011011",21748 => "11101000",21749 => "11000001",21750 => "11000100",21751 => "00100111",21752 => "01110000",21753 => "01111111",21754 => "10100001",21755 => "00100110",21756 => "00100100",21757 => "11111100",21758 => "00101001",21759 => "10110001",21760 => "11011101",21761 => "01000001",21762 => "00011011",21763 => "00110011",21764 => "00000011",21765 => "01011010",21766 => "01110101",21767 => "00011110",21768 => "01111010",21769 => "00011011",21770 => "10101011",21771 => "00101101",21772 => "00011000",21773 => "11000010",21774 => "01101111",21775 => "10011010",21776 => "10111110",21777 => "00100101",21778 => "11000010",21779 => "11010101",21780 => "01110010",21781 => "00100000",21782 => "01110111",21783 => "00011000",21784 => "01001110",21785 => "01111011",21786 => "01010001",21787 => "01111001",21788 => "11111110",21789 => "11010000",21790 => "11111011",21791 => "00110010",21792 => "11000101",21793 => "11100100",21794 => "01100011",21795 => "01111011",21796 => "11011001",21797 => "00000110",21798 => "01001110",21799 => "00111011",21800 => "11001101",21801 => "11010011",21802 => "00110011",21803 => "01001011",21804 => "01010101",21805 => "11100011",21806 => "10101000",21807 => "11110110",21808 => "10000101",21809 => "11001111",21810 => "10101010",21811 => "11101000",21812 => "00100110",21813 => "00011110",21814 => "00011111",21815 => "01010011",21816 => "10110110",21817 => "10100011",21818 => "01011101",21819 => "01111110",21820 => "11010001",21821 => "11101110",21822 => "11100111",21823 => "11001000",21824 => "11001111",21825 => "10000111",21826 => "11011001",21827 => "00100010",21828 => "11011101",21829 => "01000111",21830 => "10100111",21831 => "00111101",21832 => "01110001",21833 => "00110111",21834 => "00111011",21835 => "10001001",21836 => "01000001",21837 => "00010010",21838 => "10110001",21839 => "00011100",21840 => "00000100",21841 => "10101110",21842 => "00001110",21843 => "10101111",21844 => "01110011",21845 => "11101110",21846 => "11101111",21847 => "00011010",21848 => "00010000",21849 => "10010111",21850 => "10100110",21851 => "00011111",21852 => "11101111",21853 => "00101000",21854 => "11011101",21855 => "01010101",21856 => "00111000",21857 => "11110011",21858 => "00100110",21859 => "10011111",21860 => "11001111",21861 => "01001110",21862 => "00001100",21863 => "10000010",21864 => "00100010",21865 => "11101110",21866 => "10000001",21867 => "11111011",21868 => "11000001",21869 => "11101001",21870 => "00101000",21871 => "00000111",21872 => "01011000",21873 => "00010010",21874 => "01111110",21875 => "00111001",21876 => "01111010",21877 => "10001010",21878 => "10001001",21879 => "00100000",21880 => "01000010",21881 => "11100111",21882 => "11111001",21883 => "01001111",21884 => "01010010",21885 => "10001011",21886 => "00001010",21887 => "00111101",21888 => "10101100",21889 => "11000100",21890 => "11101010",21891 => "10011011",21892 => "10100111",21893 => "00111101",21894 => "01110101",21895 => "00101111",21896 => "10010000",21897 => "00111111",21898 => "00101110",21899 => "11111111",21900 => "11000110",21901 => "11011101",21902 => "00100010",21903 => "01001111",21904 => "11000110",21905 => "00100110",21906 => "11100101",21907 => "11111100",21908 => "01000000",21909 => "11110101",21910 => "01011100",21911 => "10001110",21912 => "10110110",21913 => "11111100",21914 => "00001111",21915 => "11111001",21916 => "01111000",21917 => "11001110",21918 => "00100111",21919 => "00010000",21920 => "00001100",21921 => "00010011",21922 => "00100001",21923 => "01100111",21924 => "10011000",21925 => "00111010",21926 => "00000000",21927 => "10100011",21928 => "01110011",21929 => "01011111",21930 => "01100010",21931 => "00001100",21932 => "00000000",21933 => "00100110",21934 => "00000100",21935 => "11000111",21936 => "00111011",21937 => "01001100",21938 => "01111100",21939 => "00001001",21940 => "10100010",21941 => "00100000",21942 => "11101010",21943 => "11101110",21944 => "01110010",21945 => "11101101",21946 => "11110000",21947 => "10111001",21948 => "01011000",21949 => "11010101",21950 => "01010101",21951 => "11111011",21952 => "10100100",21953 => "01101010",21954 => "01111111",21955 => "11011011",21956 => "00000011",21957 => "11010111",21958 => "01110011",21959 => "01010011",21960 => "10010110",21961 => "01000001",21962 => "10111010",21963 => "10111000",21964 => "11001010",21965 => "01100010",21966 => "11000101",21967 => "01100001",21968 => "11101110",21969 => "00010110",21970 => "01110001",21971 => "01010110",21972 => "11011001",21973 => "00101110",21974 => "10111100",21975 => "10011100",21976 => "00100101",21977 => "01011000",21978 => "11001010",21979 => "10010110",21980 => "01000000",21981 => "01011000",21982 => "00011101",21983 => "00001101",21984 => "10010010",21985 => "10000001",21986 => "10000110",21987 => "01100101",21988 => "01011011",21989 => "11100001",21990 => "11011111",21991 => "11011101",21992 => "00001001",21993 => "10111010",21994 => "01011110",21995 => "10110100",21996 => "10101010",21997 => "00110110",21998 => "00001111",21999 => "00100001",22000 => "11011101",22001 => "11101000",22002 => "11000110",22003 => "01001100",22004 => "11011000",22005 => "01110101",22006 => "01010101",22007 => "00101101",22008 => "01010000",22009 => "11100110",22010 => "11101001",22011 => "00111000",22012 => "11000101",22013 => "11011101",22014 => "01000000",22015 => "10000011",22016 => "10001000",22017 => "00011101",22018 => "00001110",22019 => "00010000",22020 => "11111110",22021 => "11001111",22022 => "10101110",22023 => "00010110",22024 => "10110110",22025 => "10100111",22026 => "01000000",22027 => "00111111",22028 => "11110000",22029 => "11011100",22030 => "01111100",22031 => "01100100",22032 => "00101000",22033 => "00010001",22034 => "01000000",22035 => "11110000",22036 => "00101000",22037 => "10100101",22038 => "11011100",22039 => "11011000",22040 => "10111000",22041 => "11000100",22042 => "11010011",22043 => "01001110",22044 => "11011110",22045 => "11110010",22046 => "10110010",22047 => "01111010",22048 => "00000000",22049 => "11111111",22050 => "00100011",22051 => "00000111",22052 => "10110010",22053 => "01000011",22054 => "01001000",22055 => "00101010",22056 => "10110011",22057 => "00000000",22058 => "11100000",22059 => "11000100",22060 => "11000001",22061 => "11010000",22062 => "01111111",22063 => "00001110",22064 => "01100100",22065 => "01100011",22066 => "01100100",22067 => "01011011",22068 => "00100101",22069 => "01010010",22070 => "00000011",22071 => "01110101",22072 => "10110110",22073 => "11011101",22074 => "11111100",22075 => "10101000",22076 => "00111100",22077 => "10110010",22078 => "10011111",22079 => "00011011",22080 => "01110001",22081 => "01010001",22082 => "11011010",22083 => "00000011",22084 => "01110010",22085 => "01100111",22086 => "11100001",22087 => "10011010",22088 => "10101001",22089 => "01100110",22090 => "11001110",22091 => "00010001",22092 => "01010110",22093 => "01100001",22094 => "00100010",22095 => "00110010",22096 => "10111011",22097 => "11000001",22098 => "00111101",22099 => "10001001",22100 => "10100110",22101 => "10110111",22102 => "00010110",22103 => "11000101",22104 => "11001101",22105 => "11110111",22106 => "10010010",22107 => "10100000",22108 => "11111111",22109 => "11001010",22110 => "00001110",22111 => "01100000",22112 => "00111010",22113 => "00111101",22114 => "00001000",22115 => "10110101",22116 => "01100111",22117 => "01000001",22118 => "10101110",22119 => "10100001",22120 => "01011111",22121 => "01010101",22122 => "01011011",22123 => "00000101",22124 => "01000011",22125 => "00011010",22126 => "00111001",22127 => "01000011",22128 => "00101001",22129 => "01000010",22130 => "10100011",22131 => "00001001",22132 => "00011101",22133 => "01101101",22134 => "01100001",22135 => "11101100",22136 => "11011000",22137 => "00110011",22138 => "00110111",22139 => "00011000",22140 => "01000101",22141 => "01110100",22142 => "00101110",22143 => "10000010",22144 => "10101111",22145 => "11010011",22146 => "10110010",22147 => "00100000",22148 => "10010010",22149 => "01010001",22150 => "10110000",22151 => "10000010",22152 => "10100011",22153 => "11011100",22154 => "10010111",22155 => "01010101",22156 => "11001010",22157 => "11101101",22158 => "11000111",22159 => "00101100",22160 => "00010011",22161 => "10110111",22162 => "01010011",22163 => "10100111",22164 => "01101101",22165 => "01100110",22166 => "11000111",22167 => "01111101",22168 => "01001001",22169 => "10010000",22170 => "10101000",22171 => "11011100",22172 => "11011101",22173 => "11000000",22174 => "00111011",22175 => "10011000",22176 => "11010011",22177 => "00000110",22178 => "01010101",22179 => "10001010",22180 => "00111011",22181 => "00100000",22182 => "01010101",22183 => "00100111",22184 => "10101101",22185 => "10111100",22186 => "11011111",22187 => "11100011",22188 => "01001111",22189 => "01001110",22190 => "10100100",22191 => "10011101",22192 => "01010001",22193 => "00100100",22194 => "11110100",22195 => "10000011",22196 => "10101110",22197 => "10010100",22198 => "11101001",22199 => "11101010",22200 => "00011111",22201 => "00001111",22202 => "01110101",22203 => "10001101",22204 => "11101111",22205 => "01111010",22206 => "10001110",22207 => "01010100",22208 => "10100111",22209 => "11101111",22210 => "10011001",22211 => "00010001",22212 => "11010100",22213 => "00101010",22214 => "00000010",22215 => "00110000",22216 => "00011101",22217 => "00011011",22218 => "10111101",22219 => "01110100",22220 => "10110101",22221 => "10001000",22222 => "01000101",22223 => "10001011",22224 => "10100111",22225 => "10100011",22226 => "01011011",22227 => "00010100",22228 => "10001111",22229 => "11000010",22230 => "01001010",22231 => "01100100",22232 => "10001011",22233 => "11111010",22234 => "10010100",22235 => "10010100",22236 => "01111101",22237 => "00000011",22238 => "10100011",22239 => "10011111",22240 => "01100011",22241 => "00010011",22242 => "10000000",22243 => "00010010",22244 => "00000010",22245 => "00011001",22246 => "10011100",22247 => "11001010",22248 => "01110010",22249 => "01001100",22250 => "00000101",22251 => "01111101",22252 => "11101110",22253 => "01011010",22254 => "01000010",22255 => "11000001",22256 => "01100011",22257 => "01100011",22258 => "01100100",22259 => "10010001",22260 => "11101010",22261 => "01110011",22262 => "01011100",22263 => "00110101",22264 => "10101001",22265 => "11011101",22266 => "11111010",22267 => "11111001",22268 => "11000011",22269 => "11111101",22270 => "01101101",22271 => "00011111",22272 => "01100011",22273 => "10101111",22274 => "11111010",22275 => "10000110",22276 => "00010001",22277 => "00010111",22278 => "01111011",22279 => "01111010",22280 => "00110101",22281 => "00001001",22282 => "11001111",22283 => "11110100",22284 => "10011111",22285 => "01010111",22286 => "11010110",22287 => "00011010",22288 => "01100011",22289 => "00101110",22290 => "10100011",22291 => "10001101",22292 => "10110100",22293 => "00011101",22294 => "01100110",22295 => "10011101",22296 => "01110110",22297 => "01110010",22298 => "11001010",22299 => "00010101",22300 => "01110011",22301 => "00001110",22302 => "11011001",22303 => "00011100",22304 => "11000010",22305 => "01110001",22306 => "01011111",22307 => "00010010",22308 => "00000110",22309 => "01010010",22310 => "00101011",22311 => "11100001",22312 => "00001001",22313 => "11100011",22314 => "01100110",22315 => "00000011",22316 => "00111111",22317 => "00111001",22318 => "10100001",22319 => "11101100",22320 => "11100011",22321 => "11000011",22322 => "00000011",22323 => "00000110",22324 => "10000000",22325 => "01101011",22326 => "01010000",22327 => "11110010",22328 => "00001111",22329 => "10100111",22330 => "00111011",22331 => "11011010",22332 => "11111000",22333 => "10101110",22334 => "10110001",22335 => "01100111",22336 => "11101101",22337 => "01001101",22338 => "00011010",22339 => "10001110",22340 => "00000000",22341 => "00001010",22342 => "01110111",22343 => "01111011",22344 => "10001100",22345 => "01101001",22346 => "11100101",22347 => "11000010",22348 => "01111110",22349 => "00010001",22350 => "01010111",22351 => "10101110",22352 => "00000100",22353 => "00111010",22354 => "11101111",22355 => "11000010",22356 => "11110111",22357 => "01010111",22358 => "11101010",22359 => "11110001",22360 => "01000010",22361 => "01111000",22362 => "00100110",22363 => "11010001",22364 => "00000100",22365 => "11111010",22366 => "10110110",22367 => "01100111",22368 => "00100000",22369 => "01100110",22370 => "10101111",22371 => "11010110",22372 => "11111010",22373 => "10100100",22374 => "10111000",22375 => "00010011",22376 => "01101101",22377 => "01111101",22378 => "10000011",22379 => "11101001",22380 => "11000100",22381 => "00100000",22382 => "11010101",22383 => "10011110",22384 => "10011111",22385 => "01011011",22386 => "00111111",22387 => "10011010",22388 => "00000001",22389 => "00100111",22390 => "11010110",22391 => "11110100",22392 => "00001011",22393 => "01011010",22394 => "00010011",22395 => "11110110",22396 => "11000101",22397 => "01100010",22398 => "01011100",22399 => "00110001",22400 => "01011101",22401 => "01100011",22402 => "10010010",22403 => "11010001",22404 => "00001111",22405 => "10110100",22406 => "10110110",22407 => "00110001",22408 => "00100101",22409 => "10111001",22410 => "00001100",22411 => "00100110",22412 => "00110001",22413 => "01001011",22414 => "10101110",22415 => "10000111",22416 => "10101000",22417 => "11101011",22418 => "10101010",22419 => "01100010",22420 => "11000111",22421 => "10011010",22422 => "01010000",22423 => "00011101",22424 => "10100110",22425 => "11011010",22426 => "10011000",22427 => "00010010",22428 => "00011101",22429 => "01100010",22430 => "11101001",22431 => "11010101",22432 => "00111101",22433 => "11010010",22434 => "11000000",22435 => "00100100",22436 => "11101101",22437 => "11101011",22438 => "00010011",22439 => "10110000",22440 => "10000001",22441 => "00001001",22442 => "10100101",22443 => "00110100",22444 => "11001100",22445 => "10100000",22446 => "10010100",22447 => "11100010",22448 => "11110001",22449 => "01011101",22450 => "11001000",22451 => "11010000",22452 => "10111110",22453 => "01111101",22454 => "01100011",22455 => "01011100",22456 => "00101110",22457 => "01000110",22458 => "10100010",22459 => "00111010",22460 => "01011000",22461 => "10101100",22462 => "10101101",22463 => "10001110",22464 => "00100111",22465 => "01111110",22466 => "10101011",22467 => "01111010",22468 => "00110101",22469 => "10101111",22470 => "01111101",22471 => "10111011",22472 => "01110111",22473 => "11001011",22474 => "10101010",22475 => "11111001",22476 => "11011100",22477 => "00110101",22478 => "01111000",22479 => "11011011",22480 => "00001101",22481 => "10111101",22482 => "10100111",22483 => "10111100",22484 => "01001000",22485 => "11100100",22486 => "10111100",22487 => "01010110",22488 => "01000110",22489 => "10001000",22490 => "10000000",22491 => "01110000",22492 => "00110010",22493 => "11011111",22494 => "11001011",22495 => "01101111",22496 => "11000110",22497 => "10011000",22498 => "01010100",22499 => "00011000",22500 => "11000001",22501 => "11001110",22502 => "11111111",22503 => "10000101",22504 => "10100101",22505 => "00001111",22506 => "11001011",22507 => "10001010",22508 => "10110110",22509 => "01010100",22510 => "11001110",22511 => "11011101",22512 => "01010111",22513 => "00010011",22514 => "10001011",22515 => "10100101",22516 => "11001110",22517 => "11001110",22518 => "10111010",22519 => "11101010",22520 => "01111000",22521 => "11000011",22522 => "00001000",22523 => "10000111",22524 => "01101001",22525 => "01001001",22526 => "01100101",22527 => "11101011",22528 => "01101110",22529 => "11100110",22530 => "11010100",22531 => "00001001",22532 => "00100111",22533 => "11101001",22534 => "11011000",22535 => "11011110",22536 => "11001011",22537 => "10111010",22538 => "10111110",22539 => "11000110",22540 => "01111011",22541 => "01011011",22542 => "10110101",22543 => "11000110",22544 => "00010101",22545 => "01001101",22546 => "01011010",22547 => "10110001",22548 => "11011111",22549 => "01110011",22550 => "00110100",22551 => "01111000",22552 => "01000110",22553 => "01010100",22554 => "10010101",22555 => "01001110",22556 => "01100101",22557 => "00000001",22558 => "01101000",22559 => "10010011",22560 => "01001100",22561 => "01101111",22562 => "00100100",22563 => "00000101",22564 => "10111101",22565 => "00100111",22566 => "00000011",22567 => "00011101",22568 => "00101110",22569 => "01111010",22570 => "11110100",22571 => "11000001",22572 => "10100110",22573 => "11001110",22574 => "00100101",22575 => "00010001",22576 => "10110111",22577 => "11011010",22578 => "11100101",22579 => "11000101",22580 => "01010000",22581 => "11101011",22582 => "00010110",22583 => "00110101",22584 => "00011010",22585 => "11010100",22586 => "01010001",22587 => "01001010",22588 => "01000011",22589 => "10000111",22590 => "11000101",22591 => "00100010",22592 => "01110000",22593 => "11100010",22594 => "01010100",22595 => "11100010",22596 => "10001000",22597 => "01010011",22598 => "00100110",22599 => "11001101",22600 => "10011010",22601 => "01100101",22602 => "01111000",22603 => "11011011",22604 => "01111110",22605 => "01000010",22606 => "01111001",22607 => "00110010",22608 => "01101110",22609 => "10100100",22610 => "11111011",22611 => "00100011",22612 => "01010110",22613 => "11001001",22614 => "10100011",22615 => "00001111",22616 => "00100110",22617 => "10011100",22618 => "00000101",22619 => "11010110",22620 => "00110010",22621 => "10100110",22622 => "10011010",22623 => "10100001",22624 => "10011011",22625 => "10100001",22626 => "10011011",22627 => "00011111",22628 => "11110101",22629 => "10110101",22630 => "11101100",22631 => "01101010",22632 => "00111010",22633 => "10111000",22634 => "01010010",22635 => "00100001",22636 => "01110001",22637 => "10100011",22638 => "11101110",22639 => "11101111",22640 => "00000001",22641 => "10101010",22642 => "01110010",22643 => "10010000",22644 => "11010111",22645 => "01110101",22646 => "00101110",22647 => "11001000",22648 => "00001100",22649 => "01111000",22650 => "00100100",22651 => "11101111",22652 => "01111011",22653 => "11010110",22654 => "10000110",22655 => "00010011",22656 => "11010111",22657 => "00110001",22658 => "00001110",22659 => "11101010",22660 => "01000110",22661 => "10101011",22662 => "10101000",22663 => "00110100",22664 => "00110100",22665 => "10101111",22666 => "10000000",22667 => "00001010",22668 => "10101011",22669 => "01110100",22670 => "00111001",22671 => "10000011",22672 => "11100110",22673 => "00101001",22674 => "01001011",22675 => "10101011",22676 => "00011111",22677 => "10111100",22678 => "00110001",22679 => "00010001",22680 => "01001011",22681 => "01110111",22682 => "10000111",22683 => "01111000",22684 => "10101101",22685 => "01101010",22686 => "11000011",22687 => "10110010",22688 => "11100010",22689 => "11101010",22690 => "00000011",22691 => "11110111",22692 => "01010101",22693 => "10010100",22694 => "01101000",22695 => "00101001",22696 => "10111110",22697 => "11011011",22698 => "00100000",22699 => "00011100",22700 => "11110011",22701 => "11111110",22702 => "00110011",22703 => "10111000",22704 => "10010001",22705 => "11010001",22706 => "10000110",22707 => "00111100",22708 => "11001001",22709 => "01110100",22710 => "10101001",22711 => "10001110",22712 => "11111011",22713 => "00001010",22714 => "11111111",22715 => "01100111",22716 => "10110111",22717 => "11000011",22718 => "11010000",22719 => "01101100",22720 => "11001000",22721 => "01100111",22722 => "01001100",22723 => "01111111",22724 => "10100111",22725 => "00011011",22726 => "01011110",22727 => "01010001",22728 => "11110101",22729 => "01110010",22730 => "01000100",22731 => "11111110",22732 => "01011000",22733 => "00000110",22734 => "01100101",22735 => "11100101",22736 => "10111011",22737 => "10100100",22738 => "10001111",22739 => "01111111",22740 => "01010101",22741 => "01010100",22742 => "00011000",22743 => "10101010",22744 => "11110111",22745 => "10000011",22746 => "10100000",22747 => "11101010",22748 => "00001110",22749 => "00100000",22750 => "00101001",22751 => "10010011",22752 => "10000010",22753 => "00001001",22754 => "10001101",22755 => "10001000",22756 => "10111111",22757 => "10011010",22758 => "11011100",22759 => "00110001",22760 => "11000010",22761 => "01010110",22762 => "11011101",22763 => "10010001",22764 => "01000111",22765 => "11000000",22766 => "00101101",22767 => "10001000",22768 => "11001110",22769 => "01111000",22770 => "10000001",22771 => "10100000",22772 => "10101101",22773 => "00011111",22774 => "10101001",22775 => "10001011",22776 => "01101001",22777 => "00111101",22778 => "00111100",22779 => "10010110",22780 => "11100001",22781 => "11100100",22782 => "11001010",22783 => "00110010",22784 => "00110100",22785 => "01101000",22786 => "01111001",22787 => "00010110",22788 => "10010000",22789 => "11110001",22790 => "10010100",22791 => "10011110",22792 => "01010000",22793 => "00001011",22794 => "00100100",22795 => "01110100",22796 => "00100000",22797 => "11001100",22798 => "10110111",22799 => "00111100",22800 => "00101101",22801 => "10110011",22802 => "10011111",22803 => "11011110",22804 => "00111111",22805 => "00010111",22806 => "01111010",22807 => "01110000",22808 => "01111011",22809 => "10101101",22810 => "11101111",22811 => "00001010",22812 => "01110111",22813 => "11100101",22814 => "01010111",22815 => "10101110",22816 => "10101110",22817 => "11000111",22818 => "10100010",22819 => "00010110",22820 => "11010000",22821 => "00001011",22822 => "00011011",22823 => "10110000",22824 => "11110011",22825 => "11101001",22826 => "11010010",22827 => "11100101",22828 => "11010110",22829 => "11001111",22830 => "10101101",22831 => "10000001",22832 => "01101110",22833 => "11000110",22834 => "11111010",22835 => "10100101",22836 => "01001011",22837 => "01101011",22838 => "00000110",22839 => "11000011",22840 => "00001001",22841 => "00100101",22842 => "11001010",22843 => "10010101",22844 => "01001101",22845 => "01100100",22846 => "00011101",22847 => "01110001",22848 => "00001011",22849 => "01000000",22850 => "11000011",22851 => "10110011",22852 => "11100011",22853 => "00011111",22854 => "00000010",22855 => "11101000",22856 => "00010111",22857 => "11011100",22858 => "11110100",22859 => "01100111",22860 => "10100111",22861 => "00101100",22862 => "10001010",22863 => "11010010",22864 => "00011111",22865 => "10010110",22866 => "00111110",22867 => "01101100",22868 => "01010100",22869 => "11111000",22870 => "10111111",22871 => "01011011",22872 => "11100100",22873 => "10110101",22874 => "11101000",22875 => "10100111",22876 => "10011000",22877 => "01110100",22878 => "01101110",22879 => "11000100",22880 => "01110001",22881 => "00000011",22882 => "00101111",22883 => "10101010",22884 => "00111011",22885 => "01110010",22886 => "01010000",22887 => "11101000",22888 => "10110010",22889 => "01101111",22890 => "11110011",22891 => "00000000",22892 => "10111010",22893 => "01001111",22894 => "10110101",22895 => "10000001",22896 => "11011100",22897 => "00101011",22898 => "11110101",22899 => "11000111",22900 => "00010101",22901 => "11110101",22902 => "11010011",22903 => "00010000",22904 => "01010011",22905 => "01001101",22906 => "00100111",22907 => "01010101",22908 => "10100110",22909 => "11010101",22910 => "11100011",22911 => "11010000",22912 => "00111000",22913 => "00100000",22914 => "00111100",22915 => "10111111",22916 => "01010011",22917 => "10011111",22918 => "11010111",22919 => "00001011",22920 => "10001000",22921 => "11010001",22922 => "01100101",22923 => "01111111",22924 => "01100001",22925 => "11110111",22926 => "10101001",22927 => "00110111",22928 => "10101011",22929 => "10001001",22930 => "01101001",22931 => "11111000",22932 => "01011110",22933 => "01001111",22934 => "01000000",22935 => "11001111",22936 => "01100001",22937 => "11110111",22938 => "01110010",22939 => "10100110",22940 => "00101110",22941 => "11110111",22942 => "10001110",22943 => "10010000",22944 => "01001010",22945 => "10100001",22946 => "10110000",22947 => "01011110",22948 => "01101110",22949 => "01101101",22950 => "00010000",22951 => "01100110",22952 => "11110110",22953 => "00000100",22954 => "10011100",22955 => "01100111",22956 => "11001011",22957 => "00001110",22958 => "01011101",22959 => "10010100",22960 => "11011010",22961 => "11100011",22962 => "11001101",22963 => "01101110",22964 => "01001100",22965 => "11000011",22966 => "01000000",22967 => "01011110",22968 => "01001110",22969 => "11101110",22970 => "10001110",22971 => "10100011",22972 => "00100101",22973 => "10100010",22974 => "00101111",22975 => "11000110",22976 => "11010110",22977 => "01010110",22978 => "00100111",22979 => "11010000",22980 => "00111010",22981 => "01111001",22982 => "01111010",22983 => "10000000",22984 => "00111101",22985 => "10000001",22986 => "01001000",22987 => "11101010",22988 => "10010010",22989 => "10011101",22990 => "11100100",22991 => "10100011",22992 => "01010001",22993 => "00000001",22994 => "01100011",22995 => "10110010",22996 => "10011000",22997 => "10010011",22998 => "11011100",22999 => "01000101",23000 => "00100010",23001 => "00100101",23002 => "01101000",23003 => "01101110",23004 => "01010010",23005 => "01000110",23006 => "11010000",23007 => "01010000",23008 => "10100110",23009 => "10101011",23010 => "00110101",23011 => "10011000",23012 => "11010100",23013 => "11110110",23014 => "01010100",23015 => "01010100",23016 => "00101110",23017 => "00010010",23018 => "10010111",23019 => "00010000",23020 => "11000101",23021 => "10011110",23022 => "01110010",23023 => "01001010",23024 => "11101010",23025 => "00000001",23026 => "10111010",23027 => "00111110",23028 => "10101011",23029 => "01001110",23030 => "10100100",23031 => "00000010",23032 => "00001001",23033 => "01110011",23034 => "10011101",23035 => "01110000",23036 => "01111000",23037 => "01100101",23038 => "10001000",23039 => "10111101",23040 => "00110110",23041 => "10110001",23042 => "11000101",23043 => "01000101",23044 => "11101101",23045 => "00000101",23046 => "01101101",23047 => "10011111",23048 => "00000000",23049 => "11011100",23050 => "00111111",23051 => "11001101",23052 => "00110000",23053 => "10110101",23054 => "00010100",23055 => "10110011",23056 => "01101000",23057 => "01110010",23058 => "01001111",23059 => "11000111",23060 => "11100101",23061 => "00011001",23062 => "11010100",23063 => "01111010",23064 => "00010001",23065 => "00001110",23066 => "00000011",23067 => "00001100",23068 => "11100111",23069 => "00100111",23070 => "00110001",23071 => "01110101",23072 => "10001110",23073 => "10100010",23074 => "01110100",23075 => "01100110",23076 => "10011100",23077 => "01100011",23078 => "00101010",23079 => "01001001",23080 => "01011111",23081 => "10001011",23082 => "11110110",23083 => "10010100",23084 => "11010110",23085 => "00110111",23086 => "10101100",23087 => "10100010",23088 => "01000101",23089 => "11001001",23090 => "01010011",23091 => "00000000",23092 => "00110101",23093 => "10001111",23094 => "11101000",23095 => "10000010",23096 => "00010000",23097 => "11010100",23098 => "01010011",23099 => "11101100",23100 => "10100111",23101 => "10000100",23102 => "10010100",23103 => "11000101",23104 => "01111001",23105 => "01111010",23106 => "01000001",23107 => "00011011",23108 => "00110110",23109 => "01111111",23110 => "10010000",23111 => "01111110",23112 => "10100111",23113 => "10011100",23114 => "10101011",23115 => "00001101",23116 => "11000100",23117 => "01001111",23118 => "00010110",23119 => "11111111",23120 => "01100000",23121 => "11100010",23122 => "10011001",23123 => "01011001",23124 => "10011001",23125 => "10111100",23126 => "01011100",23127 => "00100001",23128 => "11100001",23129 => "11101111",23130 => "00100101",23131 => "10110101",23132 => "00001100",23133 => "11010101",23134 => "01110111",23135 => "10100111",23136 => "00101111",23137 => "10010001",23138 => "01110011",23139 => "11110100",23140 => "00101110",23141 => "10100001",23142 => "10010110",23143 => "00101111",23144 => "11000110",23145 => "01101101",23146 => "11100000",23147 => "11001110",23148 => "10110010",23149 => "01110000",23150 => "10001011",23151 => "01011110",23152 => "11001111",23153 => "10010000",23154 => "01111100",23155 => "11001000",23156 => "00111100",23157 => "01001101",23158 => "00010001",23159 => "10100001",23160 => "01110000",23161 => "01001000",23162 => "10101111",23163 => "01011110",23164 => "00010011",23165 => "10000111",23166 => "00011100",23167 => "00100000",23168 => "01010010",23169 => "01101101",23170 => "00011010",23171 => "00011100",23172 => "10101010",23173 => "11101001",23174 => "10100101",23175 => "11101110",23176 => "01101000",23177 => "11010011",23178 => "10111001",23179 => "10001001",23180 => "00001111",23181 => "11101110",23182 => "10001101",23183 => "00111011",23184 => "01101000",23185 => "01010000",23186 => "10000010",23187 => "00011100",23188 => "10111111",23189 => "01001100",23190 => "00100000",23191 => "10001010",23192 => "00101101",23193 => "00100000",23194 => "01101010",23195 => "00000000",23196 => "01000110",23197 => "10001001",23198 => "01010100",23199 => "00010110",23200 => "00011001",23201 => "00010111",23202 => "10011001",23203 => "11101000",23204 => "11111001",23205 => "10011010",23206 => "00100110",23207 => "11000100",23208 => "00000110",23209 => "10111000",23210 => "01000110",23211 => "00101010",23212 => "11100111",23213 => "11100001",23214 => "11111110",23215 => "10010100",23216 => "11010110",23217 => "01101010",23218 => "11111111",23219 => "01000011",23220 => "01011100",23221 => "10100101",23222 => "00110011",23223 => "00000010",23224 => "11100011",23225 => "11111000",23226 => "11010001",23227 => "01110010",23228 => "10101110",23229 => "11010010",23230 => "00001000",23231 => "01000110",23232 => "00110001",23233 => "11011010",23234 => "00100000",23235 => "01100101",23236 => "11011001",23237 => "10011101",23238 => "10001110",23239 => "10001010",23240 => "11101110",23241 => "01000110",23242 => "11011101",23243 => "10001110",23244 => "01110100",23245 => "01100110",23246 => "11011101",23247 => "10011100",23248 => "10001111",23249 => "11001111",23250 => "01110100",23251 => "10000000",23252 => "11011001",23253 => "01111001",23254 => "00010000",23255 => "01101110",23256 => "11101100",23257 => "00111110",23258 => "00100010",23259 => "11011100",23260 => "00001011",23261 => "11100000",23262 => "10010010",23263 => "01000000",23264 => "00000111",23265 => "10000110",23266 => "10011000",23267 => "01101010",23268 => "10111000",23269 => "11111111",23270 => "11100010",23271 => "11110110",23272 => "10100010",23273 => "11010010",23274 => "11101110",23275 => "10011000",23276 => "00110011",23277 => "01010101",23278 => "01100011",23279 => "10101011",23280 => "11111100",23281 => "01101101",23282 => "01011110",23283 => "00001011",23284 => "10000100",23285 => "01010001",23286 => "01101110",23287 => "11101101",23288 => "01010110",23289 => "01101010",23290 => "01111010",23291 => "11101101",23292 => "11111010",23293 => "10110010",23294 => "11001111",23295 => "01101011",23296 => "11101001",23297 => "11011110",23298 => "11100001",23299 => "11010000",23300 => "01010001",23301 => "00111101",23302 => "10011000",23303 => "01110010",23304 => "11001001",23305 => "10001111",23306 => "11000010",23307 => "11101000",23308 => "01001111",23309 => "11000110",23310 => "10101000",23311 => "10000100",23312 => "10111110",23313 => "11001000",23314 => "00001001",23315 => "01001001",23316 => "01001011",23317 => "00011111",23318 => "10111011",23319 => "01101110",23320 => "11101111",23321 => "10000111",23322 => "11101010",23323 => "00011000",23324 => "01000100",23325 => "01101111",23326 => "00000100",23327 => "11010100",23328 => "00000001",23329 => "01111011",23330 => "10011100",23331 => "00101111",23332 => "10111110",23333 => "01011111",23334 => "00010100",23335 => "11110110",23336 => "11011111",23337 => "01000111",23338 => "11100111",23339 => "01111001",23340 => "10101100",23341 => "10010110",23342 => "10100110",23343 => "01000100",23344 => "00110101",23345 => "00110000",23346 => "00110111",23347 => "00010101",23348 => "11001101",23349 => "00101000",23350 => "11010011",23351 => "10111000",23352 => "11000010",23353 => "10001100",23354 => "10100010",23355 => "01110001",23356 => "01011111",23357 => "01110010",23358 => "01100100",23359 => "11001010",23360 => "01011010",23361 => "01010110",23362 => "00011001",23363 => "10001011",23364 => "11000010",23365 => "11111010",23366 => "10010010",23367 => "10000000",23368 => "01100100",23369 => "11001010",23370 => "10011011",23371 => "11010100",23372 => "00011100",23373 => "11111111",23374 => "01011111",23375 => "11110011",23376 => "11011011",23377 => "01010001",23378 => "10111110",23379 => "00000000",23380 => "00011101",23381 => "00001100",23382 => "10001011",23383 => "10100101",23384 => "10110110",23385 => "11110011",23386 => "11101000",23387 => "11110000",23388 => "11111011",23389 => "01001111",23390 => "10100100",23391 => "00100000",23392 => "01100000",23393 => "01101000",23394 => "01010100",23395 => "11101010",23396 => "10101010",23397 => "10100011",23398 => "10011110",23399 => "01000101",23400 => "00100101",23401 => "00000011",23402 => "01011001",23403 => "01101100",23404 => "10000000",23405 => "11100001",23406 => "01010010",23407 => "01111111",23408 => "11101101",23409 => "11011111",23410 => "00110100",23411 => "11001111",23412 => "01110001",23413 => "01000100",23414 => "01011101",23415 => "11101001",23416 => "01011010",23417 => "10101110",23418 => "11001101",23419 => "10000110",23420 => "00011001",23421 => "00001000",23422 => "11100100",23423 => "01100101",23424 => "01011010",23425 => "10010111",23426 => "01111010",23427 => "01111100",23428 => "00011001",23429 => "10001011",23430 => "10010010",23431 => "01110111",23432 => "11110101",23433 => "11100110",23434 => "00111001",23435 => "11010111",23436 => "01111011",23437 => "11001110",23438 => "01110100",23439 => "11110010",23440 => "10010010",23441 => "11110110",23442 => "10111011",23443 => "01011000",23444 => "00000001",23445 => "10110000",23446 => "11111011",23447 => "00010111",23448 => "00000011",23449 => "11110000",23450 => "00001110",23451 => "11001101",23452 => "11000100",23453 => "00010101",23454 => "11100101",23455 => "10101001",23456 => "11111110",23457 => "10101111",23458 => "01011011",23459 => "00111000",23460 => "00010000",23461 => "11001011",23462 => "00110110",23463 => "11100010",23464 => "01100101",23465 => "10111011",23466 => "11011101",23467 => "01101101",23468 => "10111101",23469 => "00101101",23470 => "11001010",23471 => "00101101",23472 => "00100011",23473 => "00011110",23474 => "10111100",23475 => "11000100",23476 => "01011100",23477 => "11000100",23478 => "01001110",23479 => "11010011",23480 => "01110011",23481 => "00000110",23482 => "00001011",23483 => "10100011",23484 => "11000001",23485 => "11110110",23486 => "01011011",23487 => "01100010",23488 => "10000000",23489 => "01101101",23490 => "00111101",23491 => "10000010",23492 => "00101010",23493 => "10110010",23494 => "11001001",23495 => "10011010",23496 => "11111011",23497 => "00110001",23498 => "10111001",23499 => "10110101",23500 => "10101001",23501 => "00000100",23502 => "10100110",23503 => "01000010",23504 => "11110000",23505 => "11000100",23506 => "10010111",23507 => "01001100",23508 => "10000100",23509 => "01111010",23510 => "10100001",23511 => "11010010",23512 => "01100100",23513 => "10111100",23514 => "10011010",23515 => "00001010",23516 => "11011011",23517 => "00010101",23518 => "11001110",23519 => "11100001",23520 => "10010011",23521 => "10110010",23522 => "10000011",23523 => "00100001",23524 => "00110001",23525 => "11010101",23526 => "01010111",23527 => "10111101",23528 => "01001010",23529 => "10110010",23530 => "11001011",23531 => "01011000",23532 => "01000110",23533 => "10001100",23534 => "01001000",23535 => "10011011",23536 => "00000010",23537 => "11101111",23538 => "00111111",23539 => "10001010",23540 => "01100100",23541 => "00010011",23542 => "01111111",23543 => "01000000",23544 => "01100001",23545 => "01101110",23546 => "11000100",23547 => "11011101",23548 => "11011010",23549 => "01001001",23550 => "11110101",23551 => "11100101",23552 => "01001111",23553 => "10111111",23554 => "10001001",23555 => "00010101",23556 => "10011000",23557 => "11010011",23558 => "10111001",23559 => "01000110",23560 => "01010100",23561 => "11010000",23562 => "00100010",23563 => "11101000",23564 => "01110010",23565 => "11011100",23566 => "01001010",23567 => "01110001",23568 => "11001110",23569 => "10110000",23570 => "00101001",23571 => "01110100",23572 => "00001001",23573 => "11000000",23574 => "10010001",23575 => "00101101",23576 => "11101111",23577 => "10010000",23578 => "00101111",23579 => "00110001",23580 => "01011101",23581 => "00111011",23582 => "11110000",23583 => "01011000",23584 => "10001110",23585 => "01011000",23586 => "01110011",23587 => "01100000",23588 => "11110101",23589 => "01010111",23590 => "00111010",23591 => "11001011",23592 => "11001100",23593 => "10111101",23594 => "01001100",23595 => "01011010",23596 => "01111110",23597 => "01100011",23598 => "11110000",23599 => "11101010",23600 => "10110010",23601 => "00101000",23602 => "01111100",23603 => "01011000",23604 => "00011111",23605 => "01101000",23606 => "11010101",23607 => "10000101",23608 => "10101110",23609 => "01111110",23610 => "10110001",23611 => "00010100",23612 => "11100111",23613 => "00011111",23614 => "10001011",23615 => "11010101",23616 => "00000111",23617 => "00000011",23618 => "10100111",23619 => "11111111",23620 => "01111010",23621 => "10010100",23622 => "11000111",23623 => "10100100",23624 => "10110100",23625 => "11110110",23626 => "10110000",23627 => "10001101",23628 => "00101010",23629 => "10000011",23630 => "10011001",23631 => "01110011",23632 => "01001110",23633 => "10001000",23634 => "10011011",23635 => "00010011",23636 => "00011101",23637 => "01110000",23638 => "11100110",23639 => "11010111",23640 => "00110000",23641 => "11001111",23642 => "00101100",23643 => "00000011",23644 => "00011011",23645 => "11110011",23646 => "11100001",23647 => "01010100",23648 => "10100011",23649 => "01010000",23650 => "11101010",23651 => "01010100",23652 => "11100011",23653 => "01100001",23654 => "11111101",23655 => "11100010",23656 => "11000000",23657 => "01101101",23658 => "11011000",23659 => "00110110",23660 => "01010000",23661 => "01110101",23662 => "01000001",23663 => "01111100",23664 => "10100101",23665 => "01010000",23666 => "11111001",23667 => "11000010",23668 => "10110000",23669 => "10000010",23670 => "01010010",23671 => "11101011",23672 => "01001100",23673 => "11101010",23674 => "00010011",23675 => "11010011",23676 => "11100001",23677 => "01100110",23678 => "10100011",23679 => "01000100",23680 => "10100100",23681 => "11010110",23682 => "01111000",23683 => "00110010",23684 => "00001101",23685 => "11101000",23686 => "11111010",23687 => "00101100",23688 => "11110010",23689 => "01000100",23690 => "01100110",23691 => "10010101",23692 => "10001100",23693 => "00111011",23694 => "01111111",23695 => "11000101",23696 => "01100100",23697 => "01000110",23698 => "01101001",23699 => "11101100",23700 => "11011001",23701 => "01111100",23702 => "10110000",23703 => "11000001",23704 => "01011110",23705 => "01010100",23706 => "10101010",23707 => "01010011",23708 => "10111111",23709 => "11111110",23710 => "01001101",23711 => "00000010",23712 => "10010101",23713 => "10101101",23714 => "01010000",23715 => "01110001",23716 => "10010000",23717 => "00111100",23718 => "11000111",23719 => "01001111",23720 => "11000101",23721 => "11111110",23722 => "11010001",23723 => "10000100",23724 => "11000000",23725 => "01010011",23726 => "10011011",23727 => "00110011",23728 => "00010101",23729 => "11111001",23730 => "00010100",23731 => "10101110",23732 => "01111101",23733 => "00011111",23734 => "00011001",23735 => "01100100",23736 => "01110001",23737 => "10011100",23738 => "00100101",23739 => "11100101",23740 => "00100110",23741 => "11101011",23742 => "00110011",23743 => "01001100",23744 => "10111100",23745 => "01000111",23746 => "10010010",23747 => "11101111",23748 => "00010110",23749 => "00110010",23750 => "01111100",23751 => "11010010",23752 => "11010011",23753 => "01000101",23754 => "10011100",23755 => "11000010",23756 => "10111101",23757 => "11100001",23758 => "10101001",23759 => "01101111",23760 => "01100110",23761 => "00110100",23762 => "11100010",23763 => "11101101",23764 => "10010001",23765 => "10100100",23766 => "11100100",23767 => "00001111",23768 => "10111100",23769 => "00000100",23770 => "01110110",23771 => "01001010",23772 => "11100010",23773 => "00010010",23774 => "01001011",23775 => "01101110",23776 => "00010100",23777 => "00100010",23778 => "01110000",23779 => "10110111",23780 => "01101010",23781 => "01111111",23782 => "00011111",23783 => "01011110",23784 => "01100110",23785 => "11000110",23786 => "11101111",23787 => "10000101",23788 => "10100011",23789 => "00110000",23790 => "10111010",23791 => "00101010",23792 => "00000000",23793 => "10010110",23794 => "11000000",23795 => "11111100",23796 => "01000111",23797 => "11000011",23798 => "11001010",23799 => "11101010",23800 => "01100100",23801 => "01011110",23802 => "10001001",23803 => "10110100",23804 => "10010001",23805 => "11001111",23806 => "01101110",23807 => "10101100",23808 => "10100110",23809 => "11100010",23810 => "01110000",23811 => "00111100",23812 => "11101011",23813 => "00100000",23814 => "11100100",23815 => "01000010",23816 => "00010101",23817 => "00110010",23818 => "10001110",23819 => "10011001",23820 => "01100001",23821 => "11110100",23822 => "11111100",23823 => "11011100",23824 => "10000010",23825 => "01111110",23826 => "11100010",23827 => "11110000",23828 => "01101101",23829 => "01010100",23830 => "11001011",23831 => "10010000",23832 => "00000000",23833 => "11000101",23834 => "01101011",23835 => "00100101",23836 => "11001011",23837 => "01010111",23838 => "10111001",23839 => "10000110",23840 => "11111101",23841 => "10110010",23842 => "10111011",23843 => "10110110",23844 => "00010100",23845 => "00110011",23846 => "01111111",23847 => "00010101",23848 => "11100111",23849 => "10111000",23850 => "11010000",23851 => "10000010",23852 => "10101001",23853 => "11110001",23854 => "01100011",23855 => "01100100",23856 => "00100001",23857 => "10111010",23858 => "01111100",23859 => "01010011",23860 => "01011101",23861 => "11011010",23862 => "00111000",23863 => "01011010",23864 => "10000000",23865 => "01110110",23866 => "01011110",23867 => "00011110",23868 => "11001010",23869 => "10100111",23870 => "11100001",23871 => "10110010",23872 => "01000010",23873 => "00110011",23874 => "00110001",23875 => "01001010",23876 => "10110100",23877 => "11101111",23878 => "11111111",23879 => "01010101",23880 => "10111001",23881 => "00000010",23882 => "01100011",23883 => "00011010",23884 => "01011101",23885 => "10010110",23886 => "10111001",23887 => "01010110",23888 => "11101111",23889 => "11001011",23890 => "10101010",23891 => "01101110",23892 => "00111010",23893 => "00100111",23894 => "01011001",23895 => "00100000",23896 => "00011011",23897 => "00110000",23898 => "01100101",23899 => "01001101",23900 => "10111000",23901 => "00101001",23902 => "11111010",23903 => "01110001",23904 => "10011101",23905 => "00110110",23906 => "11101011",23907 => "11011101",23908 => "10011000",23909 => "01010010",23910 => "11000011",23911 => "01001001",23912 => "01010100",23913 => "11010111",23914 => "10001000",23915 => "11110010",23916 => "01111110",23917 => "10010000",23918 => "01101001",23919 => "01011010",23920 => "11000001",23921 => "11011001",23922 => "11101101",23923 => "00011101",23924 => "01101111",23925 => "11100011",23926 => "10110110",23927 => "11001111",23928 => "11111101",23929 => "00101110",23930 => "11110010",23931 => "00100011",23932 => "01100111",23933 => "00001001",23934 => "11111101",23935 => "01010101",23936 => "11101011",23937 => "10101110",23938 => "01011100",23939 => "00001011",23940 => "00111011",23941 => "10001000",23942 => "01111000",23943 => "00101111",23944 => "11010011",23945 => "11110010",23946 => "10011010",23947 => "11011001",23948 => "10010010",23949 => "11010001",23950 => "01011000",23951 => "11011111",23952 => "01000000",23953 => "01101111",23954 => "00110100",23955 => "01000111",23956 => "11001110",23957 => "01110100",23958 => "10001110",23959 => "11101001",23960 => "11111100",23961 => "01110000",23962 => "10111110",23963 => "00011010",23964 => "10101010",23965 => "01001000",23966 => "10101010",23967 => "00000111",23968 => "01000100",23969 => "11001011",23970 => "00001000",23971 => "10011100",23972 => "11111001",23973 => "11011101",23974 => "00101100",23975 => "11101000",23976 => "10101011",23977 => "10111010",23978 => "01101101",23979 => "00001001",23980 => "00011010",23981 => "01111011",23982 => "01110101",23983 => "11101101",23984 => "11110001",23985 => "11110000",23986 => "00110101",23987 => "10111101",23988 => "10101101",23989 => "11100110",23990 => "00011001",23991 => "01111110",23992 => "00010110",23993 => "10001001",23994 => "11011100",23995 => "00111000",23996 => "00001001",23997 => "01100110",23998 => "00101101",23999 => "11110110",24000 => "11001110",24001 => "01111001",24002 => "10001101",24003 => "00001101",24004 => "01110110",24005 => "00101010",24006 => "01110000",24007 => "11100011",24008 => "00111101",24009 => "11001010",24010 => "00110100",24011 => "10000110",24012 => "00000001",24013 => "01111011",24014 => "11000011",24015 => "10010000",24016 => "01100001",24017 => "00001011",24018 => "01101010",24019 => "11101010",24020 => "01100110",24021 => "10010101",24022 => "10100111",24023 => "00001011",24024 => "00100111",24025 => "00011010",24026 => "00101100",24027 => "10000110",24028 => "11010001",24029 => "11101011",24030 => "01010100",24031 => "00011000",24032 => "10010101",24033 => "00101110",24034 => "10001001",24035 => "01000010",24036 => "00010100",24037 => "00000011",24038 => "11010001",24039 => "01100010",24040 => "00100101",24041 => "11100110",24042 => "00000010",24043 => "01000110",24044 => "11011101",24045 => "11010011",24046 => "01010110",24047 => "01111111",24048 => "01100111",24049 => "11110101",24050 => "10101011",24051 => "11100100",24052 => "01010010",24053 => "00000001",24054 => "00101101",24055 => "10110111",24056 => "01110111",24057 => "11000100",24058 => "00111100",24059 => "01001111",24060 => "00101011",24061 => "11111010",24062 => "00001101",24063 => "01001000",24064 => "10001100",24065 => "00110100",24066 => "00000110",24067 => "10100101",24068 => "10111100",24069 => "11100000",24070 => "11111111",24071 => "00100111",24072 => "00110101",24073 => "11101001",24074 => "00010101",24075 => "11010010",24076 => "11100011",24077 => "10101100",24078 => "01000000",24079 => "01111101",24080 => "10101111",24081 => "11110001",24082 => "01111111",24083 => "01100011",24084 => "11110100",24085 => "11000101",24086 => "11011101",24087 => "10111010",24088 => "00010101",24089 => "11000010",24090 => "00100000",24091 => "00100111",24092 => "01101110",24093 => "00011000",24094 => "10000111",24095 => "01001001",24096 => "11110011",24097 => "00100011",24098 => "11001000",24099 => "10000100",24100 => "01011101",24101 => "00110101",24102 => "00101101",24103 => "00010111",24104 => "00111001",24105 => "00111001",24106 => "10101100",24107 => "00111001",24108 => "11011000",24109 => "11001110",24110 => "11111000",24111 => "10010111",24112 => "10110000",24113 => "11010111",24114 => "01001011",24115 => "00011100",24116 => "11000111",24117 => "10100100",24118 => "00110011",24119 => "01010001",24120 => "10111000",24121 => "01100110",24122 => "01110001",24123 => "11010110",24124 => "01110000",24125 => "11010010",24126 => "11111111",24127 => "10010001",24128 => "11101110",24129 => "10101001",24130 => "11000100",24131 => "11101101",24132 => "11100001",24133 => "00100111",24134 => "01001010",24135 => "10000111",24136 => "01001011",24137 => "11110111",24138 => "11110111",24139 => "11001001",24140 => "10111110",24141 => "10000101",24142 => "11001111",24143 => "10110010",24144 => "11100100",24145 => "00010000",24146 => "00100100",24147 => "11111010",24148 => "11000010",24149 => "10000011",24150 => "10111110",24151 => "10100101",24152 => "10010001",24153 => "00101101",24154 => "10011011",24155 => "00011011",24156 => "00011101",24157 => "01110000",24158 => "00110011",24159 => "11100010",24160 => "11000101",24161 => "11111011",24162 => "00000100",24163 => "11011010",24164 => "00110110",24165 => "00010001",24166 => "11111100",24167 => "00100001",24168 => "10001001",24169 => "10100101",24170 => "00001100",24171 => "00001010",24172 => "10111101",24173 => "11101111",24174 => "00010011",24175 => "00010101",24176 => "00001010",24177 => "11111001",24178 => "10101001",24179 => "11101011",24180 => "11000010",24181 => "10011110",24182 => "10000111",24183 => "10100000",24184 => "10110001",24185 => "10010000",24186 => "00101101",24187 => "11100001",24188 => "11100101",24189 => "10010111",24190 => "10011111",24191 => "00001110",24192 => "10010101",24193 => "11101000",24194 => "01011000",24195 => "10110010",24196 => "10100110",24197 => "10000110",24198 => "11100001",24199 => "11100110",24200 => "01110111",24201 => "01010010",24202 => "00001011",24203 => "00000011",24204 => "11011110",24205 => "01000101",24206 => "11100101",24207 => "00010010",24208 => "11000011",24209 => "10111010",24210 => "11010100",24211 => "11101011",24212 => "11100011",24213 => "00011011",24214 => "00000100",24215 => "01000110",24216 => "11100111",24217 => "11110011",24218 => "00100111",24219 => "00011011",24220 => "11001101",24221 => "01101000",24222 => "11100101",24223 => "00000001",24224 => "01001001",24225 => "11111000",24226 => "00111110",24227 => "11101011",24228 => "11011010",24229 => "00111101",24230 => "00001100",24231 => "01111011",24232 => "00000000",24233 => "00110111",24234 => "01100101",24235 => "11101011",24236 => "11001010",24237 => "01010101",24238 => "00000011",24239 => "10111111",24240 => "10101010",24241 => "00011011",24242 => "01001010",24243 => "11001000",24244 => "11101011",24245 => "01011111",24246 => "01111000",24247 => "01010011",24248 => "00010110",24249 => "00110101",24250 => "10011101",24251 => "11000110",24252 => "10000010",24253 => "01001000",24254 => "00000111",24255 => "01100100",24256 => "00110101",24257 => "11011100",24258 => "10101010",24259 => "10110110",24260 => "10000111",24261 => "10001101",24262 => "00001011",24263 => "01011001",24264 => "00100110",24265 => "10001010",24266 => "11100101",24267 => "11110001",24268 => "10101010",24269 => "10011010",24270 => "01000101",24271 => "10000010",24272 => "00010011",24273 => "11110100",24274 => "00010101",24275 => "11100111",24276 => "11011111",24277 => "00101111",24278 => "00010110",24279 => "01110101",24280 => "10000010",24281 => "01001011",24282 => "00010001",24283 => "10101011",24284 => "01101101",24285 => "00100111",24286 => "00110011",24287 => "11100000",24288 => "01000100",24289 => "01001100",24290 => "11111111",24291 => "01110111",24292 => "10100101",24293 => "01000001",24294 => "01100011",24295 => "11011011",24296 => "01110010",24297 => "10011001",24298 => "00110011",24299 => "01110001",24300 => "00111011",24301 => "00011111",24302 => "11011001",24303 => "00111010",24304 => "00111101",24305 => "10101001",24306 => "00001000",24307 => "01001010",24308 => "10110010",24309 => "00001101",24310 => "00111111",24311 => "11000011",24312 => "11010100",24313 => "01101010",24314 => "11000111",24315 => "11000010",24316 => "11001110",24317 => "00000000",24318 => "01010101",24319 => "10001011",24320 => "10010111",24321 => "11000010",24322 => "00100111",24323 => "11101000",24324 => "01111101",24325 => "00000110",24326 => "11100111",24327 => "10000010",24328 => "01000011",24329 => "01000010",24330 => "11000001",24331 => "10110000",24332 => "10110110",24333 => "00111001",24334 => "10101010",24335 => "01111100",24336 => "10100011",24337 => "01011000",24338 => "10110010",24339 => "01010100",24340 => "00010100",24341 => "11100100",24342 => "00010100",24343 => "01100100",24344 => "00010110",24345 => "01111001",24346 => "01011000",24347 => "01011011",24348 => "01010101",24349 => "11010110",24350 => "11110000",24351 => "01110101",24352 => "10101001",24353 => "01111101",24354 => "01101001",24355 => "01101000",24356 => "00010101",24357 => "11100000",24358 => "01010011",24359 => "11111110",24360 => "01000111",24361 => "11110011",24362 => "00111110",24363 => "10101011",24364 => "10111110",24365 => "10101100",24366 => "01000100",24367 => "00011000",24368 => "11110010",24369 => "00011101",24370 => "01001101",24371 => "10110100",24372 => "01011101",24373 => "01101000",24374 => "11000010",24375 => "10101100",24376 => "01110100",24377 => "00001001",24378 => "10101001",24379 => "11101001",24380 => "01101100",24381 => "11111100",24382 => "10101000",24383 => "01001101",24384 => "01011011",24385 => "00100011",24386 => "11100011",24387 => "01110111",24388 => "10110100",24389 => "01101100",24390 => "00011000",24391 => "11100111",24392 => "10111011",24393 => "11001101",24394 => "01101101",24395 => "01001001",24396 => "11010101",24397 => "10011001",24398 => "01111011",24399 => "00010001",24400 => "10100001",24401 => "00001110",24402 => "10111100",24403 => "10101110",24404 => "11101111",24405 => "11101000",24406 => "00111110",24407 => "10011110",24408 => "01010110",24409 => "10010110",24410 => "00101011",24411 => "11001101",24412 => "10010000",24413 => "01110001",24414 => "01010111",24415 => "01010001",24416 => "11111000",24417 => "01100010",24418 => "01111010",24419 => "10111000",24420 => "10101010",24421 => "01111000",24422 => "01110110",24423 => "10100101",24424 => "11101111",24425 => "00100101",24426 => "01000010",24427 => "01011100",24428 => "01110001",24429 => "00000000",24430 => "00101010",24431 => "01101101",24432 => "11111100",24433 => "10010101",24434 => "10010011",24435 => "01001001",24436 => "11010110",24437 => "11001000",24438 => "10111111",24439 => "01110100",24440 => "01100100",24441 => "00000001",24442 => "00111101",24443 => "11110010",24444 => "10101010",24445 => "10011101",24446 => "10001000",24447 => "01011100",24448 => "00111111",24449 => "01011000",24450 => "00111110",24451 => "01100101",24452 => "00001010",24453 => "01100100",24454 => "00001001",24455 => "11010000",24456 => "10111100",24457 => "00110111",24458 => "01111100",24459 => "01010101",24460 => "10111111",24461 => "00111100",24462 => "00100001",24463 => "11100101",24464 => "01010001",24465 => "11001010",24466 => "00011111",24467 => "10111011",24468 => "00011111",24469 => "01000111",24470 => "11000000",24471 => "10000111",24472 => "11100011",24473 => "10110001",24474 => "01010001",24475 => "01001000",24476 => "11110100",24477 => "01110011",24478 => "10011101",24479 => "11011011",24480 => "00100100",24481 => "11110000",24482 => "10001011",24483 => "11000011",24484 => "11000100",24485 => "00001100",24486 => "00001000",24487 => "00111101",24488 => "00001000",24489 => "10110001",24490 => "11100100",24491 => "00000001",24492 => "11011001",24493 => "10011011",24494 => "10110001",24495 => "01000011",24496 => "01110000",24497 => "01101100",24498 => "10110110",24499 => "01011101",24500 => "11100000",24501 => "01001000",24502 => "11100011",24503 => "11110101",24504 => "10110110",24505 => "00100010",24506 => "11110111",24507 => "10001001",24508 => "11101110",24509 => "00001101",24510 => "10001111",24511 => "01000111",24512 => "00001101",24513 => "11011001",24514 => "10101001",24515 => "11101111",24516 => "11110000",24517 => "00101000",24518 => "00000111",24519 => "10111100",24520 => "00100001",24521 => "00100011",24522 => "01001110",24523 => "11000101",24524 => "01001010",24525 => "11110000",24526 => "01110011",24527 => "10111111",24528 => "00100010",24529 => "00000110",24530 => "10010000",24531 => "11000011",24532 => "10101000",24533 => "11110100",24534 => "00001100",24535 => "01000111",24536 => "11000011",24537 => "00100111",24538 => "01111110",24539 => "10111100",24540 => "11000001",24541 => "10110101",24542 => "10001000",24543 => "11100010",24544 => "00110010",24545 => "01000000",24546 => "11100001",24547 => "11101011",24548 => "10000110",24549 => "10111001",24550 => "11111000",24551 => "01110100",24552 => "01110110",24553 => "11111111",24554 => "01001011",24555 => "11010000",24556 => "00100010",24557 => "00101010",24558 => "11110101",24559 => "10100101",24560 => "11011000",24561 => "01001101",24562 => "00000010",24563 => "00000011",24564 => "00000001",24565 => "01100011",24566 => "10111111",24567 => "01111001",24568 => "11111111",24569 => "10000000",24570 => "01011100",24571 => "10001110",24572 => "00100111",24573 => "00101111",24574 => "11111001",24575 => "01010100",24576 => "01111001",24577 => "11010100",24578 => "00110111",24579 => "00110100",24580 => "10000101",24581 => "10000110",24582 => "00011001",24583 => "01010001",24584 => "01110110",24585 => "10111011",24586 => "01011010",24587 => "00000000",24588 => "00001111",24589 => "00001101",24590 => "10010001",24591 => "00000111",24592 => "10001110",24593 => "10010101",24594 => "11101011",24595 => "11110010",24596 => "00110111",24597 => "11000011",24598 => "00011111",24599 => "10011100",24600 => "00010101",24601 => "01001111",24602 => "11001011",24603 => "10010101",24604 => "01110000",24605 => "00100110",24606 => "01011110",24607 => "11011111",24608 => "00000100",24609 => "00110010",24610 => "01101000",24611 => "10101100",24612 => "01101101",24613 => "00010000",24614 => "10101100",24615 => "10101010",24616 => "01001001",24617 => "10010010",24618 => "00001100",24619 => "01000110",24620 => "01011101",24621 => "11111001",24622 => "00001110",24623 => "11010110",24624 => "00111100",24625 => "11001111",24626 => "11010001",24627 => "10001010",24628 => "00011111",24629 => "00001100",24630 => "00011101",24631 => "11000101",24632 => "00111011",24633 => "01111111",24634 => "11010010",24635 => "11110011",24636 => "00000101",24637 => "11011100",24638 => "10110000",24639 => "11001011",24640 => "11101100",24641 => "00111010",24642 => "11011111",24643 => "10110101",24644 => "00111100",24645 => "00000101",24646 => "00010110",24647 => "01000111",24648 => "00011101",24649 => "11110101",24650 => "10111110",24651 => "11001001",24652 => "11000010",24653 => "01001110",24654 => "11111010",24655 => "00011001",24656 => "11101001",24657 => "10101001",24658 => "00110100",24659 => "11001001",24660 => "10001100",24661 => "11111101",24662 => "11000100",24663 => "10000000",24664 => "11001000",24665 => "11000110",24666 => "01000000",24667 => "11100110",24668 => "11111101",24669 => "10011101",24670 => "11000011",24671 => "10010000",24672 => "00011010",24673 => "00110010",24674 => "11100011",24675 => "10111011",24676 => "11011101",24677 => "11101001",24678 => "01001000",24679 => "01011100",24680 => "11011011",24681 => "01100011",24682 => "00001010",24683 => "11100100",24684 => "11011101",24685 => "10000110",24686 => "10110110",24687 => "00011011",24688 => "01100010",24689 => "11100001",24690 => "00000111",24691 => "00000010",24692 => "10110101",24693 => "01001010",24694 => "00010010",24695 => "11101110",24696 => "01001000",24697 => "10100111",24698 => "10101111",24699 => "01011110",24700 => "00110100",24701 => "10101111",24702 => "11101011",24703 => "00110100",24704 => "01010111",24705 => "10111001",24706 => "01100001",24707 => "11011111",24708 => "01100100",24709 => "01010110",24710 => "00010111",24711 => "10110110",24712 => "01111110",24713 => "10010110",24714 => "00011111",24715 => "00101101",24716 => "10100011",24717 => "10101100",24718 => "01000100",24719 => "00100010",24720 => "10110101",24721 => "10001000",24722 => "11011001",24723 => "01010011",24724 => "11100011",24725 => "10101100",24726 => "11100011",24727 => "10011111",24728 => "01010000",24729 => "01000001",24730 => "00110100",24731 => "10010011",24732 => "11100101",24733 => "10111101",24734 => "00011101",24735 => "11000010",24736 => "10110001",24737 => "10110011",24738 => "00101011",24739 => "10000000",24740 => "10100111",24741 => "11010111",24742 => "10111011",24743 => "11110001",24744 => "00100001",24745 => "11000000",24746 => "10100110",24747 => "00011000",24748 => "01100010",24749 => "01011010",24750 => "00000001",24751 => "01111010",24752 => "00101100",24753 => "01011100",24754 => "10100111",24755 => "00110001",24756 => "10111110",24757 => "10000000",24758 => "11101111",24759 => "00100101",24760 => "00101110",24761 => "00010101",24762 => "01000110",24763 => "00100010",24764 => "11000111",24765 => "01001011",24766 => "01101001",24767 => "11011001",24768 => "11000101",24769 => "11011110",24770 => "01101011",24771 => "01101101",24772 => "01010001",24773 => "00110001",24774 => "10101111",24775 => "11101110",24776 => "10101100",24777 => "11101111",24778 => "10101110",24779 => "11100101",24780 => "01100100",24781 => "01001111",24782 => "11010010",24783 => "11100111",24784 => "01001000",24785 => "10011100",24786 => "11000001",24787 => "10100001",24788 => "10001001",24789 => "01101111",24790 => "10100111",24791 => "11100111",24792 => "10010100",24793 => "01000110",24794 => "00110111",24795 => "10010100",24796 => "00110110",24797 => "01101001",24798 => "11101101",24799 => "01101101",24800 => "11011000",24801 => "11011110",24802 => "10011010",24803 => "10010001",24804 => "10010011",24805 => "10010100",24806 => "10011101",24807 => "01100100",24808 => "00110101",24809 => "01100011",24810 => "10110000",24811 => "01010100",24812 => "00011010",24813 => "10000000",24814 => "10011111",24815 => "00001000",24816 => "01111100",24817 => "01111101",24818 => "11010000",24819 => "00101011",24820 => "11111001",24821 => "01001001",24822 => "10010001",24823 => "01100000",24824 => "10101101",24825 => "10111001",24826 => "01010111",24827 => "01000110",24828 => "01111011",24829 => "00010010",24830 => "11101110",24831 => "10010110",24832 => "00110110",24833 => "01011010",24834 => "10100011",24835 => "01100011",24836 => "01111011",24837 => "11111111",24838 => "11001001",24839 => "00011011",24840 => "11001000",24841 => "11101111",24842 => "10011101",24843 => "11001010",24844 => "00010110",24845 => "11101010",24846 => "10101101",24847 => "01000100",24848 => "01001011",24849 => "11110101",24850 => "10000111",24851 => "01001110",24852 => "10111011",24853 => "11001110",24854 => "00011011",24855 => "10010100",24856 => "00001001",24857 => "00001100",24858 => "01010001",24859 => "01100101",24860 => "00111101",24861 => "11010011",24862 => "11100010",24863 => "11100000",24864 => "00000011",24865 => "00101001",24866 => "00011100",24867 => "01001110",24868 => "11001100",24869 => "10010100",24870 => "11000111",24871 => "10000110",24872 => "10101000",24873 => "10110100",24874 => "10010010",24875 => "11100001",24876 => "01001111",24877 => "10001010",24878 => "01000110",24879 => "10000001",24880 => "01100010",24881 => "00011111",24882 => "01101101",24883 => "01110111",24884 => "00110011",24885 => "11000100",24886 => "00110001",24887 => "11110010",24888 => "10101000",24889 => "11111101",24890 => "11100000",24891 => "00100110",24892 => "10010100",24893 => "10111001",24894 => "01000111",24895 => "01100011",24896 => "10001111",24897 => "01001000",24898 => "10110011",24899 => "10000010",24900 => "10011100",24901 => "11111011",24902 => "00101011",24903 => "01011001",24904 => "10001011",24905 => "01011100",24906 => "00000011",24907 => "01001111",24908 => "11000111",24909 => "11101010",24910 => "10010111",24911 => "00010111",24912 => "00110110",24913 => "10101000",24914 => "01011011",24915 => "11101011",24916 => "11110011",24917 => "00110001",24918 => "10101101",24919 => "10111001",24920 => "00000100",24921 => "10011110",24922 => "01011110",24923 => "11101011",24924 => "01110101",24925 => "01000111",24926 => "11110011",24927 => "11001110",24928 => "11001101",24929 => "01100001",24930 => "00111011",24931 => "11100110",24932 => "01110000",24933 => "01100011",24934 => "11111010",24935 => "11001100",24936 => "01000111",24937 => "00000010",24938 => "10000100",24939 => "10001111",24940 => "10001000",24941 => "10010100",24942 => "00011001",24943 => "00000110",24944 => "11000001",24945 => "11111111",24946 => "01001010",24947 => "01000000",24948 => "10100110",24949 => "01010011",24950 => "11101101",24951 => "10111101",24952 => "11001111",24953 => "11010011",24954 => "10111100",24955 => "11101001",24956 => "00110011",24957 => "11010011",24958 => "00010101",24959 => "01111000",24960 => "10000011",24961 => "01000100",24962 => "11110101",24963 => "00011111",24964 => "11011011",24965 => "00110001",24966 => "00110100",24967 => "01010001",24968 => "10110010",24969 => "10000011",24970 => "10001000",24971 => "00111000",24972 => "00000110",24973 => "00100011",24974 => "10010010",24975 => "10111001",24976 => "01000100",24977 => "00110000",24978 => "00101101",24979 => "11110011",24980 => "10101111",24981 => "00110101",24982 => "00000011",24983 => "00010011",24984 => "10110111",24985 => "01100100",24986 => "01101010",24987 => "10010011",24988 => "11001000",24989 => "01110100",24990 => "01111111",24991 => "11011111",24992 => "10010110",24993 => "10100101",24994 => "00011001",24995 => "00011000",24996 => "01110010",24997 => "11011000",24998 => "11111011",24999 => "00001100",25000 => "11100111",25001 => "11101101",25002 => "00100001",25003 => "10011110",25004 => "01000000",25005 => "00010100",25006 => "01100101",25007 => "01100000",25008 => "01011001",25009 => "01111010",25010 => "00010001",25011 => "11010100",25012 => "00011101",25013 => "10001011",25014 => "11000000",25015 => "00001110",25016 => "01001010",25017 => "11000011",25018 => "01100010",25019 => "10101001",25020 => "01100001",25021 => "11000010",25022 => "01011111",25023 => "10110110",25024 => "00010101",25025 => "00000011",25026 => "01001001",25027 => "00100001",25028 => "11011100",25029 => "01100110",25030 => "10010000",25031 => "01010110",25032 => "00011011",25033 => "10111100",25034 => "11101001",25035 => "00110111",25036 => "00100100",25037 => "00010110",25038 => "01000100",25039 => "01100101",25040 => "01110001",25041 => "10011000",25042 => "01111100",25043 => "00111010",25044 => "00110001",25045 => "00000010",25046 => "01101000",25047 => "00010101",25048 => "00011111",25049 => "10110100",25050 => "11000101",25051 => "11011110",25052 => "11001000",25053 => "11011001",25054 => "00001000",25055 => "00101000",25056 => "01110111",25057 => "01011000",25058 => "11001011",25059 => "00111100",25060 => "01011000",25061 => "00111000",25062 => "01010001",25063 => "01101010",25064 => "00110011",25065 => "10101011",25066 => "01010010",25067 => "11001010",25068 => "00000000",25069 => "00010111",25070 => "11010001",25071 => "10001111",25072 => "01100100",25073 => "01101011",25074 => "10110011",25075 => "01011010",25076 => "11011100",25077 => "00010101",25078 => "01110110",25079 => "01110111",25080 => "11110001",25081 => "11110010",25082 => "00111111",25083 => "10100001",25084 => "00100100",25085 => "01001011",25086 => "01011111",25087 => "00101010",25088 => "11111110",25089 => "00101110",25090 => "10110000",25091 => "01000001",25092 => "00011011",25093 => "10000011",25094 => "01111111",25095 => "10001101",25096 => "10011001",25097 => "01100000",25098 => "00110010",25099 => "00011100",25100 => "11000001",25101 => "00011111",25102 => "01101000",25103 => "00001001",25104 => "11101001",25105 => "10111000",25106 => "01100110",25107 => "10001110",25108 => "11111111",25109 => "00011001",25110 => "00110011",25111 => "10101110",25112 => "00011100",25113 => "00011001",25114 => "00001000",25115 => "11110101",25116 => "11010101",25117 => "10110111",25118 => "11110001",25119 => "11100010",25120 => "11111101",25121 => "10111001",25122 => "10001110",25123 => "01100011",25124 => "01010100",25125 => "10110010",25126 => "00010100",25127 => "01010010",25128 => "10100000",25129 => "00000110",25130 => "11000110",25131 => "01010000",25132 => "11110010",25133 => "10101010",25134 => "10100011",25135 => "01000100",25136 => "00001101",25137 => "00111100",25138 => "10010001",25139 => "10011010",25140 => "10011101",25141 => "10111111",25142 => "00010100",25143 => "10001101",25144 => "11100001",25145 => "00101000",25146 => "00011011",25147 => "11101101",25148 => "01110000",25149 => "11100111",25150 => "01100001",25151 => "10011001",25152 => "00001010",25153 => "01001001",25154 => "10011010",25155 => "00010100",25156 => "11011100",25157 => "01110101",25158 => "00010000",25159 => "00011101",25160 => "11010001",25161 => "10100101",25162 => "10111001",25163 => "10100010",25164 => "10001111",25165 => "01001010",25166 => "11101010",25167 => "00101010",25168 => "11101001",25169 => "11101010",25170 => "01010100",25171 => "11011111",25172 => "10001010",25173 => "10000011",25174 => "10111010",25175 => "10011011",25176 => "11010100",25177 => "11001011",25178 => "00101110",25179 => "11110101",25180 => "01010111",25181 => "10111000",25182 => "10010001",25183 => "00110001",25184 => "00010000",25185 => "01110011",25186 => "00100110",25187 => "10010010",25188 => "11100100",25189 => "01000000",25190 => "11011000",25191 => "01011110",25192 => "01111000",25193 => "01101101",25194 => "10110100",25195 => "01001100",25196 => "10000010",25197 => "01110000",25198 => "11101100",25199 => "10110111",25200 => "11000011",25201 => "01011010",25202 => "10110011",25203 => "01010111",25204 => "10110111",25205 => "10110000",25206 => "10110110",25207 => "10011111",25208 => "00101100",25209 => "10111101",25210 => "10000110",25211 => "10011111",25212 => "01100101",25213 => "00000110",25214 => "01010010",25215 => "11001111",25216 => "10111101",25217 => "11101101",25218 => "10011011",25219 => "00110101",25220 => "01010011",25221 => "01101101",25222 => "00011011",25223 => "10101011",25224 => "11100101",25225 => "10011000",25226 => "11101101",25227 => "10000110",25228 => "11001011",25229 => "10001101",25230 => "01001010",25231 => "00001110",25232 => "10110100",25233 => "00110110",25234 => "00111001",25235 => "00000000",25236 => "01000101",25237 => "00010010",25238 => "11100001",25239 => "00011110",25240 => "10110010",25241 => "11001110",25242 => "00111010",25243 => "10101101",25244 => "11101111",25245 => "10001101",25246 => "01011011",25247 => "11000000",25248 => "11000001",25249 => "11001011",25250 => "00000100",25251 => "01101010",25252 => "11001000",25253 => "10101101",25254 => "10000000",25255 => "11011010",25256 => "00000111",25257 => "01100011",25258 => "10000011",25259 => "00111110",25260 => "10111011",25261 => "00000101",25262 => "01010100",25263 => "01000001",25264 => "11101001",25265 => "10000010",25266 => "11100111",25267 => "10100000",25268 => "00111111",25269 => "11101001",25270 => "11111100",25271 => "10010100",25272 => "11001010",25273 => "11010111",25274 => "00101111",25275 => "11000111",25276 => "00001001",25277 => "10011101",25278 => "11001010",25279 => "10010100",25280 => "01010001",25281 => "10000111",25282 => "01110000",25283 => "10110000",25284 => "01101100",25285 => "01010010",25286 => "10000111",25287 => "01010101",25288 => "10000011",25289 => "01110110",25290 => "10011111",25291 => "11100101",25292 => "10101011",25293 => "10101000",25294 => "00001100",25295 => "10100101",25296 => "00001111",25297 => "01001010",25298 => "00011111",25299 => "10110010",25300 => "00010001",25301 => "10110110",25302 => "10001100",25303 => "01001010",25304 => "01110111",25305 => "11101001",25306 => "01111101",25307 => "11111101",25308 => "00000011",25309 => "01100100",25310 => "00010111",25311 => "00100001",25312 => "00111111",25313 => "10011010",25314 => "01010010",25315 => "00111001",25316 => "01010111",25317 => "11010110",25318 => "10101111",25319 => "01110010",25320 => "01110111",25321 => "01010100",25322 => "00100110",25323 => "11100001",25324 => "00010001",25325 => "10100111",25326 => "01111110",25327 => "11001100",25328 => "01100010",25329 => "00010110",25330 => "10100110",25331 => "10111101",25332 => "01111011",25333 => "11100001",25334 => "11011101",25335 => "00011111",25336 => "01110011",25337 => "00001110",25338 => "01110110",25339 => "00100110",25340 => "00101001",25341 => "10001001",25342 => "11001101",25343 => "11110101",25344 => "11011010",25345 => "01011100",25346 => "11110000",25347 => "00010010",25348 => "00101111",25349 => "00000110",25350 => "01000001",25351 => "01111010",25352 => "10110011",25353 => "01001111",25354 => "00110011",25355 => "00100011",25356 => "11110001",25357 => "01111011",25358 => "01100111",25359 => "01011110",25360 => "11111101",25361 => "10111000",25362 => "01000011",25363 => "01101011",25364 => "00001000",25365 => "10100111",25366 => "00001010",25367 => "10001010",25368 => "10101110",25369 => "00011110",25370 => "00110000",25371 => "01010001",25372 => "01100100",25373 => "00101110",25374 => "10000000",25375 => "01100111",25376 => "11100000",25377 => "00111001",25378 => "11110001",25379 => "11111011",25380 => "00010100",25381 => "10110100",25382 => "11100111",25383 => "10011110",25384 => "11110001",25385 => "10101101",25386 => "01010011",25387 => "10011000",25388 => "10011011",25389 => "00111101",25390 => "11000010",25391 => "11010100",25392 => "10111101",25393 => "01001111",25394 => "10111111",25395 => "11011110",25396 => "00000011",25397 => "00001011",25398 => "00110011",25399 => "01110011",25400 => "00101010",25401 => "00110111",25402 => "11110110",25403 => "11110010",25404 => "10011011",25405 => "11011111",25406 => "00011010",25407 => "11000000",25408 => "01100101",25409 => "11111111",25410 => "10001100",25411 => "01101011",25412 => "01111001",25413 => "10001011",25414 => "01001011",25415 => "11111100",25416 => "10011001",25417 => "10110111",25418 => "11011010",25419 => "00000111",25420 => "00001111",25421 => "01110110",25422 => "01001001",25423 => "00000001",25424 => "11100110",25425 => "00101111",25426 => "11001111",25427 => "11011001",25428 => "01011011",25429 => "00001101",25430 => "01111100",25431 => "11110001",25432 => "10011111",25433 => "01100101",25434 => "11101110",25435 => "01101000",25436 => "01010011",25437 => "11000101",25438 => "00011000",25439 => "10100110",25440 => "11100011",25441 => "00011000",25442 => "10000110",25443 => "00100001",25444 => "10111110",25445 => "00110101",25446 => "10000110",25447 => "01010111",25448 => "00011110",25449 => "11000101",25450 => "00001001",25451 => "11111111",25452 => "10111100",25453 => "01111100",25454 => "01001111",25455 => "11100101",25456 => "11011001",25457 => "01100001",25458 => "00110010",25459 => "00010110",25460 => "11010000",25461 => "00111001",25462 => "00101100",25463 => "11100101",25464 => "11111101",25465 => "00011101",25466 => "00001010",25467 => "11100000",25468 => "01101110",25469 => "10001101",25470 => "00000101",25471 => "11010001",25472 => "11110110",25473 => "10111100",25474 => "00100010",25475 => "11100010",25476 => "00100111",25477 => "00100101",25478 => "01010011",25479 => "11101100",25480 => "01100110",25481 => "10010001",25482 => "01010101",25483 => "00001000",25484 => "10001100",25485 => "00010001",25486 => "01001001",25487 => "11100011",25488 => "00010010",25489 => "01101110",25490 => "11011110",25491 => "11101100",25492 => "00000010",25493 => "00001000",25494 => "10110100",25495 => "10111011",25496 => "11011010",25497 => "10011111",25498 => "11011010",25499 => "01110111",25500 => "11101111",25501 => "01100011",25502 => "10100001",25503 => "01111000",25504 => "00011000",25505 => "11000111",25506 => "01110111",25507 => "11111010",25508 => "00111100",25509 => "01111011",25510 => "00111011",25511 => "11010000",25512 => "11011110",25513 => "01001111",25514 => "01000101",25515 => "10101010",25516 => "00110111",25517 => "11011110",25518 => "00110100",25519 => "10100101",25520 => "11001100",25521 => "00101000",25522 => "00001111",25523 => "11111000",25524 => "00101011",25525 => "00010001",25526 => "00000011",25527 => "11010001",25528 => "11011101",25529 => "01010000",25530 => "00100110",25531 => "11000101",25532 => "01100111",25533 => "00000011",25534 => "00101110",25535 => "10101110",25536 => "00111110",25537 => "10001100",25538 => "10100001",25539 => "00001001",25540 => "10100000",25541 => "11010100",25542 => "10110101",25543 => "00111110",25544 => "00101100",25545 => "00000011",25546 => "11110101",25547 => "11001111",25548 => "01100101",25549 => "10001111",25550 => "01101110",25551 => "11111000",25552 => "00111100",25553 => "11000111",25554 => "10111000",25555 => "01001000",25556 => "11000111",25557 => "10010011",25558 => "10000100",25559 => "00010011",25560 => "01011010",25561 => "00011111",25562 => "00101010",25563 => "00011010",25564 => "01101110",25565 => "10000011",25566 => "00101001",25567 => "01000010",25568 => "00100011",25569 => "10111000",25570 => "00011100",25571 => "10101000",25572 => "10011001",25573 => "00011100",25574 => "01110110",25575 => "11101111",25576 => "01011001",25577 => "11011011",25578 => "01101001",25579 => "11010011",25580 => "01001000",25581 => "00111011",25582 => "10001100",25583 => "01000001",25584 => "00110100",25585 => "10010010",25586 => "11100010",25587 => "11111100",25588 => "00000110",25589 => "00010010",25590 => "01100011",25591 => "00011111",25592 => "01111100",25593 => "00111100",25594 => "01011011",25595 => "11011111",25596 => "01110011",25597 => "00111111",25598 => "01110110",25599 => "00001100",25600 => "01000111",25601 => "00101101",25602 => "01110001",25603 => "01100011",25604 => "10001011",25605 => "10000111",25606 => "10000011",25607 => "01101101",25608 => "00111110",25609 => "00100011",25610 => "00010111",25611 => "01101110",25612 => "10111001",25613 => "01010011",25614 => "11101010",25615 => "11001101",25616 => "01110100",25617 => "11111100",25618 => "11010011",25619 => "00010110",25620 => "10111101",25621 => "00010010",25622 => "11000010",25623 => "10010100",25624 => "01101110",25625 => "00110010",25626 => "01110100",25627 => "00000100",25628 => "00111000",25629 => "10110111",25630 => "01011111",25631 => "00001010",25632 => "00000110",25633 => "11001110",25634 => "01110010",25635 => "01110111",25636 => "10111110",25637 => "11001100",25638 => "00000001",25639 => "00000011",25640 => "10010001",25641 => "01110111",25642 => "00101011",25643 => "10100011",25644 => "00110101",25645 => "10100000",25646 => "00111110",25647 => "01010010",25648 => "00100000",25649 => "01100000",25650 => "00110111",25651 => "10000110",25652 => "10101000",25653 => "00110101",25654 => "01010101",25655 => "10000000",25656 => "00000010",25657 => "11011110",25658 => "00001111",25659 => "00001010",25660 => "10110010",25661 => "11111011",25662 => "10111111",25663 => "10111001",25664 => "00101101",25665 => "11011111",25666 => "00100101",25667 => "00111001",25668 => "01010010",25669 => "00000100",25670 => "10111110",25671 => "11010111",25672 => "11111110",25673 => "10100110",25674 => "01110001",25675 => "00110010",25676 => "10111110",25677 => "01111001",25678 => "10011110",25679 => "11010110",25680 => "11101110",25681 => "10010011",25682 => "00100101",25683 => "00000101",25684 => "01101111",25685 => "11011011",25686 => "10101000",25687 => "11101110",25688 => "10010111",25689 => "01110110",25690 => "10000001",25691 => "00101101",25692 => "10110111",25693 => "01110101",25694 => "11010101",25695 => "01101111",25696 => "00101001",25697 => "10111100",25698 => "11110100",25699 => "00010001",25700 => "11001000",25701 => "00111100",25702 => "10111101",25703 => "00010111",25704 => "01110111",25705 => "01001001",25706 => "11100011",25707 => "11000101",25708 => "00000001",25709 => "01000110",25710 => "01101110",25711 => "10011000",25712 => "11000101",25713 => "11110001",25714 => "11000101",25715 => "00010010",25716 => "00100100",25717 => "11010111",25718 => "01110110",25719 => "11100001",25720 => "01101000",25721 => "01110010",25722 => "00010011",25723 => "11111010",25724 => "11000001",25725 => "11001001",25726 => "00000000",25727 => "11011011",25728 => "10001010",25729 => "11101110",25730 => "10111001",25731 => "10100111",25732 => "11000110",25733 => "11011001",25734 => "11100011",25735 => "01101101",25736 => "01011000",25737 => "01000111",25738 => "01000011",25739 => "00000011",25740 => "11111010",25741 => "00001110",25742 => "00001010",25743 => "00011001",25744 => "01110000",25745 => "11000011",25746 => "10101100",25747 => "10110010",25748 => "01010000",25749 => "01111111",25750 => "01101011",25751 => "10000011",25752 => "00101000",25753 => "00010111",25754 => "01000011",25755 => "11000010",25756 => "10101110",25757 => "10000100",25758 => "00110011",25759 => "10000000",25760 => "01010100",25761 => "11101110",25762 => "11010100",25763 => "10011001",25764 => "11100110",25765 => "11100111",25766 => "11000011",25767 => "01100110",25768 => "10001011",25769 => "10011001",25770 => "01000111",25771 => "11111011",25772 => "01010101",25773 => "01100100",25774 => "00010001",25775 => "01010000",25776 => "00101100",25777 => "10111111",25778 => "11111010",25779 => "10011101",25780 => "10110110",25781 => "10011100",25782 => "11110001",25783 => "01101011",25784 => "00110110",25785 => "11100000",25786 => "11100111",25787 => "11101010",25788 => "00111010",25789 => "00011001",25790 => "11101011",25791 => "01100101",25792 => "01110111",25793 => "00010111",25794 => "00000100",25795 => "11101111",25796 => "11000101",25797 => "10100011",25798 => "11011100",25799 => "00111000",25800 => "10110100",25801 => "00011001",25802 => "01111101",25803 => "10001101",25804 => "01010101",25805 => "00101011",25806 => "00110100",25807 => "11000100",25808 => "01000110",25809 => "01111010",25810 => "01100101",25811 => "01000000",25812 => "00011010",25813 => "00100000",25814 => "11100010",25815 => "11011000",25816 => "00110001",25817 => "10000111",25818 => "00111101",25819 => "10100101",25820 => "11100101",25821 => "10100011",25822 => "01100000",25823 => "10101101",25824 => "00000011",25825 => "01011110",25826 => "11001110",25827 => "01001100",25828 => "01000000",25829 => "01011011",25830 => "11111110",25831 => "11110000",25832 => "01010110",25833 => "01010110",25834 => "01111100",25835 => "01010101",25836 => "00111111",25837 => "11001110",25838 => "01010011",25839 => "00100000",25840 => "00011101",25841 => "01101011",25842 => "01111100",25843 => "11100000",25844 => "00100001",25845 => "01000011",25846 => "01100110",25847 => "11001000",25848 => "11000110",25849 => "11000110",25850 => "10110100",25851 => "01111000",25852 => "11100101",25853 => "11100000",25854 => "11011111",25855 => "01100010",25856 => "10011000",25857 => "10011001",25858 => "10101100",25859 => "11011010",25860 => "01010001",25861 => "11100101",25862 => "01110111",25863 => "10111011",25864 => "01101011",25865 => "10111111",25866 => "11010010",25867 => "01011001",25868 => "01001001",25869 => "00101000",25870 => "11110101",25871 => "10011101",25872 => "10101100",25873 => "11110010",25874 => "11111100",25875 => "00000100",25876 => "00001111",25877 => "00101100",25878 => "11001101",25879 => "01101111",25880 => "11101110",25881 => "01001110",25882 => "00111101",25883 => "11110101",25884 => "01000110",25885 => "01111001",25886 => "10010011",25887 => "01110101",25888 => "01110101",25889 => "10000010",25890 => "01001101",25891 => "10100001",25892 => "11010000",25893 => "01111110",25894 => "11100001",25895 => "00010100",25896 => "10101111",25897 => "00110111",25898 => "10010000",25899 => "01101100",25900 => "10101011",25901 => "11110010",25902 => "10111101",25903 => "01000101",25904 => "01111111",25905 => "10011001",25906 => "00110101",25907 => "00111100",25908 => "00100011",25909 => "00001100",25910 => "00011111",25911 => "00100011",25912 => "10101011",25913 => "11111111",25914 => "01010111",25915 => "10000100",25916 => "00000000",25917 => "00100100",25918 => "01110000",25919 => "11100101",25920 => "01011100",25921 => "01111110",25922 => "00101101",25923 => "01111100",25924 => "10010001",25925 => "00011000",25926 => "11000000",25927 => "00011011",25928 => "01111011",25929 => "10011100",25930 => "11001101",25931 => "10101100",25932 => "01110110",25933 => "11100011",25934 => "11010011",25935 => "00101100",25936 => "01101000",25937 => "11011111",25938 => "11011001",25939 => "00101111",25940 => "01011101",25941 => "01110011",25942 => "11010011",25943 => "10011100",25944 => "00100000",25945 => "00111100",25946 => "01001100",25947 => "00111000",25948 => "10100011",25949 => "10100011",25950 => "00110000",25951 => "01001001",25952 => "10101001",25953 => "01000001",25954 => "00001100",25955 => "00010100",25956 => "00000001",25957 => "01110111",25958 => "10000100",25959 => "01001110",25960 => "00110100",25961 => "00011111",25962 => "10111001",25963 => "11010010",25964 => "00010010",25965 => "11100000",25966 => "10111110",25967 => "01000111",25968 => "00111011",25969 => "01111001",25970 => "00110010",25971 => "01000010",25972 => "11101001",25973 => "11000111",25974 => "11100011",25975 => "11001010",25976 => "10110100",25977 => "00110101",25978 => "10000100",25979 => "01001100",25980 => "01011000",25981 => "00110111",25982 => "11111010",25983 => "00110100",25984 => "11111010",25985 => "00001001",25986 => "01011101",25987 => "01110111",25988 => "11101100",25989 => "01011001",25990 => "10000001",25991 => "01010011",25992 => "10101111",25993 => "11110100",25994 => "01001000",25995 => "00111110",25996 => "00111110",25997 => "00000000",25998 => "10000100",25999 => "11100111",26000 => "01000001",26001 => "00100110",26002 => "01110111",26003 => "00101111",26004 => "01000101",26005 => "01101001",26006 => "00101110",26007 => "11010010",26008 => "11000111",26009 => "00011000",26010 => "01101111",26011 => "00110011",26012 => "10001101",26013 => "10000010",26014 => "10110010",26015 => "01110000",26016 => "10101001",26017 => "01111110",26018 => "10010011",26019 => "00100000",26020 => "00101000",26021 => "01100101",26022 => "11101111",26023 => "10101011",26024 => "10010110",26025 => "11000111",26026 => "11010100",26027 => "00011100",26028 => "00111001",26029 => "01001000",26030 => "10101011",26031 => "01101011",26032 => "11001111",26033 => "10001011",26034 => "00110011",26035 => "11010011",26036 => "11010100",26037 => "10101000",26038 => "10101001",26039 => "01000101",26040 => "00110010",26041 => "11011100",26042 => "11001010",26043 => "10000010",26044 => "01011101",26045 => "11001101",26046 => "01001111",26047 => "01000111",26048 => "10111000",26049 => "10001010",26050 => "10011001",26051 => "01111011",26052 => "11100110",26053 => "10001101",26054 => "00001101",26055 => "10001110",26056 => "01010100",26057 => "00101010",26058 => "10111101",26059 => "01110011",26060 => "10001100",26061 => "01001111",26062 => "10111110",26063 => "00100000",26064 => "11110100",26065 => "01010010",26066 => "01111110",26067 => "01010010",26068 => "01111111",26069 => "01011010",26070 => "01111011",26071 => "10100110",26072 => "10101011",26073 => "01010010",26074 => "11100101",26075 => "10010111",26076 => "10100101",26077 => "10001000",26078 => "00101100",26079 => "11110000",26080 => "10000011",26081 => "00110000",26082 => "01100100",26083 => "01111011",26084 => "00000100",26085 => "00101011",26086 => "11000010",26087 => "11011101",26088 => "11111011",26089 => "11011100",26090 => "10011010",26091 => "10001101",26092 => "10111110",26093 => "01010001",26094 => "10101000",26095 => "11110010",26096 => "10110001",26097 => "11000110",26098 => "00001011",26099 => "00010110",26100 => "11001000",26101 => "01011110",26102 => "00111011",26103 => "01000010",26104 => "01011011",26105 => "01011001",26106 => "11001001",26107 => "00010100",26108 => "11011011",26109 => "11101100",26110 => "00110010",26111 => "00011101",26112 => "11000011",26113 => "00111111",26114 => "10111101",26115 => "10101011",26116 => "00011011",26117 => "10010101",26118 => "01100000",26119 => "10101000",26120 => "01111101",26121 => "01000010",26122 => "00010010",26123 => "00000001",26124 => "00101010",26125 => "11000101",26126 => "11111100",26127 => "01000111",26128 => "01001111",26129 => "11011100",26130 => "01101010",26131 => "11110101",26132 => "11101010",26133 => "11100101",26134 => "01100011",26135 => "01110000",26136 => "10111101",26137 => "10001001",26138 => "10101001",26139 => "01101111",26140 => "11101111",26141 => "10000010",26142 => "01001111",26143 => "10101101",26144 => "01111111",26145 => "11001111",26146 => "01010111",26147 => "11100011",26148 => "01101011",26149 => "01101100",26150 => "10111011",26151 => "01110110",26152 => "01011100",26153 => "00110101",26154 => "11111101",26155 => "10000011",26156 => "11011010",26157 => "11011000",26158 => "10011101",26159 => "10111010",26160 => "00010111",26161 => "10101110",26162 => "00110100",26163 => "11110111",26164 => "11001111",26165 => "10001010",26166 => "01001011",26167 => "00101111",26168 => "11110110",26169 => "00110001",26170 => "11011011",26171 => "11100010",26172 => "01111111",26173 => "01001010",26174 => "11100110",26175 => "10001000",26176 => "10100100",26177 => "01111110",26178 => "11011010",26179 => "01111111",26180 => "11001010",26181 => "10100011",26182 => "10110000",26183 => "11111001",26184 => "01100010",26185 => "10010001",26186 => "10000100",26187 => "11010011",26188 => "00101001",26189 => "01100111",26190 => "10100011",26191 => "00100100",26192 => "10100010",26193 => "11110011",26194 => "11011000",26195 => "01011111",26196 => "10001000",26197 => "10100001",26198 => "10011110",26199 => "10101001",26200 => "11110111",26201 => "11110000",26202 => "11010000",26203 => "10100001",26204 => "11101111",26205 => "10100101",26206 => "01101100",26207 => "10010011",26208 => "01011110",26209 => "10111001",26210 => "01110101",26211 => "01000100",26212 => "11011010",26213 => "10011001",26214 => "10010001",26215 => "01000110",26216 => "10000100",26217 => "00001101",26218 => "00110110",26219 => "01011000",26220 => "01000101",26221 => "00110110",26222 => "11011011",26223 => "00001110",26224 => "00000100",26225 => "11100001",26226 => "01110011",26227 => "11000001",26228 => "11010010",26229 => "01111000",26230 => "01010010",26231 => "01001011",26232 => "10000011",26233 => "01101101",26234 => "11110101",26235 => "11000000",26236 => "00010100",26237 => "11100101",26238 => "11110100",26239 => "01001000",26240 => "00001111",26241 => "00111111",26242 => "01100100",26243 => "10001000",26244 => "00010010",26245 => "00111111",26246 => "10100001",26247 => "01000010",26248 => "01000100",26249 => "00010010",26250 => "10110001",26251 => "11011001",26252 => "00010011",26253 => "10100000",26254 => "11011101",26255 => "10000011",26256 => "01101101",26257 => "01110110",26258 => "00000010",26259 => "00001110",26260 => "01101000",26261 => "00111100",26262 => "01001111",26263 => "11010001",26264 => "10010001",26265 => "01011101",26266 => "00000111",26267 => "00101001",26268 => "11111100",26269 => "00000011",26270 => "11100000",26271 => "10111110",26272 => "11001001",26273 => "00000101",26274 => "11110100",26275 => "10011100",26276 => "00110100",26277 => "00101000",26278 => "10101101",26279 => "10000110",26280 => "00010000",26281 => "01010101",26282 => "11100111",26283 => "10110011",26284 => "00111010",26285 => "01001100",26286 => "00101011",26287 => "01001111",26288 => "01000011",26289 => "00111000",26290 => "11001001",26291 => "10110111",26292 => "00011010",26293 => "00111110",26294 => "01101100",26295 => "11111100",26296 => "10011110",26297 => "00100100",26298 => "01000101",26299 => "10101011",26300 => "11011111",26301 => "01001101",26302 => "01001101",26303 => "11010011",26304 => "10101000",26305 => "01111100",26306 => "11101111",26307 => "10000100",26308 => "10011111",26309 => "01110111",26310 => "01101011",26311 => "11011001",26312 => "10101110",26313 => "00111000",26314 => "10111100",26315 => "11010101",26316 => "10000111",26317 => "11110111",26318 => "00010000",26319 => "10000001",26320 => "01110011",26321 => "10110000",26322 => "10100011",26323 => "10110011",26324 => "01101111",26325 => "00110000",26326 => "10000110",26327 => "00011010",26328 => "10000111",26329 => "00011011",26330 => "01101100",26331 => "01010001",26332 => "01100000",26333 => "10110000",26334 => "00010010",26335 => "11110011",26336 => "10101001",26337 => "01000111",26338 => "01011110",26339 => "01011101",26340 => "10100110",26341 => "11011111",26342 => "00001010",26343 => "11000110",26344 => "01101100",26345 => "10110101",26346 => "11110111",26347 => "11001011",26348 => "11110010",26349 => "11110010",26350 => "10010011",26351 => "01000011",26352 => "10010110",26353 => "01110101",26354 => "01001100",26355 => "01110101",26356 => "10011000",26357 => "00110110",26358 => "10100010",26359 => "01011011",26360 => "01111000",26361 => "01110000",26362 => "00101100",26363 => "11001100",26364 => "10110010",26365 => "00000111",26366 => "01100110",26367 => "10100011",26368 => "11010101",26369 => "00011001",26370 => "01100111",26371 => "01010110",26372 => "11111100",26373 => "11000111",26374 => "10001111",26375 => "01001111",26376 => "01100011",26377 => "01011111",26378 => "01000011",26379 => "10100110",26380 => "01001010",26381 => "01100011",26382 => "00110010",26383 => "11011100",26384 => "11101100",26385 => "01001011",26386 => "11010010",26387 => "01111000",26388 => "01101101",26389 => "01101110",26390 => "01011101",26391 => "01100101",26392 => "10001011",26393 => "10100011",26394 => "10111101",26395 => "00011100",26396 => "11101101",26397 => "00101011",26398 => "00100111",26399 => "11111110",26400 => "11001011",26401 => "01101010",26402 => "11110010",26403 => "11110110",26404 => "01110011",26405 => "10000111",26406 => "10101000",26407 => "00110011",26408 => "11011101",26409 => "01000111",26410 => "10010010",26411 => "01101110",26412 => "01001001",26413 => "11001101",26414 => "10101000",26415 => "01001010",26416 => "01000011",26417 => "00010101",26418 => "01101010",26419 => "00000010",26420 => "01001011",26421 => "11111111",26422 => "01110100",26423 => "01001001",26424 => "11101010",26425 => "00001101",26426 => "00001101",26427 => "01000100",26428 => "01001110",26429 => "10010101",26430 => "11100100",26431 => "10011001",26432 => "00101110",26433 => "01011111",26434 => "00111101",26435 => "00111000",26436 => "10011011",26437 => "10010011",26438 => "11100101",26439 => "10001010",26440 => "10000100",26441 => "10010000",26442 => "11100111",26443 => "01011111",26444 => "01001100",26445 => "00111010",26446 => "01010101",26447 => "11101110",26448 => "10000001",26449 => "10110111",26450 => "10000010",26451 => "11000010",26452 => "11110100",26453 => "11111111",26454 => "11010001",26455 => "11000001",26456 => "11101110",26457 => "00011101",26458 => "10100111",26459 => "01000001",26460 => "10111010",26461 => "00000111",26462 => "11000011",26463 => "01010000",26464 => "11100110",26465 => "11000111",26466 => "01110101",26467 => "00000111",26468 => "00001110",26469 => "11000011",26470 => "00100100",26471 => "00011011",26472 => "00001110",26473 => "01111000",26474 => "10101111",26475 => "00100001",26476 => "11101111",26477 => "00100101",26478 => "10010010",26479 => "10001000",26480 => "10110110",26481 => "11010101",26482 => "00111100",26483 => "01111010",26484 => "00011001",26485 => "01101100",26486 => "10001100",26487 => "11000000",26488 => "10011100",26489 => "10011101",26490 => "00001010",26491 => "11111001",26492 => "11000101",26493 => "10111111",26494 => "00010001",26495 => "01011001",26496 => "00101101",26497 => "00100110",26498 => "01011000",26499 => "00111011",26500 => "00110110",26501 => "00001111",26502 => "00101101",26503 => "01111000",26504 => "11001010",26505 => "00001001",26506 => "00011101",26507 => "11011001",26508 => "11001110",26509 => "10000010",26510 => "01101000",26511 => "00001111",26512 => "10011010",26513 => "01111010",26514 => "01100001",26515 => "00011011",26516 => "11011111",26517 => "10011001",26518 => "10101010",26519 => "10111110",26520 => "10111000",26521 => "10111100",26522 => "11011000",26523 => "10111010",26524 => "11001111",26525 => "10001010",26526 => "10000110",26527 => "00101010",26528 => "11100001",26529 => "11101000",26530 => "00000101",26531 => "10011010",26532 => "01011010",26533 => "01010100",26534 => "10011111",26535 => "11001111",26536 => "11000001",26537 => "11111110",26538 => "01110001",26539 => "11000111",26540 => "10111110",26541 => "01001010",26542 => "01001111",26543 => "10001101",26544 => "11110011",26545 => "10100010",26546 => "10000111",26547 => "01011100",26548 => "10000000",26549 => "11100000",26550 => "00100111",26551 => "10110110",26552 => "01110000",26553 => "10101000",26554 => "00011101",26555 => "01000011",26556 => "11100011",26557 => "10011101",26558 => "11001111",26559 => "01010000",26560 => "00000111",26561 => "11000010",26562 => "00000100",26563 => "01000100",26564 => "10110110",26565 => "11101111",26566 => "01101000",26567 => "10001000",26568 => "00000111",26569 => "11001101",26570 => "00100001",26571 => "10100110",26572 => "10101101",26573 => "00100100",26574 => "11011011",26575 => "10100101",26576 => "10111100",26577 => "10000101",26578 => "10110011",26579 => "10011111",26580 => "01011110",26581 => "00011100",26582 => "10010011",26583 => "11010000",26584 => "10101011",26585 => "11100000",26586 => "00101001",26587 => "00001011",26588 => "10110111",26589 => "11110010",26590 => "01011000",26591 => "01110101",26592 => "01111100",26593 => "01111100",26594 => "01001100",26595 => "01101011",26596 => "11111011",26597 => "11001000",26598 => "00001001",26599 => "00111110",26600 => "10100100",26601 => "00110100",26602 => "10110100",26603 => "00001101",26604 => "01011000",26605 => "10100110",26606 => "11011010",26607 => "00000001",26608 => "01101110",26609 => "00111100",26610 => "10010110",26611 => "10011000",26612 => "10010110",26613 => "10101000",26614 => "11011110",26615 => "01101111",26616 => "01111011",26617 => "01000001",26618 => "10000010",26619 => "00010111",26620 => "10000110",26621 => "01011000",26622 => "00010000",26623 => "00101111",26624 => "00100100",26625 => "11100101",26626 => "00011011",26627 => "10010000",26628 => "10001000",26629 => "11110010",26630 => "11000010",26631 => "01101110",26632 => "10110001",26633 => "01101111",26634 => "10101010",26635 => "11010001",26636 => "01001100",26637 => "10100010",26638 => "01011111",26639 => "00010011",26640 => "01000101",26641 => "10111110",26642 => "00000100",26643 => "00010000",26644 => "11100010",26645 => "11110011",26646 => "01111101",26647 => "00111010",26648 => "00101000",26649 => "10000010",26650 => "11110110",26651 => "11100001",26652 => "01110111",26653 => "10010000",26654 => "10001100",26655 => "11110111",26656 => "10100110",26657 => "10110000",26658 => "10101110",26659 => "00000010",26660 => "00110111",26661 => "11001011",26662 => "01011110",26663 => "00000000",26664 => "10001111",26665 => "01111111",26666 => "00111011",26667 => "10101011",26668 => "10011010",26669 => "00100001",26670 => "01111010",26671 => "01000010",26672 => "10111010",26673 => "00011000",26674 => "01001001",26675 => "11111010",26676 => "11101101",26677 => "01100101",26678 => "00000110",26679 => "01011100",26680 => "10000111",26681 => "00001010",26682 => "01101110",26683 => "11000011",26684 => "11100010",26685 => "11011001",26686 => "11110000",26687 => "01101111",26688 => "00011100",26689 => "11010011",26690 => "11111110",26691 => "00111110",26692 => "00111101",26693 => "01111010",26694 => "00001101",26695 => "11010100",26696 => "10011000",26697 => "11000100",26698 => "01110100",26699 => "11111110",26700 => "10100101",26701 => "00011011",26702 => "01101110",26703 => "11110001",26704 => "10101100",26705 => "01101000",26706 => "00111001",26707 => "00000011",26708 => "11001010",26709 => "00001001",26710 => "10011100",26711 => "01101000",26712 => "11111000",26713 => "11011001",26714 => "01111100",26715 => "10001011",26716 => "00010101",26717 => "10000001",26718 => "10001001",26719 => "11011000",26720 => "10001000",26721 => "01011100",26722 => "10111001",26723 => "11010011",26724 => "11000000",26725 => "00100101",26726 => "01110011",26727 => "11001101",26728 => "11111000",26729 => "11001001",26730 => "01100100",26731 => "01101100",26732 => "01000001",26733 => "00110101",26734 => "11001110",26735 => "00100011",26736 => "10001010",26737 => "00011011",26738 => "01001101",26739 => "10000111",26740 => "10110101",26741 => "01111100",26742 => "01101110",26743 => "00101011",26744 => "11000011",26745 => "11001001",26746 => "11100111",26747 => "01001011",26748 => "11101010",26749 => "11011101",26750 => "00010010",26751 => "10100010",26752 => "10101100",26753 => "11110001",26754 => "11000000",26755 => "00001001",26756 => "11110010",26757 => "01101010",26758 => "00001110",26759 => "11001100",26760 => "10000111",26761 => "10111001",26762 => "10100100",26763 => "10011100",26764 => "11110101",26765 => "11111001",26766 => "11011001",26767 => "01011011",26768 => "10001100",26769 => "00011101",26770 => "01111001",26771 => "10011100",26772 => "00000111",26773 => "10100000",26774 => "01110010",26775 => "10111001",26776 => "00010001",26777 => "01101100",26778 => "11001001",26779 => "01011001",26780 => "10110100",26781 => "01011000",26782 => "10000101",26783 => "00000010",26784 => "10010010",26785 => "01101110",26786 => "01011010",26787 => "11100011",26788 => "01001001",26789 => "11111110",26790 => "00001001",26791 => "11011110",26792 => "11000001",26793 => "10001000",26794 => "01000111",26795 => "10000101",26796 => "01001100",26797 => "11011100",26798 => "10000101",26799 => "01000101",26800 => "01110111",26801 => "00110010",26802 => "10010011",26803 => "00000011",26804 => "11101111",26805 => "01101010",26806 => "01101001",26807 => "11111111",26808 => "00101000",26809 => "00000011",26810 => "10010001",26811 => "10001110",26812 => "01110010",26813 => "01010000",26814 => "10110100",26815 => "01101101",26816 => "10110110",26817 => "10011111",26818 => "00100001",26819 => "10010101",26820 => "01000001",26821 => "10001000",26822 => "00101110",26823 => "10001000",26824 => "10011101",26825 => "10100111",26826 => "10111100",26827 => "10101011",26828 => "01111010",26829 => "10000100",26830 => "01010111",26831 => "10110111",26832 => "01011101",26833 => "10101010",26834 => "11101010",26835 => "01011011",26836 => "01000011",26837 => "01000000",26838 => "00000110",26839 => "01000101",26840 => "11100010",26841 => "00111100",26842 => "01000000",26843 => "11001001",26844 => "01100010",26845 => "10110000",26846 => "10101011",26847 => "01001011",26848 => "11100100",26849 => "10010111",26850 => "01001000",26851 => "10111011",26852 => "11001011",26853 => "01000000",26854 => "10111011",26855 => "11011100",26856 => "10111110",26857 => "10010111",26858 => "00000000",26859 => "11101010",26860 => "10110000",26861 => "10000111",26862 => "10011110",26863 => "11101000",26864 => "10111111",26865 => "11111110",26866 => "11111111",26867 => "00000010",26868 => "11010010",26869 => "00110111",26870 => "01000000",26871 => "11001010",26872 => "00111100",26873 => "01110001",26874 => "11110110",26875 => "00100000",26876 => "01110100",26877 => "11111101",26878 => "01010101",26879 => "01010101",26880 => "11000011",26881 => "10011010",26882 => "00000100",26883 => "11101011",26884 => "01111110",26885 => "00001010",26886 => "11110101",26887 => "11011010",26888 => "00111010",26889 => "10101000",26890 => "00001000",26891 => "10100110",26892 => "01001001",26893 => "01001111",26894 => "01111000",26895 => "11011010",26896 => "10110011",26897 => "10011110",26898 => "10101011",26899 => "10100100",26900 => "11100101",26901 => "00110100",26902 => "10001010",26903 => "11110111",26904 => "11101010",26905 => "10010110",26906 => "00011001",26907 => "11000101",26908 => "10101001",26909 => "10100000",26910 => "01101001",26911 => "00001000",26912 => "01001001",26913 => "01110111",26914 => "10010110",26915 => "01001100",26916 => "11000110",26917 => "10101000",26918 => "10001001",26919 => "10100001",26920 => "10101000",26921 => "11000111",26922 => "10100100",26923 => "10010111",26924 => "00100111",26925 => "11111111",26926 => "01110100",26927 => "10010011",26928 => "01010101",26929 => "01010010",26930 => "10100011",26931 => "10111010",26932 => "00111011",26933 => "11100110",26934 => "00011010",26935 => "01111000",26936 => "11001110",26937 => "01100001",26938 => "00001111",26939 => "10000111",26940 => "01010001",26941 => "00101110",26942 => "01100111",26943 => "00110110",26944 => "11011110",26945 => "11010010",26946 => "01101001",26947 => "11011110",26948 => "00001011",26949 => "01011011",26950 => "00001000",26951 => "01011101",26952 => "10011101",26953 => "00101111",26954 => "11101111",26955 => "10111111",26956 => "10011110",26957 => "10011000",26958 => "11100110",26959 => "01111101",26960 => "10000000",26961 => "00110000",26962 => "11101000",26963 => "00000010",26964 => "00010001",26965 => "01110101",26966 => "10110110",26967 => "00011010",26968 => "11000100",26969 => "01000110",26970 => "11100100",26971 => "10101110",26972 => "01110110",26973 => "00101111",26974 => "11011110",26975 => "10000101",26976 => "01110111",26977 => "10101110",26978 => "10010000",26979 => "01011110",26980 => "11000011",26981 => "10101010",26982 => "01110111",26983 => "11101111",26984 => "10111111",26985 => "01100110",26986 => "10100101",26987 => "10011110",26988 => "11001101",26989 => "10101110",26990 => "10001011",26991 => "11010100",26992 => "10110011",26993 => "11011111",26994 => "01010010",26995 => "00011111",26996 => "01010100",26997 => "10101001",26998 => "11000110",26999 => "00111110",27000 => "01100111",27001 => "10011010",27002 => "10101110",27003 => "00100100",27004 => "01100010",27005 => "10100111",27006 => "01110101",27007 => "10110011",27008 => "10011011",27009 => "11100101",27010 => "11111110",27011 => "00010110",27012 => "11101011",27013 => "10000100",27014 => "10100110",27015 => "10100111",27016 => "10010000",27017 => "10010101",27018 => "00101110",27019 => "11100011",27020 => "11101011",27021 => "01101010",27022 => "10111001",27023 => "01111011",27024 => "10011100",27025 => "11000011",27026 => "10010101",27027 => "11000111",27028 => "01000000",27029 => "01010111",27030 => "01101110",27031 => "00100100",27032 => "00001100",27033 => "11001011",27034 => "11011001",27035 => "10001101",27036 => "00110110",27037 => "00111011",27038 => "10010100",27039 => "11100011",27040 => "11101011",27041 => "10111011",27042 => "10100111",27043 => "00110000",27044 => "01111110",27045 => "01000010",27046 => "00110111",27047 => "00101101",27048 => "01110111",27049 => "10110111",27050 => "00111110",27051 => "11000000",27052 => "00001100",27053 => "00101010",27054 => "00101010",27055 => "01001001",27056 => "10010001",27057 => "01001101",27058 => "01000000",27059 => "00000010",27060 => "01110001",27061 => "00010101",27062 => "11111001",27063 => "10111101",27064 => "10001010",27065 => "10010001",27066 => "01011001",27067 => "01011100",27068 => "11110001",27069 => "10011101",27070 => "01110011",27071 => "01110011",27072 => "11001011",27073 => "11010010",27074 => "01110011",27075 => "01011010",27076 => "10011010",27077 => "10010110",27078 => "00110101",27079 => "00001110",27080 => "10101010",27081 => "01100111",27082 => "10110111",27083 => "00110000",27084 => "10011101",27085 => "10000000",27086 => "00011000",27087 => "11100000",27088 => "11110011",27089 => "00001001",27090 => "10100100",27091 => "10110010",27092 => "10000011",27093 => "00010000",27094 => "10100111",27095 => "00101110",27096 => "11010010",27097 => "01000110",27098 => "01100101",27099 => "01000010",27100 => "00100111",27101 => "01010010",27102 => "00100010",27103 => "10001010",27104 => "00101000",27105 => "01110000",27106 => "00010110",27107 => "11010001",27108 => "11000011",27109 => "00101000",27110 => "10110011",27111 => "01001100",27112 => "00001000",27113 => "01000111",27114 => "01101100",27115 => "00110011",27116 => "01111110",27117 => "00000011",27118 => "10001100",27119 => "00011111",27120 => "11011110",27121 => "10100010",27122 => "01110100",27123 => "01111100",27124 => "01000111",27125 => "10000000",27126 => "11011011",27127 => "00111110",27128 => "00010110",27129 => "00100011",27130 => "00011011",27131 => "00000011",27132 => "00000010",27133 => "11100001",27134 => "01111001",27135 => "11010010",27136 => "01010111",27137 => "10000100",27138 => "10010110",27139 => "11101110",27140 => "10011110",27141 => "01110001",27142 => "10011010",27143 => "10100100",27144 => "10000110",27145 => "10001101",27146 => "00101010",27147 => "10011000",27148 => "00011110",27149 => "00001111",27150 => "01101010",27151 => "11011101",27152 => "00011001",27153 => "01111110",27154 => "00001001",27155 => "11011101",27156 => "11110111",27157 => "11111000",27158 => "11010010",27159 => "11010100",27160 => "11001101",27161 => "00111111",27162 => "01010101",27163 => "11000110",27164 => "00010101",27165 => "10000101",27166 => "01010001",27167 => "11000000",27168 => "11011111",27169 => "01010111",27170 => "11010000",27171 => "11011101",27172 => "10111010",27173 => "00111001",27174 => "00000011",27175 => "01001010",27176 => "01001011",27177 => "01011110",27178 => "01001001",27179 => "00010011",27180 => "01110100",27181 => "01101001",27182 => "11111011",27183 => "11010100",27184 => "01111011",27185 => "10101000",27186 => "01000011",27187 => "10111110",27188 => "00010010",27189 => "10011000",27190 => "10001101",27191 => "01101101",27192 => "01010110",27193 => "11101000",27194 => "00100001",27195 => "01101001",27196 => "10010000",27197 => "11101000",27198 => "11111100",27199 => "00010110",27200 => "11011110",27201 => "00110110",27202 => "00011101",27203 => "01011010",27204 => "00100110",27205 => "11010111",27206 => "11000011",27207 => "01101111",27208 => "00010111",27209 => "01100111",27210 => "11001110",27211 => "00010111",27212 => "11111110",27213 => "00011010",27214 => "00010111",27215 => "00110101",27216 => "01111010",27217 => "01101010",27218 => "11111101",27219 => "11010111",27220 => "11100001",27221 => "10101011",27222 => "11101001",27223 => "00110000",27224 => "11111011",27225 => "10111100",27226 => "00111001",27227 => "11110101",27228 => "11010000",27229 => "01010001",27230 => "01001100",27231 => "00000001",27232 => "01100011",27233 => "01101000",27234 => "11101001",27235 => "11100000",27236 => "11100011",27237 => "00001101",27238 => "00011110",27239 => "10011111",27240 => "01101001",27241 => "01000011",27242 => "00111000",27243 => "10000010",27244 => "10101010",27245 => "00000001",27246 => "10111101",27247 => "00010001",27248 => "10101010",27249 => "11101100",27250 => "01111010",27251 => "10011100",27252 => "01011100",27253 => "10001110",27254 => "01111100",27255 => "01010010",27256 => "11011111",27257 => "10101111",27258 => "00010100",27259 => "10111000",27260 => "00000101",27261 => "01010111",27262 => "11011100",27263 => "00110001",27264 => "11001011",27265 => "00101001",27266 => "00000001",27267 => "10000011",27268 => "00011111",27269 => "10111111",27270 => "11000000",27271 => "10000010",27272 => "01000110",27273 => "11001100",27274 => "11010111",27275 => "00010000",27276 => "11010011",27277 => "11110110",27278 => "10011001",27279 => "11111001",27280 => "11011110",27281 => "01011001",27282 => "01010111",27283 => "10110110",27284 => "01101100",27285 => "10110100",27286 => "00110010",27287 => "00111100",27288 => "10010110",27289 => "11111111",27290 => "11110100",27291 => "00000101",27292 => "01001100",27293 => "10010000",27294 => "10110111",27295 => "00010000",27296 => "10101000",27297 => "11011010",27298 => "01111110",27299 => "00000101",27300 => "01110101",27301 => "10011001",27302 => "10011010",27303 => "01110011",27304 => "11100111",27305 => "11101001",27306 => "10010011",27307 => "01010001",27308 => "11111111",27309 => "10110011",27310 => "10100111",27311 => "11001110",27312 => "10110111",27313 => "01000010",27314 => "00011010",27315 => "10001101",27316 => "10110110",27317 => "11000001",27318 => "01101010",27319 => "00100110",27320 => "11111000",27321 => "00010100",27322 => "01101010",27323 => "10010100",27324 => "00011101",27325 => "00000111",27326 => "10011100",27327 => "00100100",27328 => "01100110",27329 => "01011110",27330 => "10100001",27331 => "01011110",27332 => "01010001",27333 => "10111001",27334 => "00100101",27335 => "10011000",27336 => "10000110",27337 => "00100111",27338 => "11100111",27339 => "11010000",27340 => "11100010",27341 => "01110111",27342 => "01101010",27343 => "11101011",27344 => "11000011",27345 => "11100101",27346 => "11001101",27347 => "00100110",27348 => "00000010",27349 => "01001101",27350 => "11110110",27351 => "10011000",27352 => "11010001",27353 => "00011100",27354 => "10001111",27355 => "00001011",27356 => "00111011",27357 => "01111111",27358 => "00101101",27359 => "00110010",27360 => "01001000",27361 => "10000100",27362 => "00011111",27363 => "01101100",27364 => "11010110",27365 => "10111100",27366 => "00000100",27367 => "00001101",27368 => "11001011",27369 => "10010101",27370 => "10000011",27371 => "10101101",27372 => "01111111",27373 => "10101100",27374 => "11110001",27375 => "11100111",27376 => "00011111",27377 => "11011000",27378 => "10110001",27379 => "00001101",27380 => "10100100",27381 => "11000000",27382 => "10011001",27383 => "11110101",27384 => "01111001",27385 => "00010000",27386 => "00110001",27387 => "01010110",27388 => "10110010",27389 => "00100101",27390 => "11101110",27391 => "01101110",27392 => "00110000",27393 => "01011110",27394 => "11011100",27395 => "01110100",27396 => "10001110",27397 => "01110101",27398 => "10100100",27399 => "10101010",27400 => "01110011",27401 => "00101010",27402 => "01111101",27403 => "00100011",27404 => "10001000",27405 => "10010101",27406 => "01111110",27407 => "10001100",27408 => "01001110",27409 => "11011100",27410 => "10010010",27411 => "00110110",27412 => "10011010",27413 => "00110010",27414 => "11001011",27415 => "11000011",27416 => "11111111",27417 => "10010001",27418 => "01111111",27419 => "11011100",27420 => "01010100",27421 => "00011110",27422 => "11010000",27423 => "10001101",27424 => "10111001",27425 => "10001010",27426 => "10010110",27427 => "00010010",27428 => "11011010",27429 => "00110110",27430 => "11110101",27431 => "00000011",27432 => "01000111",27433 => "11111111",27434 => "11001101",27435 => "10100010",27436 => "11100101",27437 => "11110101",27438 => "10001110",27439 => "10101110",27440 => "00100001",27441 => "00110111",27442 => "00010100",27443 => "11000101",27444 => "00100111",27445 => "10100001",27446 => "01000001",27447 => "10000001",27448 => "00111101",27449 => "10000011",27450 => "01101001",27451 => "10001110",27452 => "10000111",27453 => "11000000",27454 => "00111000",27455 => "10111110",27456 => "10001110",27457 => "00111010",27458 => "10101010",27459 => "01000110",27460 => "01001111",27461 => "10100011",27462 => "01011100",27463 => "10000011",27464 => "10011100",27465 => "00101110",27466 => "00000001",27467 => "10000111",27468 => "10001010",27469 => "01101100",27470 => "01001111",27471 => "00011101",27472 => "10110001",27473 => "00011011",27474 => "01010010",27475 => "10101000",27476 => "01100001",27477 => "00111110",27478 => "01110001",27479 => "01110111",27480 => "11101000",27481 => "00100111",27482 => "00101001",27483 => "10000100",27484 => "10110100",27485 => "00010010",27486 => "00011110",27487 => "01101000",27488 => "10100011",27489 => "11101000",27490 => "10110111",27491 => "11010010",27492 => "00011000",27493 => "10011000",27494 => "01001011",27495 => "01000010",27496 => "10011000",27497 => "01100011",27498 => "01101100",27499 => "00111010",27500 => "10001001",27501 => "10111110",27502 => "01110011",27503 => "01110010",27504 => "10011001",27505 => "00001011",27506 => "01000011",27507 => "10010000",27508 => "11101010",27509 => "10110110",27510 => "00011101",27511 => "11000011",27512 => "10011110",27513 => "01011011",27514 => "00000000",27515 => "01101100",27516 => "00111111",27517 => "01111100",27518 => "01101110",27519 => "00101011",27520 => "11110000",27521 => "00101111",27522 => "10010111",27523 => "11001110",27524 => "01001111",27525 => "00010100",27526 => "00101011",27527 => "00100011",27528 => "00100001",27529 => "01111001",27530 => "01001100",27531 => "01011110",27532 => "01011111",27533 => "10110011",27534 => "00111111",27535 => "01110110",27536 => "10000101",27537 => "00110000",27538 => "00100011",27539 => "10110100",27540 => "11010000",27541 => "10110100",27542 => "00010101",27543 => "01001011",27544 => "01010010",27545 => "01111001",27546 => "01110111",27547 => "11011111",27548 => "01111110",27549 => "01010111",27550 => "00111101",27551 => "11100001",27552 => "10100011",27553 => "11010011",27554 => "11110101",27555 => "10110001",27556 => "01110100",27557 => "10100110",27558 => "10001110",27559 => "01000101",27560 => "10000000",27561 => "00111001",27562 => "10110111",27563 => "11100000",27564 => "10111001",27565 => "00001100",27566 => "11100101",27567 => "11011111",27568 => "11111101",27569 => "00010000",27570 => "01111011",27571 => "11101000",27572 => "01101100",27573 => "11011111",27574 => "11000111",27575 => "10001011",27576 => "11000111",27577 => "11101101",27578 => "11101011",27579 => "01001000",27580 => "11000000",27581 => "00101100",27582 => "11100101",27583 => "00010110",27584 => "01000011",27585 => "00010001",27586 => "00110111",27587 => "10111011",27588 => "10011011",27589 => "01110110",27590 => "00110001",27591 => "10010001",27592 => "00011000",27593 => "01101011",27594 => "00110010",27595 => "11101001",27596 => "11101011",27597 => "01111011",27598 => "10110111",27599 => "01110111",27600 => "11000011",27601 => "01101000",27602 => "00101000",27603 => "11000110",27604 => "01001001",27605 => "01110000",27606 => "01010011",27607 => "10010111",27608 => "10011110",27609 => "10011011",27610 => "11111111",27611 => "10101011",27612 => "00110101",27613 => "11101011",27614 => "11110010",27615 => "00001001",27616 => "11110010",27617 => "01000110",27618 => "10101000",27619 => "10100111",27620 => "00110011",27621 => "01111010",27622 => "01100101",27623 => "00001000",27624 => "10001110",27625 => "00010010",27626 => "00000011",27627 => "00011010",27628 => "01111110",27629 => "01001000",27630 => "01101010",27631 => "10111101",27632 => "01110100",27633 => "11100001",27634 => "11111100",27635 => "01111100",27636 => "10111110",27637 => "01000010",27638 => "01010000",27639 => "11011001",27640 => "01101010",27641 => "10111101",27642 => "11101101",27643 => "00000110",27644 => "10001010",27645 => "00100011",27646 => "00000010",27647 => "01100111",27648 => "10111110",27649 => "01011111",27650 => "10011000",27651 => "11000001",27652 => "11110111",27653 => "10110100",27654 => "10000001",27655 => "01000100",27656 => "11010101",27657 => "00010101",27658 => "00101100",27659 => "01010011",27660 => "00100011",27661 => "11000111",27662 => "00000010",27663 => "11111001",27664 => "10111101",27665 => "00111111",27666 => "00110100",27667 => "00010111",27668 => "10100111",27669 => "01101110",27670 => "01001000",27671 => "00110000",27672 => "01110001",27673 => "00001110",27674 => "11010001",27675 => "00011111",27676 => "11000011",27677 => "11101110",27678 => "01100011",27679 => "11010100",27680 => "01101010",27681 => "00001111",27682 => "10111100",27683 => "11011011",27684 => "11110001",27685 => "10101001",27686 => "10011000",27687 => "11011101",27688 => "11001100",27689 => "11111000",27690 => "11111110",27691 => "01011100",27692 => "00001000",27693 => "00000010",27694 => "01000110",27695 => "11001111",27696 => "10000000",27697 => "01010001",27698 => "00110110",27699 => "11110101",27700 => "11100010",27701 => "00100101",27702 => "00001101",27703 => "00011110",27704 => "00100001",27705 => "00011000",27706 => "11011010",27707 => "11010000",27708 => "01011100",27709 => "10111100",27710 => "01110010",27711 => "10001101",27712 => "10010110",27713 => "00101101",27714 => "00011010",27715 => "10100100",27716 => "01101000",27717 => "11011101",27718 => "11111110",27719 => "11001001",27720 => "11111010",27721 => "01001100",27722 => "01100010",27723 => "10110110",27724 => "10000101",27725 => "01101101",27726 => "11100001",27727 => "01101000",27728 => "01101011",27729 => "01101100",27730 => "11000111",27731 => "10011000",27732 => "11001110",27733 => "00011101",27734 => "11000100",27735 => "10010010",27736 => "00001101",27737 => "10010001",27738 => "10110001",27739 => "01011001",27740 => "10111110",27741 => "11100000",27742 => "00011110",27743 => "10101100",27744 => "10101110",27745 => "10010100",27746 => "10100001",27747 => "10101011",27748 => "00001000",27749 => "00111010",27750 => "10101000",27751 => "00101100",27752 => "01010111",27753 => "10100001",27754 => "01101001",27755 => "11110011",27756 => "10111001",27757 => "00010001",27758 => "10101000",27759 => "01011101",27760 => "11001111",27761 => "01100011",27762 => "10111011",27763 => "11101001",27764 => "00110000",27765 => "01110000",27766 => "10000101",27767 => "01001010",27768 => "11101010",27769 => "01101000",27770 => "10110000",27771 => "01101101",27772 => "11010000",27773 => "00000110",27774 => "00001101",27775 => "10110100",27776 => "01101110",27777 => "00111000",27778 => "11111111",27779 => "01011000",27780 => "10111101",27781 => "11110011",27782 => "01010101",27783 => "01010010",27784 => "10111001",27785 => "01010000",27786 => "01110001",27787 => "11111111",27788 => "10111111",27789 => "01111111",27790 => "10000111",27791 => "01001110",27792 => "01011000",27793 => "10100101",27794 => "00100111",27795 => "11001110",27796 => "00101101",27797 => "10010111",27798 => "11011000",27799 => "00001000",27800 => "10010111",27801 => "00110110",27802 => "00010001",27803 => "00110001",27804 => "10110110",27805 => "01101111",27806 => "10010000",27807 => "11111000",27808 => "10011110",27809 => "00100110",27810 => "00000010",27811 => "10001111",27812 => "01011101",27813 => "10101101",27814 => "01100010",27815 => "00101111",27816 => "00111100",27817 => "10001001",27818 => "10101011",27819 => "01011001",27820 => "00111001",27821 => "01010100",27822 => "01010001",27823 => "10100110",27824 => "10000011",27825 => "00010110",27826 => "11101000",27827 => "10011001",27828 => "00101000",27829 => "01011010",27830 => "00111100",27831 => "11010010",27832 => "00010001",27833 => "10011100",27834 => "00000001",27835 => "01111001",27836 => "11011001",27837 => "01000001",27838 => "01111100",27839 => "11101001",27840 => "00100001",27841 => "10101000",27842 => "11000101",27843 => "01111111",27844 => "11001011",27845 => "01000001",27846 => "11001011",27847 => "10001001",27848 => "01000000",27849 => "11111100",27850 => "00101010",27851 => "10000000",27852 => "11010010",27853 => "00011110",27854 => "10100101",27855 => "10100100",27856 => "11110111",27857 => "00110110",27858 => "00100000",27859 => "10011010",27860 => "01000110",27861 => "10111101",27862 => "10100101",27863 => "01100001",27864 => "10111110",27865 => "01101111",27866 => "11011000",27867 => "01010010",27868 => "11010111",27869 => "00111000",27870 => "00010010",27871 => "01011100",27872 => "10010000",27873 => "11010001",27874 => "10110001",27875 => "01100001",27876 => "01110101",27877 => "11011110",27878 => "11100101",27879 => "11110110",27880 => "10010010",27881 => "10101001",27882 => "00100111",27883 => "01110011",27884 => "10011010",27885 => "10011001",27886 => "01111000",27887 => "11111011",27888 => "00110011",27889 => "10000000",27890 => "11010011",27891 => "10000101",27892 => "11001101",27893 => "00110100",27894 => "11001001",27895 => "10100000",27896 => "10101111",27897 => "10101000",27898 => "01111110",27899 => "01010001",27900 => "00101110",27901 => "00011101",27902 => "11011101",27903 => "01110000",27904 => "00100000",27905 => "11010011",27906 => "11100111",27907 => "11101100",27908 => "00111011",27909 => "00110110",27910 => "10101100",27911 => "00001111",27912 => "01111000",27913 => "00101111",27914 => "01010110",27915 => "00001111",27916 => "10000011",27917 => "11000111",27918 => "00100100",27919 => "11101111",27920 => "10100010",27921 => "00111101",27922 => "00101001",27923 => "01100101",27924 => "11110011",27925 => "10111110",27926 => "10011110",27927 => "11110101",27928 => "10110010",27929 => "10010111",27930 => "11111011",27931 => "01000110",27932 => "11110101",27933 => "10101101",27934 => "00001011",27935 => "10011111",27936 => "00101000",27937 => "11010101",27938 => "00100010",27939 => "00110001",27940 => "11101100",27941 => "00100011",27942 => "01000000",27943 => "11100111",27944 => "11010010",27945 => "01100001",27946 => "11000111",27947 => "11101111",27948 => "00000100",27949 => "01010110",27950 => "11010000",27951 => "11000101",27952 => "01100101",27953 => "11111000",27954 => "00101101",27955 => "00110010",27956 => "11101000",27957 => "00010111",27958 => "10001011",27959 => "01100110",27960 => "11001111",27961 => "10000110",27962 => "11000001",27963 => "00001001",27964 => "11001011",27965 => "10000110",27966 => "11001001",27967 => "01111001",27968 => "00001001",27969 => "00111011",27970 => "01001111",27971 => "00010101",27972 => "01000011",27973 => "11011001",27974 => "10100101",27975 => "00101000",27976 => "00101101",27977 => "00100101",27978 => "10111100",27979 => "10001110",27980 => "00000000",27981 => "10110000",27982 => "00011101",27983 => "00010010",27984 => "01111100",27985 => "10101111",27986 => "11100110",27987 => "01111010",27988 => "01111010",27989 => "11001000",27990 => "10101001",27991 => "00011010",27992 => "11101000",27993 => "10000111",27994 => "01100111",27995 => "10001111",27996 => "01111000",27997 => "00110100",27998 => "11101110",27999 => "10110010",28000 => "00110010",28001 => "10111000",28002 => "10001100",28003 => "00000000",28004 => "01001101",28005 => "11100101",28006 => "11110001",28007 => "01101000",28008 => "00011000",28009 => "00111111",28010 => "01011101",28011 => "01111000",28012 => "01001010",28013 => "00110000",28014 => "00100101",28015 => "11111100",28016 => "00010010",28017 => "00000010",28018 => "00101001",28019 => "00110100",28020 => "10111001",28021 => "11011101",28022 => "01110000",28023 => "11000111",28024 => "11100110",28025 => "10011001",28026 => "01011111",28027 => "01111111",28028 => "01001000",28029 => "00010111",28030 => "00011101",28031 => "00010101",28032 => "11001010",28033 => "10011010",28034 => "11011111",28035 => "11000100",28036 => "11001000",28037 => "10001111",28038 => "10010011",28039 => "11101101",28040 => "11101101",28041 => "10011011",28042 => "11011110",28043 => "00101001",28044 => "10101001",28045 => "11110000",28046 => "01000110",28047 => "10001010",28048 => "11111011",28049 => "10101011",28050 => "10110001",28051 => "00110010",28052 => "00111000",28053 => "10111101",28054 => "11100001",28055 => "11100101",28056 => "10110011",28057 => "11111010",28058 => "01111011",28059 => "01101111",28060 => "11100011",28061 => "10001011",28062 => "11100001",28063 => "11111010",28064 => "10010000",28065 => "01100110",28066 => "00010100",28067 => "01101110",28068 => "10000001",28069 => "01110000",28070 => "11101001",28071 => "00010011",28072 => "10011101",28073 => "01100001",28074 => "10110110",28075 => "11010101",28076 => "10001101",28077 => "11111001",28078 => "10001101",28079 => "01111010",28080 => "00111011",28081 => "01100110",28082 => "10011110",28083 => "11010101",28084 => "01011010",28085 => "11100010",28086 => "01101111",28087 => "10110111",28088 => "01000010",28089 => "10001110",28090 => "00001100",28091 => "01001111",28092 => "10011010",28093 => "01011001",28094 => "10001100",28095 => "10010111",28096 => "10001011",28097 => "01101100",28098 => "11110110",28099 => "01010011",28100 => "01110111",28101 => "10010000",28102 => "10101100",28103 => "00111101",28104 => "11011011",28105 => "01010111",28106 => "01001101",28107 => "11011110",28108 => "01000110",28109 => "10110111",28110 => "11010110",28111 => "11110110",28112 => "01000010",28113 => "11110100",28114 => "10101101",28115 => "01111110",28116 => "11100001",28117 => "11010100",28118 => "00100000",28119 => "01000110",28120 => "11100010",28121 => "11010111",28122 => "11001110",28123 => "11011001",28124 => "11110001",28125 => "10000011",28126 => "11000010",28127 => "11100100",28128 => "11101111",28129 => "01111000",28130 => "11101011",28131 => "01000000",28132 => "00001110",28133 => "00111010",28134 => "00111110",28135 => "01111100",28136 => "01100110",28137 => "10001010",28138 => "00000011",28139 => "11100000",28140 => "00101001",28141 => "01101011",28142 => "00101100",28143 => "11001110",28144 => "11111100",28145 => "01011000",28146 => "01010100",28147 => "01010111",28148 => "01100111",28149 => "10001110",28150 => "10101001",28151 => "10101011",28152 => "11111110",28153 => "10000111",28154 => "11001010",28155 => "11110110",28156 => "11111111",28157 => "10010110",28158 => "00110101",28159 => "10000011",28160 => "00101111",28161 => "10000010",28162 => "10100111",28163 => "10111010",28164 => "01010111",28165 => "10111011",28166 => "00000010",28167 => "01111110",28168 => "11111101",28169 => "11111110",28170 => "10101101",28171 => "00111111",28172 => "00011001",28173 => "01010100",28174 => "01100010",28175 => "00101100",28176 => "10011100",28177 => "11101001",28178 => "01101000",28179 => "01110101",28180 => "00011111",28181 => "01100010",28182 => "11110100",28183 => "00011001",28184 => "10001100",28185 => "11010111",28186 => "00101001",28187 => "00111001",28188 => "11000010",28189 => "11101101",28190 => "11100101",28191 => "11001010",28192 => "10010010",28193 => "01110010",28194 => "01011010",28195 => "10111111",28196 => "10111010",28197 => "10011100",28198 => "01000001",28199 => "01101000",28200 => "01101011",28201 => "00101111",28202 => "11110100",28203 => "01111011",28204 => "00000101",28205 => "00100110",28206 => "00101001",28207 => "00111110",28208 => "11100100",28209 => "11010100",28210 => "10001110",28211 => "00011000",28212 => "01111111",28213 => "10001111",28214 => "10111010",28215 => "11101101",28216 => "11101001",28217 => "11010100",28218 => "10000111",28219 => "00111111",28220 => "11000101",28221 => "10000100",28222 => "10101010",28223 => "10011101",28224 => "10110011",28225 => "00001110",28226 => "11010101",28227 => "10100101",28228 => "11010111",28229 => "11101010",28230 => "10000111",28231 => "11111011",28232 => "01110110",28233 => "10000110",28234 => "11100000",28235 => "11001110",28236 => "11000100",28237 => "01010010",28238 => "11100000",28239 => "11011001",28240 => "11001000",28241 => "01101000",28242 => "10001000",28243 => "10010111",28244 => "00010101",28245 => "01010110",28246 => "11000001",28247 => "00100000",28248 => "00010011",28249 => "10011001",28250 => "01101101",28251 => "01111100",28252 => "00010100",28253 => "10011110",28254 => "10011101",28255 => "11101011",28256 => "00100010",28257 => "01111110",28258 => "10010010",28259 => "10111011",28260 => "10000101",28261 => "00000100",28262 => "10111000",28263 => "10010010",28264 => "11000101",28265 => "00001011",28266 => "10111111",28267 => "10111101",28268 => "00100011",28269 => "11111011",28270 => "00010101",28271 => "11011110",28272 => "00110010",28273 => "00001100",28274 => "11111110",28275 => "10110101",28276 => "10001010",28277 => "01101110",28278 => "01011101",28279 => "00100100",28280 => "00000000",28281 => "00110000",28282 => "11011011",28283 => "00101110",28284 => "00000000",28285 => "01111100",28286 => "00100000",28287 => "11000011",28288 => "11111110",28289 => "01101101",28290 => "10001111",28291 => "11110011",28292 => "00010100",28293 => "00110011",28294 => "10111001",28295 => "01111000",28296 => "00010100",28297 => "11101100",28298 => "01001001",28299 => "01101100",28300 => "01111011",28301 => "10000100",28302 => "10111001",28303 => "01111101",28304 => "10101010",28305 => "11110100",28306 => "01101100",28307 => "01111000",28308 => "11101100",28309 => "01110000",28310 => "11001010",28311 => "11111011",28312 => "01100100",28313 => "11000011",28314 => "11111000",28315 => "00111010",28316 => "00100001",28317 => "00110010",28318 => "01011111",28319 => "00001101",28320 => "00100100",28321 => "01001101",28322 => "11010000",28323 => "00111111",28324 => "01011000",28325 => "01110100",28326 => "01101110",28327 => "01000101",28328 => "11000000",28329 => "11100100",28330 => "10000101",28331 => "00010101",28332 => "00010011",28333 => "00001101",28334 => "11001111",28335 => "10001101",28336 => "11010110",28337 => "01110000",28338 => "10101011",28339 => "01100010",28340 => "00000111",28341 => "01000010",28342 => "10001001",28343 => "01010100",28344 => "01100001",28345 => "01001111",28346 => "11001111",28347 => "00101000",28348 => "01000011",28349 => "00010001",28350 => "00101111",28351 => "00100011",28352 => "11001011",28353 => "10100011",28354 => "01001000",28355 => "01101000",28356 => "10101001",28357 => "11001010",28358 => "10110101",28359 => "10101011",28360 => "00010101",28361 => "00000001",28362 => "00010001",28363 => "00011010",28364 => "00001101",28365 => "11010110",28366 => "11011001",28367 => "00101011",28368 => "11110001",28369 => "11111111",28370 => "01100100",28371 => "01000110",28372 => "10100000",28373 => "11110010",28374 => "11101010",28375 => "00000101",28376 => "01010100",28377 => "00100100",28378 => "10011111",28379 => "11111010",28380 => "00110010",28381 => "11010001",28382 => "10010011",28383 => "11000110",28384 => "10011001",28385 => "01001010",28386 => "10110010",28387 => "00100011",28388 => "11110001",28389 => "00010011",28390 => "00110101",28391 => "11111011",28392 => "00010101",28393 => "10110101",28394 => "10000110",28395 => "11100101",28396 => "01110110",28397 => "00101100",28398 => "11101000",28399 => "10111110",28400 => "11110100",28401 => "10001110",28402 => "00000010",28403 => "00111101",28404 => "11011101",28405 => "01111000",28406 => "11101000",28407 => "10011011",28408 => "10100001",28409 => "01011011",28410 => "10100011",28411 => "10010110",28412 => "11100001",28413 => "00100011",28414 => "10110111",28415 => "01110100",28416 => "10111000",28417 => "10101111",28418 => "10000101",28419 => "01010010",28420 => "11110111",28421 => "01111110",28422 => "10110010",28423 => "10101100",28424 => "00011111",28425 => "10100000",28426 => "11010100",28427 => "01110001",28428 => "00010111",28429 => "01011111",28430 => "00111101",28431 => "01000000",28432 => "10010101",28433 => "10100010",28434 => "01010101",28435 => "10001010",28436 => "11011100",28437 => "10111101",28438 => "00101001",28439 => "01010001",28440 => "00111111",28441 => "00100010",28442 => "11011001",28443 => "01100010",28444 => "00011110",28445 => "00100011",28446 => "01001010",28447 => "00010111",28448 => "01011000",28449 => "10001000",28450 => "10101110",28451 => "11010110",28452 => "00100001",28453 => "11001001",28454 => "00001010",28455 => "10100100",28456 => "11110001",28457 => "11010001",28458 => "10000011",28459 => "00110101",28460 => "10011011",28461 => "10011011",28462 => "10001010",28463 => "01010001",28464 => "00111100",28465 => "01001010",28466 => "10110100",28467 => "10010100",28468 => "01001101",28469 => "00011010",28470 => "11110111",28471 => "10011101",28472 => "00001001",28473 => "10011010",28474 => "01111100",28475 => "11010101",28476 => "10010011",28477 => "11111001",28478 => "01000100",28479 => "00100001",28480 => "10001100",28481 => "11001100",28482 => "01111001",28483 => "11000011",28484 => "00000100",28485 => "01111101",28486 => "01101110",28487 => "11000100",28488 => "10101111",28489 => "11011000",28490 => "11100100",28491 => "11100010",28492 => "01010000",28493 => "11101111",28494 => "01110111",28495 => "01100011",28496 => "10011011",28497 => "11100001",28498 => "10001011",28499 => "11000001",28500 => "01010101",28501 => "00100111",28502 => "01010110",28503 => "11111000",28504 => "11111000",28505 => "10101010",28506 => "10000111",28507 => "10110011",28508 => "11111111",28509 => "00001000",28510 => "11110010",28511 => "00111011",28512 => "01010101",28513 => "00111000",28514 => "10111001",28515 => "11100001",28516 => "10111001",28517 => "10010110",28518 => "11101111",28519 => "11010100",28520 => "11001011",28521 => "01100101",28522 => "01000110",28523 => "10000100",28524 => "10110110",28525 => "11010111",28526 => "10111101",28527 => "10010000",28528 => "10101110",28529 => "10110010",28530 => "00101011",28531 => "11000100",28532 => "00000100",28533 => "10000111",28534 => "11001100",28535 => "00011101",28536 => "10001111",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "01101111" report "FAIL high bits" severity failure;
assert RAM(0) = "01111000" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
