 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "01111000",3 => "10000001",4 => "00110110",5 => "00010111",6 => "11010100",7 => "11110000",8 => "00001010",9 => "01011111",10 => "10011001",11 => "00111100",12 => "01011111",13 => "11001000",14 => "10011001",15 => "00100010",16 => "10101011",17 => "01110010",18 => "11011010",19 => "10000111",20 => "10010001",21 => "11011010",22 => "11100010",23 => "01101111",24 => "01000111",25 => "10000000",26 => "10111110",27 => "10011000",28 => "00011000",29 => "00001111",30 => "11001110",31 => "11000110",32 => "11011000",33 => "00111001",34 => "00001000",35 => "00011001",36 => "01000011",37 => "10011100",38 => "01001111",39 => "10111001",40 => "00101100",41 => "00001001",42 => "10110001",43 => "00101001",44 => "11101110",45 => "01000101",46 => "10110010",47 => "01000001",48 => "00011000",49 => "00100111",50 => "00101111",51 => "10011111",52 => "11001001",53 => "01000100",54 => "01100000",55 => "11000111",56 => "01011011",57 => "01010110",58 => "01101111",59 => "01100111",60 => "00010010",61 => "00001000",62 => "00100111",63 => "10000011",64 => "00011110",65 => "10001111",66 => "10110011",67 => "00110000",68 => "01101100",69 => "11010000",70 => "11001011",71 => "11000011",72 => "11011001",73 => "11000110",74 => "01001101",75 => "10000111",76 => "11100010",77 => "11101001",78 => "10000010",79 => "00100110",80 => "00010101",81 => "11011000",82 => "11011110",83 => "01010100",84 => "01100011",85 => "01110111",86 => "01000101",87 => "11100010",88 => "01001010",89 => "10011111",90 => "11000011",91 => "00011001",92 => "11101001",93 => "11101001",94 => "00110010",95 => "01000001",96 => "00010101",97 => "10011110",98 => "01000000",99 => "00000110",100 => "10111001",101 => "10100101",102 => "11101000",103 => "11100010",104 => "01110101",105 => "11011111",106 => "11111001",107 => "10111110",108 => "01011101",109 => "11011110",110 => "11110011",111 => "11000111",112 => "00101101",113 => "01101001",114 => "01001101",115 => "00100001",116 => "10111101",117 => "00011000",118 => "01000101",119 => "01110111",120 => "10100111",121 => "11111100",122 => "00101110",123 => "10011110",124 => "01001101",125 => "01010111",126 => "00111110",127 => "11101111",128 => "00000000",129 => "01100011",130 => "10110000",131 => "00110111",132 => "00101011",133 => "00001010",134 => "11100010",135 => "11111001",136 => "01000001",137 => "00000111",138 => "10011111",139 => "01001010",140 => "10110011",141 => "00110100",142 => "00101011",143 => "11010100",144 => "11010110",145 => "00100110",146 => "01011010",147 => "00000110",148 => "01101011",149 => "11101111",150 => "01101001",151 => "10011100",152 => "10110111",153 => "01110101",154 => "01100010",155 => "11101111",156 => "10100010",157 => "11000110",158 => "01000000",159 => "00110010",160 => "00110111",161 => "01010000",162 => "00000100",163 => "00101100",164 => "10001010",165 => "01110100",166 => "11000101",167 => "01111000",168 => "11001010",169 => "00001111",170 => "00000101",171 => "00111000",172 => "01000101",173 => "00101111",174 => "00010010",175 => "10110000",176 => "11111011",177 => "00101100",178 => "10010000",179 => "10110101",180 => "10100101",181 => "10101111",182 => "00010011",183 => "10100111",184 => "01011011",185 => "10111110",186 => "00000001",187 => "10000101",188 => "10010010",189 => "01100011",190 => "11111011",191 => "11011000",192 => "11010110",193 => "11001001",194 => "10111101",195 => "01110101",196 => "01001100",197 => "00101101",198 => "00011101",199 => "00101101",200 => "11110110",201 => "00101010",202 => "11100001",203 => "11001010",204 => "10111111",205 => "11011000",206 => "10000000",207 => "11110100",208 => "00000111",209 => "11010110",210 => "01101011",211 => "01110011",212 => "10011010",213 => "01111011",214 => "11000100",215 => "10000101",216 => "00101110",217 => "11101100",218 => "10000111",219 => "10001100",220 => "11110100",221 => "01010010",222 => "01110010",223 => "00110001",224 => "01101000",225 => "10001100",226 => "11001111",227 => "11011001",228 => "00001100",229 => "01010111",230 => "00000010",231 => "11001011",232 => "01011111",233 => "01010100",234 => "01100111",235 => "10011011",236 => "01010100",237 => "00000001",238 => "00110011",239 => "10001111",240 => "01111101",241 => "01001011",242 => "10111100",243 => "01011111",244 => "11101011",245 => "11100011",246 => "01000001",247 => "11001001",248 => "00000001",249 => "11010110",250 => "00101100",251 => "00000101",252 => "10010111",253 => "10000110",254 => "11010100",255 => "01100111",256 => "01111010",257 => "01001100",258 => "00110110",259 => "01011000",260 => "00110101",261 => "11001100",262 => "01101101",263 => "00011000",264 => "00010010",265 => "01001000",266 => "11000101",267 => "10001110",268 => "10010100",269 => "00101000",270 => "00100110",271 => "01110110",272 => "11100001",273 => "00000101",274 => "00111110",275 => "01101000",276 => "11111001",277 => "01101000",278 => "01011001",279 => "00111010",280 => "10001011",281 => "00001000",282 => "11110100",283 => "01110000",284 => "00110001",285 => "10101010",286 => "11011100",287 => "01001100",288 => "11101101",289 => "11011001",290 => "00011010",291 => "11000011",292 => "10101101",293 => "00101100",294 => "10000001",295 => "10011000",296 => "10100101",297 => "10100111",298 => "01010000",299 => "01000010",300 => "00110111",301 => "11101111",302 => "10101100",303 => "00110110",304 => "11010111",305 => "11011000",306 => "00100111",307 => "10000101",308 => "00010110",309 => "00010101",310 => "10111110",311 => "11001111",312 => "01111001",313 => "10001011",314 => "01011011",315 => "01111010",316 => "01011010",317 => "10101110",318 => "10001111",319 => "01010001",320 => "10101110",321 => "10101111",322 => "01000001",323 => "00011111",324 => "00000101",325 => "10011100",326 => "11101010",327 => "00111101",328 => "01110110",329 => "01001111",330 => "11011110",331 => "00111011",332 => "01001111",333 => "01100100",334 => "10101011",335 => "10111010",336 => "00111110",337 => "10110010",338 => "01111111",339 => "00101011",340 => "01011011",341 => "11010000",342 => "11100100",343 => "11001101",344 => "01111001",345 => "01100111",346 => "10111101",347 => "01111000",348 => "00111000",349 => "10101011",350 => "10000101",351 => "01111001",352 => "11101010",353 => "11011111",354 => "01100101",355 => "11111101",356 => "00111111",357 => "11001001",358 => "10110101",359 => "01010010",360 => "00000101",361 => "11000100",362 => "01011011",363 => "11010100",364 => "11010100",365 => "10000000",366 => "01000000",367 => "00001001",368 => "10110100",369 => "01000011",370 => "00110001",371 => "10001100",372 => "11101010",373 => "01010111",374 => "10000111",375 => "11001101",376 => "00001010",377 => "01010000",378 => "00000011",379 => "11111101",380 => "11101001",381 => "01101000",382 => "11100001",383 => "01100011",384 => "00110000",385 => "01001110",386 => "01010001",387 => "10110101",388 => "10101110",389 => "00100011",390 => "01110111",391 => "10111111",392 => "10100010",393 => "11011011",394 => "10101010",395 => "11011001",396 => "11101000",397 => "11001001",398 => "00100100",399 => "11111100",400 => "01011101",401 => "00001010",402 => "00001000",403 => "00010011",404 => "00000010",405 => "11000111",406 => "10001000",407 => "00001100",408 => "01101110",409 => "11111001",410 => "11111110",411 => "10110011",412 => "11001011",413 => "01110010",414 => "10000110",415 => "10011011",416 => "01101011",417 => "00011100",418 => "00000111",419 => "10000011",420 => "01110110",421 => "00010011",422 => "00110111",423 => "10010110",424 => "11001000",425 => "10001000",426 => "01100001",427 => "00001110",428 => "00011111",429 => "10001010",430 => "10001100",431 => "10110100",432 => "01001110",433 => "10010101",434 => "01011011",435 => "11001000",436 => "11011001",437 => "11010010",438 => "01001111",439 => "00000111",440 => "00001111",441 => "11010011",442 => "00110001",443 => "00111001",444 => "01110100",445 => "01000100",446 => "10100010",447 => "11101111",448 => "01011110",449 => "10010111",450 => "10001111",451 => "00011000",452 => "00001010",453 => "01000100",454 => "00110001",455 => "10010110",456 => "11110000",457 => "01110001",458 => "00111001",459 => "00111001",460 => "10001101",461 => "00111111",462 => "10000010",463 => "00110111",464 => "00010010",465 => "10011000",466 => "11000100",467 => "10101101",468 => "11110101",469 => "11110100",470 => "11000001",471 => "01111101",472 => "11001111",473 => "11100100",474 => "11111010",475 => "01010001",476 => "01011111",477 => "11100011",478 => "00001111",479 => "10010111",480 => "11110010",481 => "10010001",482 => "10000010",483 => "01000010",484 => "10100011",485 => "10011000",486 => "00001101",487 => "01001111",488 => "00111000",489 => "00001000",490 => "11110100",491 => "00101011",492 => "11101001",493 => "10001010",494 => "11000100",495 => "10001110",496 => "00001001",497 => "01101101",498 => "00011110",499 => "11101101",500 => "11000100",501 => "10100001",502 => "10010100",503 => "10111111",504 => "11101000",505 => "01000001",506 => "10000000",507 => "10010001",508 => "00100110",509 => "10010011",510 => "01110110",511 => "11000100",512 => "00001111",513 => "01001001",514 => "11110101",515 => "11000000",516 => "11100000",517 => "10010000",518 => "10110100",519 => "10101010",520 => "11000000",521 => "10111110",522 => "10111011",523 => "11101010",524 => "01001001",525 => "11101100",526 => "10100011",527 => "11001111",528 => "11011111",529 => "00110100",530 => "10100101",531 => "00011011",532 => "10010100",533 => "00100000",534 => "01000000",535 => "10000111",536 => "11101101",537 => "01110111",538 => "10000100",539 => "00000011",540 => "01001010",541 => "00011001",542 => "01111110",543 => "01110010",544 => "01010100",545 => "00011000",546 => "00111001",547 => "00111111",548 => "11111111",549 => "01001001",550 => "01110011",551 => "11110111",552 => "11111011",553 => "01111100",554 => "11101110",555 => "01100100",556 => "11000010",557 => "01100000",558 => "10011010",559 => "01001010",560 => "11111000",561 => "10011011",562 => "01100011",563 => "11110010",564 => "11110001",565 => "11100000",566 => "10011101",567 => "00010101",568 => "11111000",569 => "00001110",570 => "01111000",571 => "11100110",572 => "01111111",573 => "11110001",574 => "00101001",575 => "00100001",576 => "11001000",577 => "01111001",578 => "10100000",579 => "00000001",580 => "10111001",581 => "01000100",582 => "11000000",583 => "00100000",584 => "00100111",585 => "00101011",586 => "11101100",587 => "00011100",588 => "01000100",589 => "01100011",590 => "00101010",591 => "10001100",592 => "01010000",593 => "01111110",594 => "10100000",595 => "11111010",596 => "11111101",597 => "10101100",598 => "00101101",599 => "01011011",600 => "11000110",601 => "01010001",602 => "00001011",603 => "01001110",604 => "01100000",605 => "10111001",606 => "10110101",607 => "11001111",608 => "00110101",609 => "10010010",610 => "01100010",611 => "11001000",612 => "11110001",613 => "00111101",614 => "10110011",615 => "11001101",616 => "10110111",617 => "11110110",618 => "11111011",619 => "00110101",620 => "00011011",621 => "00000101",622 => "00100001",623 => "01100100",624 => "00100100",625 => "00101100",626 => "00111111",627 => "10101101",628 => "10011011",629 => "00001011",630 => "00010010",631 => "11000001",632 => "00011001",633 => "11010011",634 => "00111101",635 => "00110000",636 => "01010010",637 => "00000011",638 => "01101010",639 => "11011011",640 => "00010011",641 => "00001100",642 => "00011100",643 => "11000000",644 => "10110011",645 => "11000011",646 => "11101010",647 => "01001100",648 => "10000101",649 => "11000111",650 => "01011010",651 => "10001101",652 => "01010100",653 => "01100101",654 => "01101010",655 => "01001111",656 => "11101001",657 => "00100111",658 => "01111001",659 => "01000011",660 => "10011111",661 => "11000111",662 => "01110110",663 => "00010101",664 => "11100110",665 => "10110100",666 => "01110110",667 => "11001110",668 => "01000110",669 => "11000111",670 => "01001100",671 => "11100100",672 => "10111101",673 => "10110010",674 => "01110100",675 => "11110110",676 => "00110001",677 => "01001011",678 => "00101111",679 => "01000101",680 => "10111101",681 => "00110110",682 => "10110101",683 => "00011101",684 => "01000000",685 => "01010000",686 => "10011000",687 => "10101011",688 => "10011100",689 => "10011010",690 => "10111000",691 => "10100011",692 => "00010011",693 => "01101101",694 => "11000000",695 => "11000000",696 => "10110001",697 => "11111101",698 => "11010101",699 => "00111110",700 => "11011010",701 => "11010001",702 => "10100101",703 => "00110011",704 => "11101100",705 => "11010011",706 => "01011001",707 => "10011110",708 => "00011000",709 => "10011010",710 => "00110010",711 => "00000001",712 => "00100000",713 => "11100011",714 => "01001110",715 => "01101101",716 => "10001011",717 => "10110011",718 => "11011110",719 => "11100110",720 => "11110101",721 => "00000000",722 => "10001010",723 => "11000001",724 => "10000010",725 => "01100111",726 => "10110001",727 => "00000101",728 => "00011100",729 => "11010001",730 => "01101011",731 => "11000100",732 => "10001101",733 => "01110111",734 => "01011101",735 => "01000001",736 => "00111000",737 => "11011000",738 => "11110011",739 => "10100111",740 => "00111010",741 => "01110010",742 => "00001110",743 => "00111011",744 => "01101101",745 => "11111011",746 => "10100111",747 => "10101001",748 => "10111100",749 => "10000000",750 => "01110011",751 => "01101100",752 => "00101100",753 => "11100001",754 => "10001001",755 => "10110000",756 => "01101100",757 => "01100010",758 => "10000000",759 => "00011111",760 => "11011010",761 => "11000101",762 => "11010001",763 => "10001001",764 => "10110111",765 => "01001000",766 => "11110100",767 => "11111111",768 => "11000011",769 => "00100110",770 => "10001100",771 => "11111101",772 => "01000011",773 => "10001110",774 => "11001101",775 => "00111010",776 => "10010111",777 => "11111011",778 => "10011100",779 => "01010110",780 => "10101000",781 => "01000101",782 => "10001101",783 => "10010010",784 => "11100010",785 => "10111000",786 => "01000111",787 => "01011100",788 => "01101100",789 => "00100011",790 => "00001100",791 => "11111011",792 => "11000111",793 => "01111100",794 => "01110001",795 => "00001100",796 => "11100001",797 => "01111010",798 => "11111011",799 => "11011110",800 => "00010000",801 => "00011000",802 => "11111001",803 => "01000001",804 => "10010010",805 => "11010000",806 => "00101011",807 => "01101101",808 => "00010111",809 => "11001101",810 => "11100000",811 => "10101101",812 => "01011111",813 => "01011110",814 => "01000001",815 => "00101000",816 => "11000100",817 => "11111001",818 => "00110111",819 => "00100101",820 => "10001100",821 => "00001110",822 => "10011100",823 => "10101111",824 => "00000001",825 => "00111001",826 => "01001001",827 => "01110011",828 => "10001000",829 => "11110000",830 => "10001010",831 => "00010001",832 => "00101001",833 => "00111110",834 => "00101100",835 => "11100111",836 => "11011001",837 => "00100010",838 => "11000010",839 => "01111010",840 => "10100001",841 => "01100011",842 => "11000111",843 => "00011001",844 => "11000101",845 => "00100001",846 => "10010110",847 => "01100000",848 => "00101000",849 => "01111110",850 => "11110101",851 => "01110110",852 => "01101010",853 => "00100111",854 => "11000111",855 => "11000111",856 => "11011111",857 => "00101000",858 => "10000010",859 => "01101011",860 => "11001111",861 => "10001101",862 => "01110101",863 => "00010111",864 => "11101100",865 => "01111011",866 => "01001010",867 => "00110001",868 => "01000100",869 => "11100111",870 => "10011010",871 => "01000111",872 => "00100100",873 => "00100010",874 => "01110000",875 => "01111100",876 => "11101101",877 => "00110010",878 => "10100111",879 => "00101000",880 => "01000010",881 => "00111010",882 => "00000110",883 => "10110011",884 => "00101111",885 => "10101110",886 => "01000001",887 => "00101111",888 => "00011010",889 => "00011001",890 => "10111010",891 => "11001111",892 => "11001001",893 => "11100100",894 => "10110010",895 => "01011011",896 => "01011000",897 => "11000111",898 => "00101001",899 => "11101101",900 => "01011100",901 => "00000111",902 => "10111110",903 => "00111101",904 => "10110101",905 => "11001111",906 => "10010110",907 => "01000111",908 => "01000011",909 => "10010101",910 => "11111111",911 => "00110101",912 => "11111110",913 => "11011100",914 => "00000000",915 => "10001111",916 => "00001001",917 => "00000111",918 => "00100010",919 => "11110111",920 => "01000110",921 => "10110011",922 => "11011100",923 => "11100010",924 => "10000110",925 => "01110000",926 => "01110100",927 => "00101001",928 => "10000011",929 => "11101111",930 => "01000100",931 => "10101010",932 => "01011100",933 => "10110101",934 => "11100101",935 => "01000101",936 => "01110001",937 => "10110110",938 => "10111110",939 => "01100010",940 => "11011100",941 => "10011110",942 => "01011101",943 => "01110010",944 => "10101000",945 => "10111001",946 => "01001011",947 => "10101000",948 => "00001111",949 => "00101011",950 => "11010111",951 => "00001110",952 => "10110101",953 => "11010110",954 => "10101000",955 => "00111111",956 => "01110010",957 => "11010000",958 => "01011111",959 => "11010101",960 => "01011101",961 => "11111011",962 => "11011110",963 => "00110110",964 => "11110110",965 => "00001001",966 => "11101111",967 => "10011000",968 => "01110111",969 => "10001010",970 => "01001100",971 => "01000010",972 => "01111000",973 => "10000111",974 => "00010001",975 => "01010110",976 => "10010110",977 => "10111011",978 => "00010110",979 => "01011100",980 => "11110111",981 => "01000011",982 => "10001001",983 => "11010110",984 => "11000111",985 => "10100010",986 => "00011010",987 => "00111001",988 => "10100110",989 => "11101010",990 => "01000000",991 => "10101011",992 => "00000001",993 => "01101010",994 => "01011100",995 => "10111111",996 => "01001110",997 => "00001010",998 => "11001100",999 => "00111100",1000 => "00001100",1001 => "11111011",1002 => "01111110",1003 => "10010010",1004 => "10010000",1005 => "10000110",1006 => "10100011",1007 => "00101011",1008 => "11000011",1009 => "00111001",1010 => "00100010",1011 => "11111101",1012 => "11100010",1013 => "10101000",1014 => "01111011",1015 => "00010101",1016 => "01000111",1017 => "00001100",1018 => "11011000",1019 => "01100110",1020 => "11000101",1021 => "01001001",1022 => "11001100",1023 => "00100010",1024 => "10000101",1025 => "01010100",1026 => "00101001",1027 => "10000100",1028 => "00100111",1029 => "11010010",1030 => "00011111",1031 => "01111000",1032 => "01011110",1033 => "01111001",1034 => "00011000",1035 => "01001010",1036 => "10111101",1037 => "00010000",1038 => "00111111",1039 => "10110011",1040 => "11011001",1041 => "11111100",1042 => "00111110",1043 => "01001111",1044 => "10110000",1045 => "11000110",1046 => "00111010",1047 => "01110111",1048 => "00010000",1049 => "01111100",1050 => "00010010",1051 => "10111000",1052 => "11101100",1053 => "01001100",1054 => "11000110",1055 => "11000001",1056 => "00111110",1057 => "00001100",1058 => "10001010",1059 => "01001011",1060 => "10111001",1061 => "01011011",1062 => "10100110",1063 => "11001110",1064 => "10101011",1065 => "01101101",1066 => "10111001",1067 => "10010001",1068 => "00100001",1069 => "10100000",1070 => "01111111",1071 => "11100100",1072 => "11000001",1073 => "01011111",1074 => "10001110",1075 => "10000110",1076 => "00010001",1077 => "11110101",1078 => "10111110",1079 => "00000001",1080 => "00000010",1081 => "11100110",1082 => "11010000",1083 => "01101011",1084 => "11101100",1085 => "10011111",1086 => "11000101",1087 => "00010010",1088 => "00001010",1089 => "00001111",1090 => "10011001",1091 => "00011010",1092 => "01111011",1093 => "11110011",1094 => "10100010",1095 => "01110011",1096 => "00111110",1097 => "01001010",1098 => "01011001",1099 => "00001111",1100 => "10011011",1101 => "10110100",1102 => "00101000",1103 => "10100101",1104 => "11110000",1105 => "10101000",1106 => "00000111",1107 => "00111010",1108 => "10000011",1109 => "01000110",1110 => "11110101",1111 => "01101100",1112 => "00011000",1113 => "01001110",1114 => "00100011",1115 => "11000011",1116 => "00101011",1117 => "00011001",1118 => "00100111",1119 => "01010101",1120 => "11000011",1121 => "10110001",1122 => "11111011",1123 => "00101110",1124 => "11101011",1125 => "01000001",1126 => "10010000",1127 => "00100110",1128 => "00111110",1129 => "11010001",1130 => "01111101",1131 => "01010110",1132 => "00000110",1133 => "01100111",1134 => "10110011",1135 => "10101001",1136 => "10011010",1137 => "00110000",1138 => "10110111",1139 => "10011100",1140 => "00001000",1141 => "00101001",1142 => "01011111",1143 => "01011001",1144 => "00100101",1145 => "10001110",1146 => "01100111",1147 => "01010101",1148 => "11011010",1149 => "10111100",1150 => "01001100",1151 => "11011111",1152 => "01010011",1153 => "00000110",1154 => "11101001",1155 => "01101111",1156 => "11011010",1157 => "10110101",1158 => "11111011",1159 => "10011000",1160 => "01111100",1161 => "10110101",1162 => "10110010",1163 => "01010001",1164 => "00101001",1165 => "01000000",1166 => "11000101",1167 => "01010100",1168 => "01010001",1169 => "10110000",1170 => "10101110",1171 => "01010110",1172 => "00000000",1173 => "10010101",1174 => "10110010",1175 => "00110100",1176 => "11101010",1177 => "01101000",1178 => "11111001",1179 => "11010101",1180 => "11000100",1181 => "01100111",1182 => "11000001",1183 => "01010010",1184 => "00010010",1185 => "11101000",1186 => "01101101",1187 => "00111111",1188 => "11101000",1189 => "00110110",1190 => "00011111",1191 => "10101001",1192 => "11011000",1193 => "10100000",1194 => "11011100",1195 => "10100001",1196 => "00100101",1197 => "11011010",1198 => "00111101",1199 => "11011011",1200 => "00110000",1201 => "01111011",1202 => "11011110",1203 => "01110100",1204 => "10100011",1205 => "01001110",1206 => "11110001",1207 => "11101000",1208 => "11001000",1209 => "11011001",1210 => "01101010",1211 => "00010110",1212 => "01001111",1213 => "00100000",1214 => "11000110",1215 => "10001001",1216 => "11000011",1217 => "11010011",1218 => "11100101",1219 => "11000110",1220 => "10010011",1221 => "11110001",1222 => "00010000",1223 => "01111010",1224 => "00000011",1225 => "01011001",1226 => "11100111",1227 => "01101001",1228 => "01011101",1229 => "11010011",1230 => "11011000",1231 => "01101110",1232 => "10101110",1233 => "11010110",1234 => "00010011",1235 => "01000101",1236 => "01110101",1237 => "11011011",1238 => "11010100",1239 => "11100110",1240 => "01111100",1241 => "01100000",1242 => "01101010",1243 => "11000010",1244 => "10100011",1245 => "00011011",1246 => "01011000",1247 => "10110001",1248 => "01111010",1249 => "11001010",1250 => "10000000",1251 => "11000100",1252 => "01101010",1253 => "10111101",1254 => "00001100",1255 => "01010001",1256 => "10011111",1257 => "10000101",1258 => "10010101",1259 => "01011100",1260 => "11110010",1261 => "10011011",1262 => "10000010",1263 => "11100111",1264 => "11011011",1265 => "01110000",1266 => "10110101",1267 => "11001001",1268 => "00111011",1269 => "01101100",1270 => "00001010",1271 => "00111111",1272 => "11001101",1273 => "00011100",1274 => "11111011",1275 => "10011101",1276 => "11000111",1277 => "10101010",1278 => "01010001",1279 => "01101100",1280 => "10010000",1281 => "11000011",1282 => "01011101",1283 => "11011100",1284 => "10111010",1285 => "01010101",1286 => "00000101",1287 => "10000101",1288 => "10000011",1289 => "11111000",1290 => "10100111",1291 => "01010000",1292 => "10101001",1293 => "11000111",1294 => "11010101",1295 => "00100101",1296 => "00110000",1297 => "11010100",1298 => "01101010",1299 => "00011010",1300 => "11100001",1301 => "10011110",1302 => "00010000",1303 => "10010100",1304 => "11000001",1305 => "00001000",1306 => "00100011",1307 => "11001110",1308 => "00010000",1309 => "11101100",1310 => "01100111",1311 => "10100001",1312 => "00010100",1313 => "10101011",1314 => "10111111",1315 => "00110010",1316 => "01110111",1317 => "10001111",1318 => "11101000",1319 => "01001101",1320 => "10001101",1321 => "10101010",1322 => "11111010",1323 => "00111001",1324 => "11100101",1325 => "01011010",1326 => "11110100",1327 => "11001011",1328 => "01101000",1329 => "11111011",1330 => "00100110",1331 => "10011001",1332 => "01011001",1333 => "01111010",1334 => "10000011",1335 => "01010100",1336 => "10101101",1337 => "10111100",1338 => "10010101",1339 => "10000000",1340 => "11110100",1341 => "11101100",1342 => "00100111",1343 => "11110101",1344 => "01000010",1345 => "11011011",1346 => "11101000",1347 => "01101111",1348 => "01101100",1349 => "00011010",1350 => "01001111",1351 => "01100001",1352 => "11101110",1353 => "01011011",1354 => "10101101",1355 => "01101001",1356 => "00101101",1357 => "00111101",1358 => "00100110",1359 => "00010101",1360 => "00010100",1361 => "10110101",1362 => "00100001",1363 => "10111001",1364 => "10110010",1365 => "00001110",1366 => "10000000",1367 => "11000000",1368 => "11100011",1369 => "01101011",1370 => "11000001",1371 => "01011101",1372 => "00001000",1373 => "01111101",1374 => "10001101",1375 => "11011100",1376 => "10011001",1377 => "00011100",1378 => "01111110",1379 => "01010110",1380 => "10100000",1381 => "01110101",1382 => "10010000",1383 => "01011101",1384 => "00100110",1385 => "00010101",1386 => "10011100",1387 => "10111100",1388 => "10010000",1389 => "01010101",1390 => "10011100",1391 => "01001010",1392 => "11010100",1393 => "10010011",1394 => "11000011",1395 => "10110001",1396 => "10111101",1397 => "01101111",1398 => "00100100",1399 => "10010010",1400 => "10100101",1401 => "01011010",1402 => "11001000",1403 => "00110011",1404 => "01000011",1405 => "11100100",1406 => "01001001",1407 => "11111000",1408 => "11111011",1409 => "00100100",1410 => "10101111",1411 => "00010010",1412 => "00101001",1413 => "10000011",1414 => "01011001",1415 => "00111001",1416 => "00111111",1417 => "00011100",1418 => "00010110",1419 => "10010110",1420 => "11111101",1421 => "11101110",1422 => "00000100",1423 => "10010110",1424 => "00111011",1425 => "10101111",1426 => "11011001",1427 => "10010010",1428 => "00101111",1429 => "01000011",1430 => "00011111",1431 => "00100100",1432 => "01010110",1433 => "00110001",1434 => "00000100",1435 => "10000110",1436 => "01000000",1437 => "10100100",1438 => "00110100",1439 => "01111001",1440 => "10010100",1441 => "01100010",1442 => "11111010",1443 => "11000100",1444 => "01000010",1445 => "10010111",1446 => "00010111",1447 => "00011110",1448 => "00111000",1449 => "00010000",1450 => "00101010",1451 => "01000011",1452 => "11100011",1453 => "11101110",1454 => "10001001",1455 => "10001010",1456 => "11011010",1457 => "01011001",1458 => "00011001",1459 => "11101111",1460 => "10100000",1461 => "01111000",1462 => "00100010",1463 => "00010100",1464 => "11100101",1465 => "10100111",1466 => "00101011",1467 => "10111111",1468 => "10101011",1469 => "10110010",1470 => "10111000",1471 => "10111001",1472 => "00110101",1473 => "01110011",1474 => "00010100",1475 => "01111110",1476 => "11100100",1477 => "11110100",1478 => "00111100",1479 => "11010110",1480 => "00001100",1481 => "00010000",1482 => "10100000",1483 => "01011000",1484 => "01000110",1485 => "01101101",1486 => "01100110",1487 => "10001010",1488 => "10000001",1489 => "10110001",1490 => "11110110",1491 => "01110111",1492 => "11010010",1493 => "01001001",1494 => "10100111",1495 => "11000101",1496 => "01100100",1497 => "01000001",1498 => "10100110",1499 => "11100100",1500 => "00000101",1501 => "10101100",1502 => "10111011",1503 => "10010011",1504 => "11000111",1505 => "11111101",1506 => "00010100",1507 => "01001100",1508 => "11001111",1509 => "10011110",1510 => "00011000",1511 => "10010110",1512 => "11001110",1513 => "00000110",1514 => "10000010",1515 => "10010101",1516 => "10101111",1517 => "01110111",1518 => "10110011",1519 => "01100000",1520 => "01111011",1521 => "10110111",1522 => "01010111",1523 => "00111001",1524 => "01100001",1525 => "01000110",1526 => "11000011",1527 => "00101100",1528 => "10100000",1529 => "11100110",1530 => "00011100",1531 => "01111000",1532 => "11011100",1533 => "10110011",1534 => "11011110",1535 => "01110110",1536 => "11101101",1537 => "01100010",1538 => "10010011",1539 => "01101010",1540 => "11010011",1541 => "11011010",1542 => "11111011",1543 => "00010000",1544 => "11100100",1545 => "10001000",1546 => "01010001",1547 => "00010111",1548 => "11111000",1549 => "11100101",1550 => "00111111",1551 => "11001100",1552 => "10110100",1553 => "01111001",1554 => "11111111",1555 => "00001111",1556 => "00110001",1557 => "01010111",1558 => "01110111",1559 => "11010010",1560 => "11000001",1561 => "01110011",1562 => "10011000",1563 => "11110100",1564 => "00010101",1565 => "00100110",1566 => "01011001",1567 => "01101111",1568 => "10111100",1569 => "01111000",1570 => "10101011",1571 => "00001100",1572 => "00001011",1573 => "01100101",1574 => "11100101",1575 => "10000111",1576 => "01010110",1577 => "00111001",1578 => "00000111",1579 => "00000001",1580 => "11001010",1581 => "10101010",1582 => "00011110",1583 => "11011000",1584 => "01110110",1585 => "11101000",1586 => "01101011",1587 => "00111101",1588 => "10100110",1589 => "10101101",1590 => "11010101",1591 => "11000101",1592 => "00000001",1593 => "11110110",1594 => "00000010",1595 => "10101010",1596 => "10100101",1597 => "10110110",1598 => "00111111",1599 => "01001001",1600 => "00100001",1601 => "11101001",1602 => "10010101",1603 => "11000111",1604 => "01100101",1605 => "11011000",1606 => "01010111",1607 => "00101010",1608 => "11100011",1609 => "00100000",1610 => "10010101",1611 => "01111010",1612 => "11000010",1613 => "10111110",1614 => "10011011",1615 => "10001100",1616 => "01110111",1617 => "11110001",1618 => "11111110",1619 => "00101011",1620 => "00000011",1621 => "00001110",1622 => "10100111",1623 => "10011100",1624 => "11101101",1625 => "11101100",1626 => "01001011",1627 => "10011010",1628 => "01110011",1629 => "00101100",1630 => "01000111",1631 => "01101101",1632 => "11000000",1633 => "10110101",1634 => "10001010",1635 => "10001101",1636 => "01110010",1637 => "10011101",1638 => "01000111",1639 => "01110101",1640 => "11001110",1641 => "10110101",1642 => "11000111",1643 => "11010000",1644 => "00010100",1645 => "11000101",1646 => "00001110",1647 => "00011000",1648 => "11010010",1649 => "10011111",1650 => "00101000",1651 => "11100101",1652 => "01010000",1653 => "01101010",1654 => "10000101",1655 => "10110010",1656 => "10010110",1657 => "00100000",1658 => "10101110",1659 => "00011101",1660 => "00111011",1661 => "00010101",1662 => "01000011",1663 => "00111101",1664 => "01110111",1665 => "00110111",1666 => "00110010",1667 => "01100111",1668 => "01010010",1669 => "00101111",1670 => "00010111",1671 => "10110100",1672 => "10100000",1673 => "01100001",1674 => "00110110",1675 => "10001000",1676 => "01101010",1677 => "01111101",1678 => "01011011",1679 => "00000010",1680 => "10111000",1681 => "00110111",1682 => "01011010",1683 => "01101000",1684 => "00101100",1685 => "00101101",1686 => "11010010",1687 => "00011110",1688 => "10100100",1689 => "11000111",1690 => "00011000",1691 => "01001101",1692 => "01110000",1693 => "10001010",1694 => "11101010",1695 => "10101001",1696 => "11101010",1697 => "10110101",1698 => "11010110",1699 => "01001001",1700 => "11111011",1701 => "11100111",1702 => "01100111",1703 => "11000000",1704 => "00011101",1705 => "10110100",1706 => "11111101",1707 => "11011100",1708 => "10000111",1709 => "11111001",1710 => "11000100",1711 => "01110001",1712 => "01110001",1713 => "11010100",1714 => "10110000",1715 => "10010110",1716 => "10001110",1717 => "10011010",1718 => "10011000",1719 => "11000011",1720 => "01100101",1721 => "10110011",1722 => "11100111",1723 => "00110010",1724 => "00110110",1725 => "00111101",1726 => "11110100",1727 => "01000010",1728 => "01010111",1729 => "00000001",1730 => "00100100",1731 => "10010010",1732 => "00110011",1733 => "11101110",1734 => "00100110",1735 => "10101000",1736 => "01010010",1737 => "10000001",1738 => "10010010",1739 => "00100101",1740 => "01100111",1741 => "11110101",1742 => "00010101",1743 => "10010100",1744 => "10101101",1745 => "10000010",1746 => "11101111",1747 => "10000110",1748 => "10100011",1749 => "11110010",1750 => "00011011",1751 => "10001010",1752 => "10001111",1753 => "01001101",1754 => "00000100",1755 => "11010110",1756 => "00100101",1757 => "11111101",1758 => "01011011",1759 => "01100011",1760 => "01001011",1761 => "01011011",1762 => "10010101",1763 => "10110010",1764 => "01101101",1765 => "11110111",1766 => "10110000",1767 => "11110110",1768 => "10000110",1769 => "01000000",1770 => "10011110",1771 => "10111100",1772 => "00001111",1773 => "11010100",1774 => "00111101",1775 => "01011101",1776 => "01010110",1777 => "01011101",1778 => "00111001",1779 => "00101010",1780 => "00101111",1781 => "01010000",1782 => "01101001",1783 => "00000110",1784 => "01010101",1785 => "11100001",1786 => "01000111",1787 => "11101100",1788 => "00010100",1789 => "00101100",1790 => "10101110",1791 => "10011010",1792 => "11111110",1793 => "01001010",1794 => "01101101",1795 => "01110100",1796 => "10110100",1797 => "01110110",1798 => "11011100",1799 => "00100110",1800 => "00110001",1801 => "10001110",1802 => "00111101",1803 => "11001000",1804 => "00000011",1805 => "10001010",1806 => "00101101",1807 => "01100110",1808 => "10011011",1809 => "11001100",1810 => "11110011",1811 => "10011010",1812 => "01001001",1813 => "10110000",1814 => "11111100",1815 => "00101111",1816 => "00110010",1817 => "10001111",1818 => "01010000",1819 => "10011000",1820 => "00110100",1821 => "10000100",1822 => "01101000",1823 => "00111001",1824 => "00000000",1825 => "10110000",1826 => "11110000",1827 => "00011111",1828 => "10011110",1829 => "01111001",1830 => "01010101",1831 => "10111000",1832 => "10111110",1833 => "00010010",1834 => "10100101",1835 => "11110010",1836 => "00111101",1837 => "00101110",1838 => "10001111",1839 => "00010101",1840 => "11110111",1841 => "00000010",1842 => "11111110",1843 => "00111000",1844 => "00011011",1845 => "10010101",1846 => "01110111",1847 => "00001001",1848 => "10111001",1849 => "01011001",1850 => "01011001",1851 => "01010011",1852 => "01001001",1853 => "11001101",1854 => "11110101",1855 => "01110110",1856 => "01110000",1857 => "00111111",1858 => "01011000",1859 => "11111011",1860 => "01101011",1861 => "01011100",1862 => "10001001",1863 => "11111000",1864 => "01001010",1865 => "10001100",1866 => "01011101",1867 => "01111010",1868 => "11100111",1869 => "00010001",1870 => "10101101",1871 => "01100111",1872 => "01011001",1873 => "11000111",1874 => "11101111",1875 => "01110001",1876 => "01111111",1877 => "10001011",1878 => "01001111",1879 => "10110010",1880 => "00000001",1881 => "10001000",1882 => "10111001",1883 => "11001001",1884 => "00101010",1885 => "10111011",1886 => "00111001",1887 => "10100110",1888 => "11011110",1889 => "11100011",1890 => "01101001",1891 => "00101001",1892 => "10101101",1893 => "11101000",1894 => "10110011",1895 => "11100110",1896 => "11100101",1897 => "11000101",1898 => "11100010",1899 => "00001111",1900 => "11101110",1901 => "01010001",1902 => "11110000",1903 => "01101100",1904 => "10010110",1905 => "10100101",1906 => "01101101",1907 => "11110010",1908 => "10000010",1909 => "11100011",1910 => "01011111",1911 => "10100001",1912 => "00111001",1913 => "10111010",1914 => "01100000",1915 => "01010011",1916 => "00111111",1917 => "00111000",1918 => "10011011",1919 => "10001000",1920 => "10001111",1921 => "01001110",1922 => "00001110",1923 => "00100110",1924 => "00000101",1925 => "00001001",1926 => "11100111",1927 => "01100101",1928 => "11110010",1929 => "00111011",1930 => "11101101",1931 => "10000000",1932 => "00100010",1933 => "10010001",1934 => "00111111",1935 => "00001000",1936 => "01011111",1937 => "10001001",1938 => "01110011",1939 => "10101101",1940 => "10010111",1941 => "00001101",1942 => "10110100",1943 => "11011000",1944 => "01001010",1945 => "01101001",1946 => "01100011",1947 => "10010011",1948 => "11000111",1949 => "10010100",1950 => "11011000",1951 => "00001101",1952 => "11011001",1953 => "10011100",1954 => "00010111",1955 => "11000000",1956 => "00100001",1957 => "00011110",1958 => "01100010",1959 => "10010011",1960 => "01110101",1961 => "00101110",1962 => "01000111",1963 => "00001101",1964 => "00110011",1965 => "01110111",1966 => "10000011",1967 => "11010000",1968 => "11001011",1969 => "00010100",1970 => "01011101",1971 => "00010111",1972 => "11010001",1973 => "10010000",1974 => "00011111",1975 => "00111001",1976 => "11001010",1977 => "10001000",1978 => "00111001",1979 => "00110101",1980 => "00011110",1981 => "10001110",1982 => "11111010",1983 => "01001111",1984 => "00001111",1985 => "11101111",1986 => "01000100",1987 => "01001100",1988 => "01101111",1989 => "00111100",1990 => "10100010",1991 => "10011001",1992 => "01100110",1993 => "11111010",1994 => "00110010",1995 => "00111110",1996 => "11101110",1997 => "10001101",1998 => "11011001",1999 => "01001111",2000 => "11110010",2001 => "01001000",2002 => "10110001",2003 => "10010110",2004 => "00100110",2005 => "00101101",2006 => "01010010",2007 => "00001010",2008 => "11011100",2009 => "10000010",2010 => "11010111",2011 => "11001110",2012 => "01011001",2013 => "00110101",2014 => "01100110",2015 => "11011010",2016 => "00111100",2017 => "01000111",2018 => "01010010",2019 => "00111100",2020 => "00010010",2021 => "00101011",2022 => "01111100",2023 => "00000001",2024 => "11010000",2025 => "00011001",2026 => "11000100",2027 => "10111101",2028 => "01101100",2029 => "10101001",2030 => "01100111",2031 => "00010011",2032 => "11100111",2033 => "00100001",2034 => "01000010",2035 => "00110010",2036 => "10000000",2037 => "10000111",2038 => "11111111",2039 => "00101111",2040 => "00011111",2041 => "01011110",2042 => "10010111",2043 => "11101111",2044 => "00100010",2045 => "11100011",2046 => "11010111",2047 => "01011100",2048 => "01000000",2049 => "00000100",2050 => "00001111",2051 => "11001111",2052 => "01110111",2053 => "10100001",2054 => "11010011",2055 => "01111101",2056 => "10110000",2057 => "10111110",2058 => "11001111",2059 => "11000110",2060 => "11110001",2061 => "11000000",2062 => "10011001",2063 => "00001110",2064 => "11001100",2065 => "01001001",2066 => "00100011",2067 => "00001000",2068 => "00001101",2069 => "01101111",2070 => "10011011",2071 => "11001011",2072 => "00011111",2073 => "10111000",2074 => "11001001",2075 => "11101101",2076 => "00111110",2077 => "01001111",2078 => "01001111",2079 => "00110101",2080 => "01010111",2081 => "10110111",2082 => "11110000",2083 => "01001101",2084 => "11100011",2085 => "00101111",2086 => "11111100",2087 => "01110001",2088 => "10010001",2089 => "01111010",2090 => "10011110",2091 => "01011111",2092 => "01101011",2093 => "11001000",2094 => "00110101",2095 => "00100101",2096 => "01110100",2097 => "00011111",2098 => "11101101",2099 => "00001001",2100 => "10000101",2101 => "01101001",2102 => "00101101",2103 => "01101001",2104 => "11010000",2105 => "00110001",2106 => "01011000",2107 => "00111111",2108 => "10101101",2109 => "11011110",2110 => "10110000",2111 => "10111000",2112 => "10100111",2113 => "10101000",2114 => "10010101",2115 => "00110001",2116 => "11010010",2117 => "11111000",2118 => "01111100",2119 => "11011101",2120 => "00110010",2121 => "00111000",2122 => "00111111",2123 => "10110000",2124 => "10110010",2125 => "01111010",2126 => "11100010",2127 => "10000000",2128 => "01011110",2129 => "00101011",2130 => "10000010",2131 => "01011011",2132 => "00111110",2133 => "11000000",2134 => "00101100",2135 => "01001010",2136 => "11101101",2137 => "00110110",2138 => "00111001",2139 => "00110000",2140 => "11111010",2141 => "01111010",2142 => "11010100",2143 => "10000010",2144 => "11010000",2145 => "00010011",2146 => "10111101",2147 => "10000001",2148 => "00000101",2149 => "11000111",2150 => "10010000",2151 => "11001101",2152 => "00001100",2153 => "01010111",2154 => "11011011",2155 => "00000001",2156 => "10011101",2157 => "11110100",2158 => "10100010",2159 => "01010011",2160 => "10010101",2161 => "10001001",2162 => "10111100",2163 => "00001000",2164 => "01111110",2165 => "11100100",2166 => "01000011",2167 => "01110101",2168 => "01011001",2169 => "01000110",2170 => "01111100",2171 => "11010111",2172 => "00001011",2173 => "11110000",2174 => "11000100",2175 => "01100100",2176 => "11011000",2177 => "10011010",2178 => "00010010",2179 => "00111110",2180 => "01010100",2181 => "01111100",2182 => "01011110",2183 => "10101101",2184 => "00101001",2185 => "10101111",2186 => "00011001",2187 => "10110100",2188 => "00101000",2189 => "01011111",2190 => "11010001",2191 => "10111001",2192 => "01010101",2193 => "01101111",2194 => "11101110",2195 => "01001001",2196 => "11011001",2197 => "10101110",2198 => "11010000",2199 => "01000010",2200 => "01101010",2201 => "01010000",2202 => "00011010",2203 => "11011011",2204 => "00110100",2205 => "01110000",2206 => "00100110",2207 => "00001101",2208 => "11011010",2209 => "10010100",2210 => "01100011",2211 => "11010110",2212 => "00100110",2213 => "01010110",2214 => "00010011",2215 => "10111010",2216 => "11101010",2217 => "11101100",2218 => "01100110",2219 => "00101101",2220 => "10100001",2221 => "10001101",2222 => "00001101",2223 => "11010010",2224 => "00001101",2225 => "11010110",2226 => "11110111",2227 => "11011110",2228 => "01111001",2229 => "10110011",2230 => "01100011",2231 => "01111101",2232 => "01000101",2233 => "10000001",2234 => "11001011",2235 => "11110110",2236 => "00000011",2237 => "00110101",2238 => "00101111",2239 => "01101100",2240 => "00101011",2241 => "11001000",2242 => "01010011",2243 => "11011011",2244 => "10001000",2245 => "11011001",2246 => "10101101",2247 => "11001110",2248 => "00110001",2249 => "11001110",2250 => "01011100",2251 => "10001101",2252 => "00010111",2253 => "00111101",2254 => "10100011",2255 => "01010000",2256 => "11001111",2257 => "10001010",2258 => "00001000",2259 => "01111110",2260 => "11000100",2261 => "11101010",2262 => "00100010",2263 => "10111010",2264 => "11000010",2265 => "10000011",2266 => "00111110",2267 => "00000100",2268 => "10110010",2269 => "00110000",2270 => "00000111",2271 => "11101000",2272 => "10110011",2273 => "01001100",2274 => "00100010",2275 => "11011000",2276 => "11101110",2277 => "10001000",2278 => "10111101",2279 => "11110011",2280 => "01011101",2281 => "11111001",2282 => "00001010",2283 => "10101111",2284 => "00010110",2285 => "11111010",2286 => "11010000",2287 => "11101010",2288 => "00101101",2289 => "10101010",2290 => "01111010",2291 => "11111101",2292 => "00101000",2293 => "11001011",2294 => "01011111",2295 => "11001111",2296 => "00101100",2297 => "00111000",2298 => "10111111",2299 => "01101011",2300 => "10100100",2301 => "11101000",2302 => "00101111",2303 => "00001001",2304 => "00110110",2305 => "01110111",2306 => "11100100",2307 => "11000000",2308 => "01010101",2309 => "11101111",2310 => "00001011",2311 => "11000000",2312 => "10100101",2313 => "01001010",2314 => "01011110",2315 => "01101010",2316 => "11001011",2317 => "00110101",2318 => "01000011",2319 => "11001101",2320 => "10101010",2321 => "01111000",2322 => "01111000",2323 => "11011000",2324 => "00000110",2325 => "01101110",2326 => "11001110",2327 => "01001001",2328 => "00101010",2329 => "11010010",2330 => "11100000",2331 => "00000101",2332 => "11100001",2333 => "11100100",2334 => "01011101",2335 => "00110100",2336 => "10010111",2337 => "10100110",2338 => "01101110",2339 => "10011011",2340 => "01000011",2341 => "10111000",2342 => "01100011",2343 => "00111000",2344 => "00110000",2345 => "00010111",2346 => "01110110",2347 => "11101111",2348 => "11110110",2349 => "00100001",2350 => "01111011",2351 => "11100100",2352 => "00000101",2353 => "00100101",2354 => "00110010",2355 => "10010001",2356 => "11001111",2357 => "10011000",2358 => "01001111",2359 => "00000110",2360 => "10101100",2361 => "01110110",2362 => "11101101",2363 => "11000010",2364 => "11111101",2365 => "01110011",2366 => "10001101",2367 => "00100111",2368 => "00101010",2369 => "00011110",2370 => "00001100",2371 => "01100101",2372 => "01000101",2373 => "01110101",2374 => "10010101",2375 => "11101010",2376 => "01111000",2377 => "00000110",2378 => "10001101",2379 => "01111010",2380 => "10111111",2381 => "01011100",2382 => "00000010",2383 => "01000000",2384 => "10110001",2385 => "10011011",2386 => "01010100",2387 => "11100001",2388 => "01001010",2389 => "00101110",2390 => "00100100",2391 => "00001101",2392 => "10011100",2393 => "01010010",2394 => "10111101",2395 => "01100000",2396 => "11001000",2397 => "00010101",2398 => "00001101",2399 => "11000011",2400 => "10111111",2401 => "01011011",2402 => "11010100",2403 => "10011000",2404 => "00010111",2405 => "01110000",2406 => "01001101",2407 => "01010111",2408 => "11001111",2409 => "11101101",2410 => "01101111",2411 => "10101110",2412 => "10111000",2413 => "10010011",2414 => "00101111",2415 => "00111111",2416 => "11000101",2417 => "00110001",2418 => "10000101",2419 => "00011000",2420 => "11011011",2421 => "01000011",2422 => "01101010",2423 => "01101111",2424 => "11001111",2425 => "00100100",2426 => "10011000",2427 => "00111100",2428 => "11100000",2429 => "01101010",2430 => "01101101",2431 => "11001100",2432 => "01000011",2433 => "00110101",2434 => "00001000",2435 => "10001001",2436 => "10100110",2437 => "10110010",2438 => "10000100",2439 => "10001010",2440 => "10101011",2441 => "10010011",2442 => "11111111",2443 => "01011101",2444 => "01010101",2445 => "10011011",2446 => "11000100",2447 => "11110011",2448 => "00001000",2449 => "11111010",2450 => "10001111",2451 => "00110001",2452 => "10010101",2453 => "00111010",2454 => "11000001",2455 => "10100001",2456 => "01000110",2457 => "00110000",2458 => "11000010",2459 => "10010000",2460 => "11110000",2461 => "01010000",2462 => "11110000",2463 => "10100111",2464 => "00101001",2465 => "11000101",2466 => "11000000",2467 => "10101000",2468 => "01011011",2469 => "01110100",2470 => "01110000",2471 => "11001010",2472 => "10100101",2473 => "01001001",2474 => "11010000",2475 => "11101001",2476 => "01000110",2477 => "00001001",2478 => "10101110",2479 => "01111110",2480 => "01111110",2481 => "01101111",2482 => "00001101",2483 => "01000110",2484 => "11100000",2485 => "01110110",2486 => "01100001",2487 => "01010010",2488 => "10111100",2489 => "01110011",2490 => "11000000",2491 => "01111000",2492 => "10001101",2493 => "11000111",2494 => "00001000",2495 => "11011010",2496 => "01101111",2497 => "11011010",2498 => "01111111",2499 => "11001000",2500 => "10001100",2501 => "01111011",2502 => "10010100",2503 => "00000001",2504 => "01110101",2505 => "01001001",2506 => "00001110",2507 => "11011100",2508 => "10111010",2509 => "01101111",2510 => "11110110",2511 => "10101111",2512 => "01111111",2513 => "00100001",2514 => "01001101",2515 => "11001111",2516 => "10110101",2517 => "00101010",2518 => "01001111",2519 => "10000010",2520 => "01111001",2521 => "11100110",2522 => "10010100",2523 => "11001010",2524 => "00010101",2525 => "10111111",2526 => "01010001",2527 => "01011110",2528 => "10000000",2529 => "11101010",2530 => "10110000",2531 => "00111111",2532 => "10110011",2533 => "01111000",2534 => "01011110",2535 => "10011011",2536 => "11000001",2537 => "01111011",2538 => "10011110",2539 => "01101011",2540 => "11001010",2541 => "01010101",2542 => "11011001",2543 => "00001000",2544 => "10000110",2545 => "00010001",2546 => "10111011",2547 => "00100011",2548 => "01001100",2549 => "00101110",2550 => "00101010",2551 => "10011001",2552 => "01100011",2553 => "10110110",2554 => "00100111",2555 => "10010101",2556 => "11110110",2557 => "00001101",2558 => "01011011",2559 => "00010000",2560 => "11011011",2561 => "11001000",2562 => "01100111",2563 => "10000001",2564 => "01011001",2565 => "00100111",2566 => "00111110",2567 => "10110001",2568 => "11000110",2569 => "10001010",2570 => "11000111",2571 => "10100010",2572 => "00000110",2573 => "00000101",2574 => "10010001",2575 => "11000010",2576 => "11000010",2577 => "11010110",2578 => "10100011",2579 => "01111011",2580 => "11000001",2581 => "01010101",2582 => "11100001",2583 => "00111010",2584 => "00100100",2585 => "11000011",2586 => "00001110",2587 => "01010110",2588 => "00010111",2589 => "00000100",2590 => "00100101",2591 => "11110001",2592 => "11001010",2593 => "11110010",2594 => "11111001",2595 => "00000001",2596 => "01100101",2597 => "11000110",2598 => "01010001",2599 => "11110100",2600 => "10111001",2601 => "10011011",2602 => "11011010",2603 => "01110010",2604 => "00101110",2605 => "11001011",2606 => "11011111",2607 => "11101111",2608 => "10011001",2609 => "01111101",2610 => "10101101",2611 => "01110010",2612 => "01010101",2613 => "00000010",2614 => "01110111",2615 => "11011001",2616 => "01000001",2617 => "11111011",2618 => "10000100",2619 => "01100001",2620 => "00101111",2621 => "10000001",2622 => "10001101",2623 => "00011011",2624 => "01100101",2625 => "01011111",2626 => "11100111",2627 => "10110011",2628 => "00001111",2629 => "00001000",2630 => "01110010",2631 => "11100111",2632 => "01010111",2633 => "10000101",2634 => "10100000",2635 => "01110001",2636 => "01001110",2637 => "01001101",2638 => "10100001",2639 => "01100010",2640 => "00111101",2641 => "00110011",2642 => "10111010",2643 => "10011100",2644 => "10001110",2645 => "00001101",2646 => "10001111",2647 => "11110011",2648 => "11110110",2649 => "11011010",2650 => "00101011",2651 => "11110111",2652 => "01010111",2653 => "11110110",2654 => "11001101",2655 => "01000011",2656 => "01100101",2657 => "00101001",2658 => "00110101",2659 => "11001010",2660 => "11010010",2661 => "11100011",2662 => "10010101",2663 => "00010100",2664 => "10100000",2665 => "10101011",2666 => "10001110",2667 => "01001101",2668 => "01101011",2669 => "00100011",2670 => "10100100",2671 => "10100100",2672 => "00101001",2673 => "11001010",2674 => "00001110",2675 => "00110000",2676 => "11011101",2677 => "10010010",2678 => "11110100",2679 => "10000001",2680 => "10111000",2681 => "10010000",2682 => "01011111",2683 => "00101100",2684 => "01001011",2685 => "00010110",2686 => "11001010",2687 => "11101100",2688 => "00001011",2689 => "01001100",2690 => "01110010",2691 => "11010101",2692 => "10001011",2693 => "11100011",2694 => "01101011",2695 => "11101100",2696 => "00011011",2697 => "11000100",2698 => "10101011",2699 => "00110000",2700 => "10100111",2701 => "11110011",2702 => "10011111",2703 => "00000011",2704 => "01111100",2705 => "10111000",2706 => "01010111",2707 => "01000000",2708 => "10001101",2709 => "01001000",2710 => "10001000",2711 => "11111011",2712 => "10011010",2713 => "00100100",2714 => "01010010",2715 => "01000010",2716 => "11100011",2717 => "00010110",2718 => "00000100",2719 => "01010001",2720 => "01110010",2721 => "10010011",2722 => "10000111",2723 => "01000001",2724 => "11011111",2725 => "11100101",2726 => "11111111",2727 => "00001100",2728 => "10101111",2729 => "01001101",2730 => "01010101",2731 => "11000000",2732 => "01101000",2733 => "00100000",2734 => "11000100",2735 => "10110001",2736 => "00011110",2737 => "10010110",2738 => "01110111",2739 => "01111111",2740 => "11110000",2741 => "11001001",2742 => "11100111",2743 => "10111100",2744 => "00111111",2745 => "01100110",2746 => "01101001",2747 => "01001100",2748 => "01100110",2749 => "11010111",2750 => "10110001",2751 => "00111100",2752 => "01111001",2753 => "01010110",2754 => "00010101",2755 => "10001011",2756 => "10000000",2757 => "00110010",2758 => "11110011",2759 => "11001110",2760 => "11001110",2761 => "01000000",2762 => "00100010",2763 => "10011111",2764 => "01111011",2765 => "01110110",2766 => "00111010",2767 => "10110111",2768 => "11001101",2769 => "11101100",2770 => "01111011",2771 => "10110110",2772 => "10000111",2773 => "10001111",2774 => "11111011",2775 => "11111101",2776 => "11111111",2777 => "00001011",2778 => "01111010",2779 => "00010011",2780 => "10101000",2781 => "10010011",2782 => "00001001",2783 => "01000010",2784 => "01100011",2785 => "10000001",2786 => "01010011",2787 => "10110001",2788 => "00010101",2789 => "10101000",2790 => "01100001",2791 => "00001111",2792 => "00110000",2793 => "00011010",2794 => "11101001",2795 => "11101100",2796 => "10100010",2797 => "01001011",2798 => "00101010",2799 => "11100001",2800 => "10100011",2801 => "01001100",2802 => "10001010",2803 => "10000011",2804 => "10111010",2805 => "00101000",2806 => "10000011",2807 => "00010000",2808 => "01100111",2809 => "00001111",2810 => "10111101",2811 => "01100011",2812 => "11101100",2813 => "00011001",2814 => "00100110",2815 => "11001101",2816 => "00001111",2817 => "00101111",2818 => "01001000",2819 => "10111101",2820 => "11011110",2821 => "11100111",2822 => "10100110",2823 => "11000010",2824 => "00001000",2825 => "10100111",2826 => "11010001",2827 => "10100110",2828 => "00100001",2829 => "01111010",2830 => "00110110",2831 => "10110110",2832 => "01010010",2833 => "00011100",2834 => "00101011",2835 => "10100101",2836 => "01110101",2837 => "11000010",2838 => "01101110",2839 => "00101100",2840 => "00010001",2841 => "11001111",2842 => "10111000",2843 => "11001001",2844 => "00000001",2845 => "01001010",2846 => "01101001",2847 => "11100110",2848 => "00110110",2849 => "11011001",2850 => "00000110",2851 => "00010000",2852 => "01111100",2853 => "11111011",2854 => "01000101",2855 => "11101011",2856 => "01111000",2857 => "01001011",2858 => "11011110",2859 => "10010010",2860 => "00111101",2861 => "01100001",2862 => "10001011",2863 => "00111100",2864 => "01100111",2865 => "10011101",2866 => "10000111",2867 => "01000110",2868 => "10011000",2869 => "10100001",2870 => "11011111",2871 => "00101100",2872 => "00110010",2873 => "11010010",2874 => "11110011",2875 => "00111001",2876 => "01010001",2877 => "11001001",2878 => "00010001",2879 => "10000000",2880 => "01111010",2881 => "11010101",2882 => "11000010",2883 => "00101001",2884 => "11111010",2885 => "01110000",2886 => "10000001",2887 => "11000001",2888 => "11110011",2889 => "01001101",2890 => "01011001",2891 => "01110101",2892 => "10100110",2893 => "00111001",2894 => "11010101",2895 => "01011010",2896 => "10111111",2897 => "01001000",2898 => "01101000",2899 => "01000011",2900 => "10010010",2901 => "10001111",2902 => "10111101",2903 => "10000111",2904 => "10000111",2905 => "10001111",2906 => "00101001",2907 => "10100001",2908 => "00100111",2909 => "10011000",2910 => "10000011",2911 => "11001001",2912 => "11000100",2913 => "10111110",2914 => "10101100",2915 => "01000001",2916 => "00111110",2917 => "10100001",2918 => "00100100",2919 => "01001010",2920 => "01010100",2921 => "11110010",2922 => "11111011",2923 => "11001001",2924 => "01111010",2925 => "10111111",2926 => "11111101",2927 => "00111001",2928 => "11001111",2929 => "00100000",2930 => "11001101",2931 => "00010100",2932 => "00101110",2933 => "10111010",2934 => "00101010",2935 => "01011010",2936 => "11000100",2937 => "10111100",2938 => "11111001",2939 => "10010100",2940 => "10001101",2941 => "00111110",2942 => "01110101",2943 => "01010111",2944 => "11001010",2945 => "01100111",2946 => "10001101",2947 => "01000010",2948 => "01100100",2949 => "11100110",2950 => "01111110",2951 => "01001100",2952 => "11101010",2953 => "00001011",2954 => "10110000",2955 => "01100101",2956 => "00111100",2957 => "01010000",2958 => "11000011",2959 => "11001011",2960 => "01101000",2961 => "11000110",2962 => "00001101",2963 => "11111101",2964 => "00000001",2965 => "11001001",2966 => "01000001",2967 => "00101010",2968 => "00000100",2969 => "01001000",2970 => "11001110",2971 => "00011110",2972 => "01010001",2973 => "11000011",2974 => "00011011",2975 => "01001001",2976 => "00111101",2977 => "11000001",2978 => "10111000",2979 => "01011111",2980 => "01011100",2981 => "00111000",2982 => "00101101",2983 => "01110001",2984 => "01100001",2985 => "11111110",2986 => "11111111",2987 => "00001011",2988 => "00010111",2989 => "00011100",2990 => "10101110",2991 => "11000110",2992 => "00100111",2993 => "11001001",2994 => "11100110",2995 => "11010000",2996 => "11110001",2997 => "10010110",2998 => "11110001",2999 => "01111100",3000 => "00110011",3001 => "00000001",3002 => "01000111",3003 => "11101011",3004 => "00101111",3005 => "01110111",3006 => "01110100",3007 => "10101110",3008 => "11010110",3009 => "00111101",3010 => "00100111",3011 => "11010000",3012 => "10011111",3013 => "01011010",3014 => "11110100",3015 => "11110011",3016 => "10010000",3017 => "00011111",3018 => "10101011",3019 => "01100001",3020 => "00101101",3021 => "11010100",3022 => "00010101",3023 => "10000001",3024 => "11010101",3025 => "01111110",3026 => "00101110",3027 => "11101111",3028 => "11000100",3029 => "01100010",3030 => "11001010",3031 => "11010000",3032 => "01010100",3033 => "00010010",3034 => "11100100",3035 => "10111000",3036 => "11001000",3037 => "11010110",3038 => "01011011",3039 => "10110001",3040 => "00110111",3041 => "10110001",3042 => "10100011",3043 => "11011000",3044 => "10010110",3045 => "01101001",3046 => "11000000",3047 => "01001101",3048 => "00011100",3049 => "10101001",3050 => "10101001",3051 => "11111001",3052 => "10100001",3053 => "11010101",3054 => "10010010",3055 => "01101110",3056 => "00000010",3057 => "00000101",3058 => "00101101",3059 => "00111011",3060 => "00100001",3061 => "00011111",3062 => "11011101",3063 => "01011000",3064 => "01111101",3065 => "01011001",3066 => "10101101",3067 => "10000110",3068 => "11110110",3069 => "10100111",3070 => "11001001",3071 => "00100000",3072 => "10100110",3073 => "01000110",3074 => "00001111",3075 => "00010101",3076 => "00111000",3077 => "10100111",3078 => "00001111",3079 => "00000101",3080 => "01100111",3081 => "10000001",3082 => "00110000",3083 => "00000000",3084 => "00111001",3085 => "01101110",3086 => "00001010",3087 => "10111010",3088 => "00100001",3089 => "01011010",3090 => "11001010",3091 => "10100000",3092 => "00011001",3093 => "10011010",3094 => "01100001",3095 => "01101111",3096 => "10100011",3097 => "10101101",3098 => "01000000",3099 => "00000111",3100 => "11100001",3101 => "11011110",3102 => "11110000",3103 => "01010001",3104 => "10010110",3105 => "00001111",3106 => "10010100",3107 => "00011111",3108 => "11011010",3109 => "00110010",3110 => "10100110",3111 => "10111101",3112 => "00100101",3113 => "11011000",3114 => "10000101",3115 => "10110100",3116 => "10010001",3117 => "11011110",3118 => "11010001",3119 => "00110010",3120 => "00000001",3121 => "10001000",3122 => "11110100",3123 => "10001000",3124 => "10010000",3125 => "00100011",3126 => "00011110",3127 => "10111011",3128 => "00001101",3129 => "10010011",3130 => "01010000",3131 => "10110001",3132 => "10101111",3133 => "10000101",3134 => "01011011",3135 => "01000010",3136 => "11111111",3137 => "00001110",3138 => "10011010",3139 => "10100111",3140 => "00110100",3141 => "01110101",3142 => "00011001",3143 => "11101000",3144 => "10001011",3145 => "00011000",3146 => "00001110",3147 => "00000111",3148 => "11001010",3149 => "01100000",3150 => "11011001",3151 => "10010101",3152 => "00001101",3153 => "01000110",3154 => "00010000",3155 => "11111110",3156 => "01000111",3157 => "00100111",3158 => "00011011",3159 => "01111011",3160 => "00101101",3161 => "00010101",3162 => "01001000",3163 => "11011010",3164 => "11010110",3165 => "00001000",3166 => "01001100",3167 => "00011111",3168 => "11000011",3169 => "10101000",3170 => "10101101",3171 => "10101101",3172 => "00010000",3173 => "00011000",3174 => "10011101",3175 => "01001001",3176 => "10011110",3177 => "10000011",3178 => "11001011",3179 => "01000000",3180 => "11011000",3181 => "00101111",3182 => "11001010",3183 => "01001000",3184 => "11001010",3185 => "11111101",3186 => "10010101",3187 => "01110100",3188 => "10011101",3189 => "11110111",3190 => "10100110",3191 => "01000100",3192 => "00001101",3193 => "00001001",3194 => "11011110",3195 => "00010010",3196 => "01110110",3197 => "00011111",3198 => "10000010",3199 => "01101011",3200 => "00001101",3201 => "00111101",3202 => "10110101",3203 => "11100010",3204 => "11110011",3205 => "11001000",3206 => "10011110",3207 => "10110001",3208 => "01111110",3209 => "11010111",3210 => "11010010",3211 => "11101010",3212 => "00010001",3213 => "00101001",3214 => "01111011",3215 => "11010011",3216 => "11001110",3217 => "01111011",3218 => "00000001",3219 => "01100110",3220 => "10110100",3221 => "11110100",3222 => "01110101",3223 => "11101111",3224 => "11111101",3225 => "00111101",3226 => "00011011",3227 => "01011101",3228 => "00100000",3229 => "00000000",3230 => "00001101",3231 => "00110110",3232 => "01100111",3233 => "01101001",3234 => "11011001",3235 => "11011001",3236 => "01101010",3237 => "10100111",3238 => "11011101",3239 => "11100010",3240 => "00110100",3241 => "11110011",3242 => "00010101",3243 => "01110110",3244 => "11010110",3245 => "00010100",3246 => "10101110",3247 => "10110110",3248 => "11010011",3249 => "01101100",3250 => "00001001",3251 => "10101010",3252 => "01010000",3253 => "11011100",3254 => "11100101",3255 => "00000111",3256 => "11011100",3257 => "10110111",3258 => "11001101",3259 => "01101110",3260 => "10001000",3261 => "11110000",3262 => "10001111",3263 => "11100111",3264 => "11110111",3265 => "11101110",3266 => "00011100",3267 => "01010110",3268 => "11001111",3269 => "10101000",3270 => "11110101",3271 => "11010000",3272 => "00110000",3273 => "11100111",3274 => "01100111",3275 => "10001111",3276 => "11111010",3277 => "10111010",3278 => "10110110",3279 => "00011001",3280 => "11000010",3281 => "00010000",3282 => "00111101",3283 => "11110001",3284 => "01000010",3285 => "01111101",3286 => "11011101",3287 => "11100101",3288 => "11100010",3289 => "10000001",3290 => "10010100",3291 => "00001100",3292 => "00101101",3293 => "01101011",3294 => "01111000",3295 => "11000001",3296 => "10111110",3297 => "10110101",3298 => "10111110",3299 => "01011010",3300 => "00100100",3301 => "11000000",3302 => "10110001",3303 => "00111010",3304 => "00111100",3305 => "11111010",3306 => "01011100",3307 => "11100010",3308 => "10111010",3309 => "01011000",3310 => "11000000",3311 => "00110010",3312 => "00010000",3313 => "10111001",3314 => "00001001",3315 => "10111001",3316 => "11101010",3317 => "00001100",3318 => "01010011",3319 => "00011110",3320 => "01101001",3321 => "00110010",3322 => "10110000",3323 => "10100000",3324 => "11110110",3325 => "01011100",3326 => "11000011",3327 => "00010000",3328 => "00101101",3329 => "11011011",3330 => "10100010",3331 => "00000000",3332 => "10111111",3333 => "00000001",3334 => "00111100",3335 => "00010110",3336 => "01111100",3337 => "11000110",3338 => "01011111",3339 => "10011110",3340 => "00001111",3341 => "00110001",3342 => "11100111",3343 => "01001010",3344 => "00101111",3345 => "00100111",3346 => "01110101",3347 => "10101000",3348 => "01011010",3349 => "01101110",3350 => "01101000",3351 => "00110011",3352 => "01111101",3353 => "11011001",3354 => "01110011",3355 => "01100000",3356 => "01110010",3357 => "11000110",3358 => "00000101",3359 => "11111110",3360 => "01011110",3361 => "00010111",3362 => "01010010",3363 => "01011111",3364 => "10010111",3365 => "10110011",3366 => "11010001",3367 => "10100010",3368 => "01000000",3369 => "00111101",3370 => "11101100",3371 => "00000100",3372 => "00011101",3373 => "11010011",3374 => "10101001",3375 => "10111110",3376 => "11100010",3377 => "11000001",3378 => "11000100",3379 => "01010101",3380 => "01010110",3381 => "00000111",3382 => "10101011",3383 => "10000011",3384 => "00000110",3385 => "11000000",3386 => "01011101",3387 => "10011000",3388 => "01010101",3389 => "11111101",3390 => "11101011",3391 => "11111011",3392 => "01010110",3393 => "00011111",3394 => "11101010",3395 => "11011001",3396 => "01010111",3397 => "00010100",3398 => "00110001",3399 => "11001001",3400 => "00100001",3401 => "10011110",3402 => "01001011",3403 => "01010101",3404 => "11011001",3405 => "01001010",3406 => "01011111",3407 => "10111111",3408 => "01001010",3409 => "10101111",3410 => "00101010",3411 => "01101001",3412 => "11010010",3413 => "01100000",3414 => "01111100",3415 => "11010001",3416 => "00111101",3417 => "11011010",3418 => "11011101",3419 => "10011111",3420 => "11101100",3421 => "10101101",3422 => "11101111",3423 => "10011001",3424 => "00000101",3425 => "01111001",3426 => "01001110",3427 => "01000011",3428 => "00000011",3429 => "11001001",3430 => "11101001",3431 => "01101101",3432 => "00011101",3433 => "11111001",3434 => "11011001",3435 => "10100101",3436 => "11001010",3437 => "00011001",3438 => "11011001",3439 => "01000000",3440 => "00100111",3441 => "11010000",3442 => "01000100",3443 => "01110111",3444 => "10111100",3445 => "00111011",3446 => "10010000",3447 => "11001001",3448 => "11101110",3449 => "00011000",3450 => "11001000",3451 => "10010000",3452 => "10111001",3453 => "00110101",3454 => "00100010",3455 => "10101011",3456 => "10001001",3457 => "11001001",3458 => "11010101",3459 => "01111010",3460 => "10000111",3461 => "00100011",3462 => "10111000",3463 => "10111101",3464 => "10011111",3465 => "10111101",3466 => "01011111",3467 => "10101110",3468 => "11101001",3469 => "01111010",3470 => "10001111",3471 => "10011110",3472 => "10111100",3473 => "00000100",3474 => "10111111",3475 => "10011011",3476 => "01101100",3477 => "10100001",3478 => "01111101",3479 => "00110011",3480 => "00001010",3481 => "11110111",3482 => "01101101",3483 => "10101000",3484 => "11010000",3485 => "11010010",3486 => "00110000",3487 => "10111010",3488 => "10100011",3489 => "10001010",3490 => "00101101",3491 => "10010000",3492 => "10101110",3493 => "01010001",3494 => "11100101",3495 => "10101001",3496 => "01100111",3497 => "10110111",3498 => "10000110",3499 => "00001101",3500 => "11001111",3501 => "11111000",3502 => "01000001",3503 => "00000101",3504 => "11100110",3505 => "10110000",3506 => "11001100",3507 => "10101101",3508 => "01101001",3509 => "10111101",3510 => "01011001",3511 => "11011000",3512 => "10010101",3513 => "00111111",3514 => "00100000",3515 => "11111110",3516 => "11001010",3517 => "00000001",3518 => "01010101",3519 => "10010011",3520 => "11110110",3521 => "11100011",3522 => "00001111",3523 => "11100110",3524 => "01010011",3525 => "01101000",3526 => "10100111",3527 => "01001110",3528 => "10001000",3529 => "01111101",3530 => "10101110",3531 => "01011101",3532 => "01000110",3533 => "01010111",3534 => "11110110",3535 => "00110010",3536 => "01010010",3537 => "10000001",3538 => "10001010",3539 => "11010000",3540 => "01000000",3541 => "00011110",3542 => "00011001",3543 => "11101011",3544 => "01011001",3545 => "01111100",3546 => "00000110",3547 => "10001101",3548 => "10110000",3549 => "00010101",3550 => "11100110",3551 => "01100000",3552 => "10010110",3553 => "01101111",3554 => "01011001",3555 => "10110110",3556 => "00011111",3557 => "01111010",3558 => "00110101",3559 => "00100110",3560 => "01111011",3561 => "10011000",3562 => "11011101",3563 => "10000001",3564 => "11010101",3565 => "10100111",3566 => "10110111",3567 => "10101110",3568 => "00001001",3569 => "11000010",3570 => "00010110",3571 => "00010011",3572 => "00010100",3573 => "01010101",3574 => "00000101",3575 => "11101100",3576 => "00011100",3577 => "01100001",3578 => "10100010",3579 => "10000101",3580 => "11001101",3581 => "11100111",3582 => "11100101",3583 => "11011100",3584 => "11000000",3585 => "11011111",3586 => "10110000",3587 => "10011111",3588 => "10010000",3589 => "00110010",3590 => "11000011",3591 => "10000011",3592 => "10100000",3593 => "00010111",3594 => "01101100",3595 => "10001010",3596 => "11001101",3597 => "10000011",3598 => "11010001",3599 => "01000111",3600 => "10011101",3601 => "10000010",3602 => "10011000",3603 => "11010110",3604 => "11100100",3605 => "00000001",3606 => "10100011",3607 => "11110011",3608 => "00011100",3609 => "10110101",3610 => "10110101",3611 => "10011101",3612 => "10011011",3613 => "11100100",3614 => "10000110",3615 => "00101001",3616 => "11001010",3617 => "11010010",3618 => "11001000",3619 => "00000100",3620 => "01110100",3621 => "00000101",3622 => "11111101",3623 => "11111000",3624 => "01101010",3625 => "10100101",3626 => "10000110",3627 => "01101000",3628 => "01111110",3629 => "10010011",3630 => "10100100",3631 => "11111010",3632 => "00111101",3633 => "00100100",3634 => "10100001",3635 => "01010011",3636 => "10011000",3637 => "11110100",3638 => "11000011",3639 => "01000101",3640 => "11110100",3641 => "11101001",3642 => "00101011",3643 => "00010111",3644 => "11111100",3645 => "10111110",3646 => "11001110",3647 => "00001001",3648 => "01100101",3649 => "00001100",3650 => "00101001",3651 => "11010111",3652 => "11011011",3653 => "11010100",3654 => "10000000",3655 => "00111010",3656 => "11010010",3657 => "11100000",3658 => "01101101",3659 => "01100011",3660 => "11010010",3661 => "01010101",3662 => "11100010",3663 => "00100100",3664 => "01110101",3665 => "01001100",3666 => "11101010",3667 => "11011101",3668 => "01101100",3669 => "01100111",3670 => "00001001",3671 => "10001111",3672 => "10000001",3673 => "00011000",3674 => "00001101",3675 => "01101100",3676 => "10101010",3677 => "10101110",3678 => "01100000",3679 => "11110110",3680 => "01001101",3681 => "10000011",3682 => "10001011",3683 => "01010010",3684 => "01101011",3685 => "10000101",3686 => "00110100",3687 => "01111110",3688 => "11000100",3689 => "00001000",3690 => "11101011",3691 => "00110011",3692 => "01100100",3693 => "11110100",3694 => "11011010",3695 => "00000011",3696 => "00111111",3697 => "01111110",3698 => "00000010",3699 => "01011111",3700 => "10010110",3701 => "11000010",3702 => "01101000",3703 => "01100001",3704 => "10100100",3705 => "11001111",3706 => "01110110",3707 => "10100111",3708 => "00011011",3709 => "11000011",3710 => "10101010",3711 => "01000101",3712 => "11110010",3713 => "01110000",3714 => "11100110",3715 => "10100011",3716 => "00010101",3717 => "10000001",3718 => "00010010",3719 => "10011110",3720 => "00101011",3721 => "10110001",3722 => "00000011",3723 => "01011110",3724 => "10010010",3725 => "01000101",3726 => "00100010",3727 => "00110010",3728 => "00011011",3729 => "01001101",3730 => "10010110",3731 => "10111011",3732 => "10010011",3733 => "00010001",3734 => "10110001",3735 => "10001000",3736 => "01000000",3737 => "11110101",3738 => "01100001",3739 => "00111011",3740 => "10011000",3741 => "00101000",3742 => "10000011",3743 => "00110100",3744 => "11101010",3745 => "11111010",3746 => "11011001",3747 => "01111111",3748 => "01100100",3749 => "01111100",3750 => "11110001",3751 => "11100101",3752 => "10001001",3753 => "11010100",3754 => "10101101",3755 => "01001010",3756 => "10011011",3757 => "00001111",3758 => "10010010",3759 => "11101110",3760 => "11101001",3761 => "00111110",3762 => "00011000",3763 => "11100011",3764 => "01000100",3765 => "11001000",3766 => "01000010",3767 => "10110111",3768 => "10001111",3769 => "00100001",3770 => "10100000",3771 => "01000100",3772 => "01000101",3773 => "00001100",3774 => "11011000",3775 => "01001011",3776 => "01111101",3777 => "00010011",3778 => "01100000",3779 => "10000000",3780 => "01101001",3781 => "01010011",3782 => "00111101",3783 => "11100100",3784 => "00110011",3785 => "11101001",3786 => "11110110",3787 => "10110000",3788 => "00110011",3789 => "01100100",3790 => "11000010",3791 => "11110011",3792 => "10000100",3793 => "00111000",3794 => "01111000",3795 => "11011111",3796 => "01001111",3797 => "11110101",3798 => "01110111",3799 => "10101111",3800 => "00101000",3801 => "00001001",3802 => "10010010",3803 => "11111101",3804 => "10100111",3805 => "01001011",3806 => "11101100",3807 => "11000011",3808 => "00111100",3809 => "10111000",3810 => "11010110",3811 => "11011010",3812 => "00001110",3813 => "11010010",3814 => "00000111",3815 => "01010001",3816 => "11001101",3817 => "11011000",3818 => "11101100",3819 => "00000000",3820 => "11101011",3821 => "01000000",3822 => "11111011",3823 => "01101101",3824 => "00001000",3825 => "00011011",3826 => "10100010",3827 => "00011111",3828 => "00001000",3829 => "10110100",3830 => "00100111",3831 => "00101110",3832 => "11000000",3833 => "10000100",3834 => "01011101",3835 => "10001001",3836 => "11100000",3837 => "01110001",3838 => "11001010",3839 => "11110010",3840 => "00001101",3841 => "11011100",3842 => "10010110",3843 => "11111000",3844 => "01010011",3845 => "10001001",3846 => "11110011",3847 => "00001100",3848 => "01000000",3849 => "11111000",3850 => "11011000",3851 => "01110110",3852 => "00110110",3853 => "11111110",3854 => "01111000",3855 => "10010111",3856 => "11000111",3857 => "11100010",3858 => "01000010",3859 => "10110100",3860 => "00100110",3861 => "10010100",3862 => "01010101",3863 => "10000001",3864 => "11101110",3865 => "10111101",3866 => "01000111",3867 => "01001011",3868 => "10011111",3869 => "11101011",3870 => "11110110",3871 => "01011000",3872 => "00111001",3873 => "01010001",3874 => "00101010",3875 => "11011010",3876 => "00101011",3877 => "11100111",3878 => "10101010",3879 => "10101000",3880 => "11110101",3881 => "00010110",3882 => "01100111",3883 => "10100100",3884 => "11110010",3885 => "10010010",3886 => "01011000",3887 => "01110010",3888 => "11010010",3889 => "01011011",3890 => "11110101",3891 => "11111011",3892 => "10010001",3893 => "00000001",3894 => "01001010",3895 => "01111100",3896 => "11000011",3897 => "00001111",3898 => "00110110",3899 => "10010001",3900 => "01000100",3901 => "10010011",3902 => "11000101",3903 => "11000101",3904 => "01011100",3905 => "01101000",3906 => "10000010",3907 => "00000111",3908 => "11001000",3909 => "10000010",3910 => "00100110",3911 => "11100010",3912 => "01010111",3913 => "10110111",3914 => "00111000",3915 => "01101101",3916 => "01001101",3917 => "10111111",3918 => "10111111",3919 => "10000110",3920 => "10000110",3921 => "11001110",3922 => "10110000",3923 => "11000101",3924 => "00101101",3925 => "00011010",3926 => "10001010",3927 => "00110010",3928 => "01111100",3929 => "10001001",3930 => "11101100",3931 => "00000101",3932 => "10000010",3933 => "01111110",3934 => "11000100",3935 => "11111011",3936 => "11100011",3937 => "11101011",3938 => "10100011",3939 => "11001110",3940 => "10011101",3941 => "00110111",3942 => "11100110",3943 => "00101110",3944 => "10001110",3945 => "01011001",3946 => "11001111",3947 => "01101000",3948 => "01000101",3949 => "00011111",3950 => "10100010",3951 => "10110101",3952 => "01010011",3953 => "01101100",3954 => "11011010",3955 => "11110100",3956 => "10111010",3957 => "11101101",3958 => "01101101",3959 => "00011101",3960 => "01101111",3961 => "01111001",3962 => "10111000",3963 => "11111000",3964 => "11000010",3965 => "00111000",3966 => "10100010",3967 => "10110011",3968 => "10001101",3969 => "10101111",3970 => "10000011",3971 => "10001111",3972 => "01010010",3973 => "10101010",3974 => "01101000",3975 => "00111110",3976 => "00011111",3977 => "00101111",3978 => "11100000",3979 => "11001010",3980 => "00110111",3981 => "10011100",3982 => "01000100",3983 => "11011001",3984 => "00010111",3985 => "10001100",3986 => "01010110",3987 => "00010000",3988 => "10001111",3989 => "11011110",3990 => "00101100",3991 => "10100100",3992 => "10011101",3993 => "01010010",3994 => "10010000",3995 => "11100101",3996 => "10000111",3997 => "01100010",3998 => "01111010",3999 => "00001100",4000 => "01000011",4001 => "00011111",4002 => "01001100",4003 => "01001100",4004 => "10101110",4005 => "00111001",4006 => "01000011",4007 => "00110011",4008 => "01000001",4009 => "00011100",4010 => "00111100",4011 => "01000000",4012 => "11001110",4013 => "11011000",4014 => "10110100",4015 => "01111010",4016 => "11000000",4017 => "10010010",4018 => "00011000",4019 => "10000010",4020 => "10000100",4021 => "11101110",4022 => "10011110",4023 => "00000001",4024 => "10111101",4025 => "10000111",4026 => "01100000",4027 => "11100001",4028 => "00110011",4029 => "11100011",4030 => "01010010",4031 => "10111001",4032 => "00110011",4033 => "10010010",4034 => "01111001",4035 => "10111000",4036 => "00001011",4037 => "00110110",4038 => "00001000",4039 => "00111000",4040 => "10001101",4041 => "01100111",4042 => "11010010",4043 => "01110010",4044 => "11000100",4045 => "10000111",4046 => "01110010",4047 => "00101001",4048 => "11011010",4049 => "10010100",4050 => "01101010",4051 => "10000100",4052 => "10000001",4053 => "11111101",4054 => "10110100",4055 => "00101001",4056 => "11110011",4057 => "00100110",4058 => "00111101",4059 => "00111101",4060 => "00011101",4061 => "11100011",4062 => "11011100",4063 => "01100011",4064 => "10010010",4065 => "11111100",4066 => "11011010",4067 => "00110111",4068 => "10001000",4069 => "01101111",4070 => "10111110",4071 => "10100100",4072 => "11011011",4073 => "10011101",4074 => "01001110",4075 => "00000101",4076 => "00111010",4077 => "01010100",4078 => "10000001",4079 => "01010101",4080 => "01000111",4081 => "11110001",4082 => "01111101",4083 => "00011111",4084 => "00001001",4085 => "00010110",4086 => "10011100",4087 => "01010011",4088 => "10100100",4089 => "01100100",4090 => "10011100",4091 => "11101100",4092 => "11011111",4093 => "00101101",4094 => "10000101",4095 => "01111101",4096 => "11110001",4097 => "11011000",4098 => "11110010",4099 => "01110010",4100 => "10111000",4101 => "00001001",4102 => "00111110",4103 => "00111011",4104 => "00010110",4105 => "01001011",4106 => "00010000",4107 => "00100111",4108 => "10010000",4109 => "10111111",4110 => "00110110",4111 => "01111001",4112 => "01100100",4113 => "01000010",4114 => "10100111",4115 => "00110101",4116 => "10011011",4117 => "11110001",4118 => "01111100",4119 => "00010011",4120 => "00111100",4121 => "01110001",4122 => "00101000",4123 => "11000101",4124 => "11001001",4125 => "11000001",4126 => "11111101",4127 => "01001001",4128 => "11101011",4129 => "10010001",4130 => "01001111",4131 => "00001011",4132 => "00000111",4133 => "00111011",4134 => "11110100",4135 => "10010011",4136 => "00100011",4137 => "10110110",4138 => "01101010",4139 => "01000000",4140 => "11010000",4141 => "10101011",4142 => "10101110",4143 => "01001111",4144 => "11000111",4145 => "00111000",4146 => "01001010",4147 => "10110010",4148 => "10010100",4149 => "11110000",4150 => "10101101",4151 => "10100011",4152 => "10001010",4153 => "00010000",4154 => "01001101",4155 => "01000010",4156 => "01111101",4157 => "10110111",4158 => "11101011",4159 => "11100110",4160 => "01010000",4161 => "01011111",4162 => "01011001",4163 => "10001001",4164 => "01110101",4165 => "11111011",4166 => "10111101",4167 => "00001011",4168 => "11000110",4169 => "10000000",4170 => "01101111",4171 => "00111100",4172 => "10110011",4173 => "01010101",4174 => "00101100",4175 => "11101010",4176 => "11001111",4177 => "01111010",4178 => "11110011",4179 => "01001100",4180 => "11100011",4181 => "11001101",4182 => "11111010",4183 => "00011111",4184 => "11110111",4185 => "10110000",4186 => "00010011",4187 => "01111100",4188 => "01010011",4189 => "10111110",4190 => "11011010",4191 => "10100001",4192 => "00100001",4193 => "01010011",4194 => "01011111",4195 => "11001111",4196 => "11010000",4197 => "01101100",4198 => "10001001",4199 => "11001110",4200 => "01010011",4201 => "00111011",4202 => "00000000",4203 => "10100010",4204 => "00101001",4205 => "11101001",4206 => "00010101",4207 => "01100001",4208 => "01101110",4209 => "00100101",4210 => "10110110",4211 => "01011111",4212 => "00010110",4213 => "11010100",4214 => "00001011",4215 => "00100101",4216 => "11110110",4217 => "11110010",4218 => "10110011",4219 => "01001111",4220 => "00110110",4221 => "11100010",4222 => "10010110",4223 => "11111110",4224 => "00011100",4225 => "10000101",4226 => "11011001",4227 => "01100111",4228 => "01110011",4229 => "10011110",4230 => "10101011",4231 => "10101101",4232 => "11100010",4233 => "11011001",4234 => "10101011",4235 => "11110111",4236 => "00101100",4237 => "11110111",4238 => "11001000",4239 => "11110111",4240 => "01111000",4241 => "00101100",4242 => "10011001",4243 => "01011000",4244 => "10111110",4245 => "00110110",4246 => "00000101",4247 => "11110100",4248 => "01101010",4249 => "00100000",4250 => "10110101",4251 => "01100000",4252 => "00011111",4253 => "00000011",4254 => "01000101",4255 => "11001011",4256 => "10000110",4257 => "01001101",4258 => "10100001",4259 => "11000110",4260 => "11001011",4261 => "01100011",4262 => "10101100",4263 => "10100101",4264 => "11110000",4265 => "11101001",4266 => "01101110",4267 => "10001010",4268 => "01011100",4269 => "01110111",4270 => "01111000",4271 => "11101000",4272 => "00100111",4273 => "10001001",4274 => "10111110",4275 => "10101110",4276 => "11010000",4277 => "11111010",4278 => "00111111",4279 => "10011010",4280 => "00010100",4281 => "01011110",4282 => "10000100",4283 => "00111111",4284 => "01010010",4285 => "11101110",4286 => "00101011",4287 => "10110111",4288 => "11100010",4289 => "11101101",4290 => "01011110",4291 => "00100110",4292 => "10111111",4293 => "10100011",4294 => "10011001",4295 => "10011101",4296 => "11100111",4297 => "01111011",4298 => "11010001",4299 => "10010001",4300 => "10000000",4301 => "10000011",4302 => "10001101",4303 => "10111011",4304 => "11100001",4305 => "10011011",4306 => "10011101",4307 => "11110111",4308 => "01010011",4309 => "11011011",4310 => "01110110",4311 => "00011011",4312 => "10110100",4313 => "01110011",4314 => "10111011",4315 => "01100101",4316 => "01110101",4317 => "00111110",4318 => "10000100",4319 => "10100000",4320 => "11100000",4321 => "11110100",4322 => "01100001",4323 => "00010000",4324 => "11100000",4325 => "00011000",4326 => "11011111",4327 => "11100110",4328 => "10010010",4329 => "00001100",4330 => "00010101",4331 => "00000000",4332 => "00010101",4333 => "01111111",4334 => "10111000",4335 => "01001100",4336 => "11010110",4337 => "10111101",4338 => "00001000",4339 => "11100100",4340 => "00100111",4341 => "01010100",4342 => "01010011",4343 => "11011101",4344 => "11010001",4345 => "11101100",4346 => "01101110",4347 => "11100101",4348 => "10111100",4349 => "01111100",4350 => "01011100",4351 => "11101001",4352 => "01101010",4353 => "00011100",4354 => "01011111",4355 => "00001100",4356 => "00101011",4357 => "00010101",4358 => "11011111",4359 => "00010100",4360 => "00110100",4361 => "00110000",4362 => "00100011",4363 => "01010010",4364 => "10101010",4365 => "11101100",4366 => "00100010",4367 => "01000010",4368 => "01001001",4369 => "11110000",4370 => "10011001",4371 => "10110100",4372 => "11111010",4373 => "10010000",4374 => "01010100",4375 => "01111101",4376 => "01011111",4377 => "01001101",4378 => "10000110",4379 => "01101100",4380 => "11001111",4381 => "00001001",4382 => "00010000",4383 => "00110110",4384 => "11101110",4385 => "00011110",4386 => "01111010",4387 => "01000010",4388 => "01111001",4389 => "01100001",4390 => "00010010",4391 => "00100001",4392 => "11001111",4393 => "10111010",4394 => "10001001",4395 => "10110001",4396 => "11000101",4397 => "01110010",4398 => "11011100",4399 => "10000001",4400 => "00011001",4401 => "00101001",4402 => "11110101",4403 => "10101011",4404 => "10101101",4405 => "01110010",4406 => "10100010",4407 => "10000010",4408 => "01010101",4409 => "00010101",4410 => "10001011",4411 => "00100000",4412 => "10001010",4413 => "01010001",4414 => "10000000",4415 => "01111001",4416 => "11001110",4417 => "01100110",4418 => "11100000",4419 => "01110111",4420 => "11011101",4421 => "11101111",4422 => "00110010",4423 => "10100110",4424 => "01011000",4425 => "11010101",4426 => "01111101",4427 => "11001101",4428 => "10011011",4429 => "01101001",4430 => "11011101",4431 => "10101001",4432 => "11010111",4433 => "01001011",4434 => "01001001",4435 => "00100011",4436 => "00101000",4437 => "01001010",4438 => "01110100",4439 => "11101011",4440 => "10101111",4441 => "11000000",4442 => "10001110",4443 => "10010110",4444 => "11110010",4445 => "10110101",4446 => "10111011",4447 => "00100001",4448 => "10101011",4449 => "11001010",4450 => "00011011",4451 => "00011111",4452 => "00110111",4453 => "10110101",4454 => "10100110",4455 => "11011001",4456 => "10010010",4457 => "01000100",4458 => "11000110",4459 => "01101001",4460 => "01000110",4461 => "01100100",4462 => "11110111",4463 => "01111010",4464 => "11101100",4465 => "00011101",4466 => "11101101",4467 => "11110000",4468 => "11110000",4469 => "10010101",4470 => "01111110",4471 => "10110010",4472 => "00001100",4473 => "10000000",4474 => "11010100",4475 => "00101110",4476 => "11010110",4477 => "11011110",4478 => "01101100",4479 => "01110101",4480 => "00011010",4481 => "10010110",4482 => "01001101",4483 => "00011000",4484 => "01101010",4485 => "11101001",4486 => "11111000",4487 => "10010010",4488 => "11001100",4489 => "01001010",4490 => "10100100",4491 => "11000100",4492 => "01111111",4493 => "01111100",4494 => "00100001",4495 => "00000000",4496 => "01111010",4497 => "11100011",4498 => "00000101",4499 => "00001011",4500 => "00010110",4501 => "11010100",4502 => "10001110",4503 => "10010111",4504 => "10100000",4505 => "01010010",4506 => "00011100",4507 => "00110111",4508 => "10100011",4509 => "11101000",4510 => "00001111",4511 => "11011001",4512 => "01111101",4513 => "11100111",4514 => "10001110",4515 => "01011001",4516 => "01000110",4517 => "00001011",4518 => "10010110",4519 => "01011000",4520 => "11111010",4521 => "01110010",4522 => "01100101",4523 => "00110110",4524 => "11001100",4525 => "10000001",4526 => "10110010",4527 => "10100001",4528 => "00111010",4529 => "11000111",4530 => "10001001",4531 => "10010000",4532 => "00111011",4533 => "01100111",4534 => "00010111",4535 => "00001101",4536 => "00110010",4537 => "11111011",4538 => "01100001",4539 => "10101011",4540 => "11011010",4541 => "01010010",4542 => "01010000",4543 => "00111011",4544 => "11111101",4545 => "11011100",4546 => "01110100",4547 => "00101000",4548 => "11011100",4549 => "10110011",4550 => "10101011",4551 => "10101111",4552 => "00010001",4553 => "01001000",4554 => "00100000",4555 => "01011001",4556 => "11010101",4557 => "01011010",4558 => "00111010",4559 => "00101010",4560 => "00110000",4561 => "11111110",4562 => "11101111",4563 => "10001101",4564 => "11101111",4565 => "01100100",4566 => "00010001",4567 => "01000010",4568 => "10100110",4569 => "11000001",4570 => "01000010",4571 => "10010000",4572 => "00100011",4573 => "01001001",4574 => "00110101",4575 => "11100001",4576 => "10101101",4577 => "00001000",4578 => "00111010",4579 => "10001111",4580 => "00110100",4581 => "01111100",4582 => "10101011",4583 => "10101110",4584 => "10011011",4585 => "10110011",4586 => "00000101",4587 => "10000101",4588 => "01011111",4589 => "10101101",4590 => "11010000",4591 => "00101010",4592 => "11110010",4593 => "01110110",4594 => "11110010",4595 => "00001001",4596 => "10001000",4597 => "01000010",4598 => "01001010",4599 => "00100010",4600 => "10110001",4601 => "01110111",4602 => "10000001",4603 => "01100001",4604 => "11010111",4605 => "00010000",4606 => "11011001",4607 => "00010000",4608 => "01000001",4609 => "11011011",4610 => "10000110",4611 => "11011110",4612 => "00011010",4613 => "01010111",4614 => "00101010",4615 => "01001001",4616 => "11000101",4617 => "11101011",4618 => "11011001",4619 => "01101110",4620 => "10100100",4621 => "11000010",4622 => "00000001",4623 => "11100010",4624 => "11111101",4625 => "00100010",4626 => "01000111",4627 => "10001010",4628 => "01011011",4629 => "11001101",4630 => "00011101",4631 => "10111111",4632 => "00100000",4633 => "00011011",4634 => "01101000",4635 => "11101000",4636 => "00011000",4637 => "10111100",4638 => "00011000",4639 => "11101100",4640 => "01111111",4641 => "11000000",4642 => "00010010",4643 => "10111011",4644 => "10111110",4645 => "11010101",4646 => "11100001",4647 => "01111100",4648 => "10101101",4649 => "11111110",4650 => "01111111",4651 => "10001011",4652 => "00110001",4653 => "11010000",4654 => "10110010",4655 => "11110001",4656 => "00001101",4657 => "01111000",4658 => "11010110",4659 => "00110100",4660 => "01011101",4661 => "10010010",4662 => "10000011",4663 => "01110101",4664 => "10010011",4665 => "10010110",4666 => "01111111",4667 => "10000011",4668 => "10011100",4669 => "01001110",4670 => "11011100",4671 => "10100100",4672 => "00011010",4673 => "10011001",4674 => "11000101",4675 => "01100111",4676 => "01100001",4677 => "10111010",4678 => "01010010",4679 => "11110101",4680 => "01010000",4681 => "01100110",4682 => "00010100",4683 => "10101101",4684 => "10001000",4685 => "10111101",4686 => "01111000",4687 => "01010000",4688 => "10011000",4689 => "11001000",4690 => "11000011",4691 => "11010000",4692 => "10110101",4693 => "11001010",4694 => "01011111",4695 => "01000011",4696 => "10111101",4697 => "11011011",4698 => "00001000",4699 => "10101010",4700 => "10110101",4701 => "01101010",4702 => "10111111",4703 => "01111100",4704 => "11111100",4705 => "10101011",4706 => "01111011",4707 => "10101000",4708 => "10100111",4709 => "00011110",4710 => "01011110",4711 => "11110101",4712 => "10010010",4713 => "01110111",4714 => "10010101",4715 => "10111010",4716 => "10011100",4717 => "10011010",4718 => "00001100",4719 => "10010000",4720 => "00001101",4721 => "10101101",4722 => "00011011",4723 => "10001001",4724 => "11101001",4725 => "11010100",4726 => "00000100",4727 => "00110001",4728 => "10110011",4729 => "01110101",4730 => "11001010",4731 => "11101000",4732 => "11001110",4733 => "01001111",4734 => "00010000",4735 => "00101001",4736 => "01101001",4737 => "11100001",4738 => "01000111",4739 => "10111110",4740 => "10100010",4741 => "01010011",4742 => "10101110",4743 => "01001100",4744 => "10010000",4745 => "10101100",4746 => "01001000",4747 => "11000000",4748 => "01110000",4749 => "11010011",4750 => "00110011",4751 => "11100001",4752 => "11101101",4753 => "01010000",4754 => "10000010",4755 => "01101100",4756 => "00010010",4757 => "00110110",4758 => "10111111",4759 => "01001001",4760 => "11001000",4761 => "00010010",4762 => "11001001",4763 => "11111111",4764 => "01100011",4765 => "11011111",4766 => "00101011",4767 => "10101010",4768 => "01011101",4769 => "00110011",4770 => "10101001",4771 => "01110101",4772 => "01100110",4773 => "11001111",4774 => "11001011",4775 => "11101001",4776 => "11001000",4777 => "01010100",4778 => "10100111",4779 => "11111011",4780 => "11001001",4781 => "01011010",4782 => "10000111",4783 => "11001101",4784 => "00001101",4785 => "11100110",4786 => "10111110",4787 => "11110110",4788 => "01000111",4789 => "10011011",4790 => "10101110",4791 => "11001011",4792 => "10010101",4793 => "00100011",4794 => "01011101",4795 => "10100101",4796 => "01111111",4797 => "00001001",4798 => "00100111",4799 => "10011010",4800 => "10101011",4801 => "11000011",4802 => "01100100",4803 => "11100011",4804 => "10001101",4805 => "00000100",4806 => "10001010",4807 => "00001110",4808 => "00110000",4809 => "11111010",4810 => "01101110",4811 => "01010110",4812 => "00011001",4813 => "10101001",4814 => "11111111",4815 => "00000001",4816 => "11001110",4817 => "00100111",4818 => "10001000",4819 => "10000010",4820 => "00000001",4821 => "11101100",4822 => "11010111",4823 => "11100101",4824 => "11100111",4825 => "11111101",4826 => "00011111",4827 => "11111101",4828 => "10111100",4829 => "10000110",4830 => "00110000",4831 => "01011100",4832 => "00100011",4833 => "10011000",4834 => "10011000",4835 => "11101111",4836 => "01010000",4837 => "10000010",4838 => "11111011",4839 => "11100010",4840 => "10011101",4841 => "10010010",4842 => "10001111",4843 => "01111110",4844 => "01011010",4845 => "11001100",4846 => "10010001",4847 => "10011110",4848 => "01011100",4849 => "10010000",4850 => "11010100",4851 => "10001101",4852 => "00001000",4853 => "00101101",4854 => "11100100",4855 => "10110011",4856 => "00011011",4857 => "00011110",4858 => "10101101",4859 => "00011111",4860 => "11010011",4861 => "01000011",4862 => "10101000",4863 => "11000010",4864 => "01110000",4865 => "01111010",4866 => "11000101",4867 => "10010010",4868 => "01111000",4869 => "10011000",4870 => "00101010",4871 => "01100100",4872 => "01000100",4873 => "10110001",4874 => "11100100",4875 => "10000001",4876 => "01101111",4877 => "01000011",4878 => "00100101",4879 => "01110001",4880 => "10011110",4881 => "11101001",4882 => "01000000",4883 => "10100100",4884 => "00110011",4885 => "11011110",4886 => "10010001",4887 => "10111001",4888 => "10010010",4889 => "01101010",4890 => "01011110",4891 => "00011111",4892 => "00010100",4893 => "01110101",4894 => "10010001",4895 => "10110100",4896 => "11101101",4897 => "11001010",4898 => "11000111",4899 => "00110011",4900 => "10100111",4901 => "00011011",4902 => "00000110",4903 => "10100110",4904 => "10101000",4905 => "11000101",4906 => "10110010",4907 => "10111000",4908 => "00011110",4909 => "01100011",4910 => "01010001",4911 => "11111011",4912 => "11111111",4913 => "10001010",4914 => "11110101",4915 => "01000111",4916 => "11010010",4917 => "10111111",4918 => "01101000",4919 => "11101110",4920 => "11000001",4921 => "11110010",4922 => "11100100",4923 => "00100101",4924 => "10001001",4925 => "01000101",4926 => "01010011",4927 => "01001100",4928 => "11100110",4929 => "11110100",4930 => "00110001",4931 => "11000011",4932 => "11100001",4933 => "00000000",4934 => "00011111",4935 => "00111101",4936 => "01011101",4937 => "11000000",4938 => "00110001",4939 => "01010001",4940 => "00100100",4941 => "01001101",4942 => "11010111",4943 => "10101101",4944 => "11111011",4945 => "01001000",4946 => "11000001",4947 => "01000101",4948 => "10100111",4949 => "01011000",4950 => "11100011",4951 => "11110110",4952 => "10100101",4953 => "01111110",4954 => "11111001",4955 => "10001000",4956 => "10001111",4957 => "01101101",4958 => "10001000",4959 => "01101000",4960 => "10111110",4961 => "10110001",4962 => "11110000",4963 => "00011000",4964 => "01111000",4965 => "00000001",4966 => "11000001",4967 => "10000011",4968 => "00111001",4969 => "00010111",4970 => "00101101",4971 => "01100111",4972 => "11110111",4973 => "01010101",4974 => "00001111",4975 => "01010010",4976 => "10101011",4977 => "01000111",4978 => "10010101",4979 => "11000101",4980 => "01101111",4981 => "01111001",4982 => "10000100",4983 => "11010010",4984 => "00111000",4985 => "10110101",4986 => "11110110",4987 => "01000011",4988 => "00101100",4989 => "00001011",4990 => "00101110",4991 => "01000110",4992 => "00110001",4993 => "00101101",4994 => "10100000",4995 => "01100010",4996 => "10011101",4997 => "10101000",4998 => "01100011",4999 => "00111101",5000 => "00100101",5001 => "01000011",5002 => "11011010",5003 => "01010001",5004 => "11000111",5005 => "01000110",5006 => "11100010",5007 => "00001000",5008 => "10011100",5009 => "11110101",5010 => "00111100",5011 => "01011001",5012 => "01000111",5013 => "11111101",5014 => "00000011",5015 => "01101010",5016 => "11011101",5017 => "11100111",5018 => "01100111",5019 => "01100100",5020 => "10100000",5021 => "00010110",5022 => "01101100",5023 => "00101000",5024 => "00001110",5025 => "01100111",5026 => "10110111",5027 => "01101100",5028 => "10000111",5029 => "01111100",5030 => "01010111",5031 => "01010001",5032 => "01100010",5033 => "11011001",5034 => "11001011",5035 => "11111011",5036 => "10101001",5037 => "11110010",5038 => "11000111",5039 => "11011111",5040 => "11000111",5041 => "00011100",5042 => "00100010",5043 => "10100100",5044 => "00001001",5045 => "01110000",5046 => "01101100",5047 => "00000010",5048 => "01000110",5049 => "11101110",5050 => "01011001",5051 => "11001000",5052 => "11000011",5053 => "11110000",5054 => "00001100",5055 => "00011000",5056 => "10010111",5057 => "10010000",5058 => "01110011",5059 => "00011101",5060 => "10110010",5061 => "00111001",5062 => "10000110",5063 => "11001001",5064 => "00110001",5065 => "11010000",5066 => "10101011",5067 => "00001110",5068 => "00101000",5069 => "10110010",5070 => "11101111",5071 => "10010111",5072 => "00111111",5073 => "11101100",5074 => "01010100",5075 => "11001001",5076 => "11001100",5077 => "01010100",5078 => "10001001",5079 => "11101001",5080 => "10011101",5081 => "10110001",5082 => "00011111",5083 => "11000100",5084 => "00000101",5085 => "11010010",5086 => "11111111",5087 => "11011000",5088 => "11011101",5089 => "00100110",5090 => "10101101",5091 => "00010011",5092 => "01110011",5093 => "11000111",5094 => "00110100",5095 => "00011101",5096 => "10000111",5097 => "00000010",5098 => "10110011",5099 => "00110111",5100 => "00100111",5101 => "01011011",5102 => "10101010",5103 => "10110011",5104 => "00011101",5105 => "01001011",5106 => "00010100",5107 => "00001000",5108 => "11010110",5109 => "11111101",5110 => "01101011",5111 => "10000111",5112 => "01001000",5113 => "01011101",5114 => "11011011",5115 => "11001110",5116 => "00001100",5117 => "11101001",5118 => "00001000",5119 => "10011001",5120 => "10111110",5121 => "00010110",5122 => "10110000",5123 => "01001101",5124 => "00101110",5125 => "10111100",5126 => "10011110",5127 => "11011011",5128 => "00010100",5129 => "10000001",5130 => "11001111",5131 => "10110111",5132 => "01111011",5133 => "01000111",5134 => "00101010",5135 => "00110101",5136 => "11110000",5137 => "01011011",5138 => "01000110",5139 => "00001000",5140 => "11111110",5141 => "11001101",5142 => "11100100",5143 => "11010000",5144 => "01010001",5145 => "01011000",5146 => "00001000",5147 => "11100101",5148 => "10101011",5149 => "10011101",5150 => "00011110",5151 => "00101010",5152 => "00100100",5153 => "11011101",5154 => "01011101",5155 => "00111011",5156 => "00000100",5157 => "01110111",5158 => "11011110",5159 => "11010101",5160 => "10100111",5161 => "01011000",5162 => "00010111",5163 => "01101000",5164 => "00100111",5165 => "01000110",5166 => "11001111",5167 => "10100111",5168 => "01100101",5169 => "11100011",5170 => "00011001",5171 => "10110010",5172 => "00000000",5173 => "10010110",5174 => "10000001",5175 => "01110010",5176 => "11010010",5177 => "01100011",5178 => "11101111",5179 => "00001001",5180 => "01001111",5181 => "10101001",5182 => "10110100",5183 => "00111010",5184 => "00100111",5185 => "01001110",5186 => "10011101",5187 => "10001010",5188 => "01101110",5189 => "11011101",5190 => "00101111",5191 => "11000010",5192 => "01100100",5193 => "10011110",5194 => "00100001",5195 => "11001110",5196 => "01010000",5197 => "01100111",5198 => "10100110",5199 => "11010111",5200 => "11100011",5201 => "01101111",5202 => "01101111",5203 => "01100011",5204 => "01101111",5205 => "10001110",5206 => "11111010",5207 => "01001011",5208 => "01001100",5209 => "11000111",5210 => "00001101",5211 => "00100010",5212 => "01100100",5213 => "11111101",5214 => "11000001",5215 => "11011000",5216 => "10010011",5217 => "00010011",5218 => "01100010",5219 => "01001111",5220 => "00010101",5221 => "10010000",5222 => "10011001",5223 => "10100000",5224 => "00111001",5225 => "01110110",5226 => "10011110",5227 => "11000000",5228 => "11110010",5229 => "11100011",5230 => "01000010",5231 => "10001011",5232 => "01000110",5233 => "00110000",5234 => "01001100",5235 => "10111011",5236 => "01101010",5237 => "00001110",5238 => "00001011",5239 => "10100111",5240 => "10000111",5241 => "10001010",5242 => "11010010",5243 => "11000000",5244 => "01000001",5245 => "00000101",5246 => "01110101",5247 => "01001000",5248 => "11010001",5249 => "01100000",5250 => "11111100",5251 => "10001101",5252 => "00101011",5253 => "00000011",5254 => "01101101",5255 => "11011111",5256 => "11000111",5257 => "11001000",5258 => "10010001",5259 => "00001110",5260 => "01111000",5261 => "00000100",5262 => "11010001",5263 => "10011001",5264 => "00100000",5265 => "11110000",5266 => "10100111",5267 => "10110101",5268 => "10000010",5269 => "00000011",5270 => "01001101",5271 => "00111101",5272 => "10111111",5273 => "10001101",5274 => "01111101",5275 => "10010011",5276 => "00011100",5277 => "01000101",5278 => "11011111",5279 => "01010110",5280 => "10111100",5281 => "10111000",5282 => "11111101",5283 => "00101011",5284 => "10010001",5285 => "10001111",5286 => "00111010",5287 => "00100110",5288 => "01010111",5289 => "01110100",5290 => "01110100",5291 => "10011000",5292 => "11011010",5293 => "11111010",5294 => "11100010",5295 => "11000011",5296 => "01001011",5297 => "01000010",5298 => "11100111",5299 => "11111110",5300 => "10011100",5301 => "11100000",5302 => "00010111",5303 => "01000100",5304 => "10011111",5305 => "01111000",5306 => "00100101",5307 => "10110100",5308 => "00001101",5309 => "10011000",5310 => "00010111",5311 => "11110000",5312 => "00011011",5313 => "10000111",5314 => "00000101",5315 => "10011000",5316 => "01010100",5317 => "01110110",5318 => "10101000",5319 => "10110001",5320 => "10110110",5321 => "00111000",5322 => "10110010",5323 => "11010101",5324 => "11001010",5325 => "01001010",5326 => "00110010",5327 => "11111010",5328 => "11011001",5329 => "00110101",5330 => "01001001",5331 => "01001010",5332 => "11001010",5333 => "10010010",5334 => "10000001",5335 => "01001101",5336 => "01110110",5337 => "10111010",5338 => "10001000",5339 => "00010110",5340 => "00101000",5341 => "00001100",5342 => "10100000",5343 => "01101001",5344 => "01111011",5345 => "00111011",5346 => "00001011",5347 => "01100001",5348 => "01001001",5349 => "10011010",5350 => "00110110",5351 => "00110010",5352 => "00010010",5353 => "11110001",5354 => "10000111",5355 => "10010111",5356 => "10101001",5357 => "01010111",5358 => "01011011",5359 => "11110110",5360 => "11111111",5361 => "01010110",5362 => "11111011",5363 => "00100100",5364 => "00000001",5365 => "00111101",5366 => "01100110",5367 => "00101100",5368 => "10100111",5369 => "00101000",5370 => "11111010",5371 => "00110100",5372 => "00010110",5373 => "10101001",5374 => "11010110",5375 => "11000001",5376 => "11101010",5377 => "10110010",5378 => "01101111",5379 => "01110100",5380 => "10110111",5381 => "01100100",5382 => "10100101",5383 => "11111011",5384 => "00011010",5385 => "11001110",5386 => "00010000",5387 => "00100011",5388 => "01101001",5389 => "10100001",5390 => "01001110",5391 => "10000011",5392 => "01011011",5393 => "00000001",5394 => "11011100",5395 => "01111010",5396 => "01000000",5397 => "01011010",5398 => "00011001",5399 => "10001001",5400 => "00000010",5401 => "10001010",5402 => "01001010",5403 => "01011001",5404 => "01111111",5405 => "00010011",5406 => "01110100",5407 => "10111000",5408 => "00100010",5409 => "10110000",5410 => "01001100",5411 => "11100101",5412 => "00001110",5413 => "01011101",5414 => "10110000",5415 => "10011111",5416 => "11000111",5417 => "01111011",5418 => "01010001",5419 => "11101100",5420 => "01100000",5421 => "11010001",5422 => "10011011",5423 => "11100111",5424 => "10111001",5425 => "10111111",5426 => "11111110",5427 => "10110000",5428 => "11110111",5429 => "00110101",5430 => "01011011",5431 => "10111101",5432 => "10010001",5433 => "11000101",5434 => "01101011",5435 => "11001001",5436 => "10100010",5437 => "00111000",5438 => "10001010",5439 => "11100110",5440 => "00001101",5441 => "00001110",5442 => "01111101",5443 => "10101110",5444 => "10010110",5445 => "01010100",5446 => "11100001",5447 => "00111111",5448 => "00010100",5449 => "11100110",5450 => "11100111",5451 => "01111000",5452 => "01110000",5453 => "11110101",5454 => "10000101",5455 => "10111100",5456 => "11111111",5457 => "01100101",5458 => "11010000",5459 => "10110101",5460 => "11011111",5461 => "01011100",5462 => "11001111",5463 => "01010011",5464 => "10000000",5465 => "00110100",5466 => "01111001",5467 => "00001001",5468 => "10111011",5469 => "01011010",5470 => "01110101",5471 => "10110001",5472 => "01110110",5473 => "10010110",5474 => "01100110",5475 => "01101101",5476 => "01001111",5477 => "10111100",5478 => "10010011",5479 => "10101111",5480 => "00101100",5481 => "10110110",5482 => "01110101",5483 => "11000101",5484 => "10111100",5485 => "10010001",5486 => "10110010",5487 => "01111100",5488 => "01100111",5489 => "11000101",5490 => "00100110",5491 => "10100001",5492 => "01010000",5493 => "01101011",5494 => "10010001",5495 => "01110000",5496 => "01000111",5497 => "01100001",5498 => "01101110",5499 => "01100111",5500 => "10110101",5501 => "10110111",5502 => "01110110",5503 => "01010000",5504 => "00110110",5505 => "00001001",5506 => "00101100",5507 => "11100101",5508 => "01101111",5509 => "11010011",5510 => "10000100",5511 => "11001000",5512 => "00001001",5513 => "00100000",5514 => "10101000",5515 => "11000100",5516 => "00011011",5517 => "11101111",5518 => "00111100",5519 => "11110101",5520 => "01000111",5521 => "01010111",5522 => "00010111",5523 => "00110101",5524 => "10110100",5525 => "11110110",5526 => "11010100",5527 => "01100100",5528 => "10000101",5529 => "00110010",5530 => "10100010",5531 => "10010001",5532 => "10100010",5533 => "11110011",5534 => "00100111",5535 => "00010011",5536 => "01111111",5537 => "10100111",5538 => "00010010",5539 => "10110100",5540 => "00101101",5541 => "10101101",5542 => "00000001",5543 => "11011010",5544 => "01101111",5545 => "10000101",5546 => "00000001",5547 => "01100100",5548 => "11110000",5549 => "10010001",5550 => "11101100",5551 => "01001011",5552 => "11010101",5553 => "01010001",5554 => "11000111",5555 => "00010111",5556 => "10100011",5557 => "00111100",5558 => "00001111",5559 => "00100001",5560 => "01000101",5561 => "00010101",5562 => "00011011",5563 => "01001101",5564 => "00001111",5565 => "10011001",5566 => "10010100",5567 => "11001011",5568 => "11111111",5569 => "11110011",5570 => "01000100",5571 => "01000000",5572 => "00010100",5573 => "00001000",5574 => "00011110",5575 => "11000000",5576 => "11010101",5577 => "10000010",5578 => "01110110",5579 => "11111110",5580 => "00011101",5581 => "10111110",5582 => "10111001",5583 => "10001010",5584 => "00011111",5585 => "00101001",5586 => "11111011",5587 => "11000011",5588 => "11101010",5589 => "00100010",5590 => "00000010",5591 => "00010011",5592 => "11010110",5593 => "11100111",5594 => "01111011",5595 => "01001111",5596 => "01011001",5597 => "00110010",5598 => "10011111",5599 => "10010101",5600 => "11000111",5601 => "10001010",5602 => "00101001",5603 => "01100111",5604 => "01010001",5605 => "10011100",5606 => "00001100",5607 => "10011101",5608 => "11100010",5609 => "10001001",5610 => "01011011",5611 => "10100011",5612 => "10100110",5613 => "11110100",5614 => "10001011",5615 => "00111101",5616 => "00010110",5617 => "00110111",5618 => "01111110",5619 => "01010001",5620 => "01110011",5621 => "11110110",5622 => "00100010",5623 => "00101110",5624 => "10111001",5625 => "01100000",5626 => "00110110",5627 => "01100100",5628 => "11100000",5629 => "01010111",5630 => "10000011",5631 => "10001100",5632 => "00101100",5633 => "11010011",5634 => "01101010",5635 => "00110010",5636 => "10001111",5637 => "10001001",5638 => "01000110",5639 => "11011011",5640 => "11000110",5641 => "00001000",5642 => "10101001",5643 => "00100111",5644 => "10111100",5645 => "11011100",5646 => "01101001",5647 => "10001010",5648 => "10001110",5649 => "01100011",5650 => "01111100",5651 => "10111011",5652 => "01010010",5653 => "11001010",5654 => "00001111",5655 => "11110111",5656 => "10110110",5657 => "00111011",5658 => "01001010",5659 => "01111101",5660 => "11111101",5661 => "10010011",5662 => "01011000",5663 => "00101100",5664 => "10000110",5665 => "01101100",5666 => "01100110",5667 => "11101000",5668 => "01001011",5669 => "01111000",5670 => "00110111",5671 => "10100011",5672 => "00101100",5673 => "01010100",5674 => "00001010",5675 => "11111101",5676 => "11000011",5677 => "01110001",5678 => "01101001",5679 => "11001010",5680 => "11110100",5681 => "11111011",5682 => "00011101",5683 => "10101001",5684 => "01001110",5685 => "10101101",5686 => "00110111",5687 => "01011000",5688 => "10111010",5689 => "01111001",5690 => "11001011",5691 => "11101010",5692 => "11100001",5693 => "10001101",5694 => "01101101",5695 => "11110101",5696 => "00000101",5697 => "11010011",5698 => "00000011",5699 => "11000001",5700 => "00111101",5701 => "10111000",5702 => "01111000",5703 => "11010110",5704 => "01010011",5705 => "11111110",5706 => "11101111",5707 => "10000010",5708 => "01001110",5709 => "10111100",5710 => "00001100",5711 => "00011101",5712 => "00001101",5713 => "10000011",5714 => "01100000",5715 => "10001001",5716 => "01101001",5717 => "00100110",5718 => "10011011",5719 => "10101100",5720 => "10101000",5721 => "11001100",5722 => "00011011",5723 => "10011101",5724 => "00000000",5725 => "01001100",5726 => "01111010",5727 => "11000010",5728 => "01000010",5729 => "11010001",5730 => "10000001",5731 => "11100110",5732 => "10101110",5733 => "00101111",5734 => "10011000",5735 => "01101010",5736 => "11101001",5737 => "10001001",5738 => "11010110",5739 => "00110111",5740 => "10101001",5741 => "00001010",5742 => "10111111",5743 => "10011011",5744 => "10000001",5745 => "11100110",5746 => "00000100",5747 => "00101001",5748 => "11111001",5749 => "11011110",5750 => "01011101",5751 => "10000111",5752 => "10011001",5753 => "01001011",5754 => "10000101",5755 => "10110001",5756 => "10110001",5757 => "01001100",5758 => "01001011",5759 => "11000100",5760 => "00111010",5761 => "11110111",5762 => "10110010",5763 => "00011010",5764 => "00100100",5765 => "00000000",5766 => "10111010",5767 => "00011101",5768 => "00000010",5769 => "01001010",5770 => "11010001",5771 => "01000000",5772 => "00110010",5773 => "11010011",5774 => "00001011",5775 => "10011001",5776 => "11111100",5777 => "10101001",5778 => "01100011",5779 => "10101000",5780 => "11000110",5781 => "00100101",5782 => "00011011",5783 => "10000111",5784 => "00011000",5785 => "11011000",5786 => "11010000",5787 => "11001111",5788 => "10000101",5789 => "01001000",5790 => "00011101",5791 => "00001001",5792 => "11111001",5793 => "11010111",5794 => "01101100",5795 => "00001110",5796 => "01110110",5797 => "10110001",5798 => "10000000",5799 => "00000110",5800 => "00101001",5801 => "11111010",5802 => "01100011",5803 => "01110111",5804 => "01001011",5805 => "10000100",5806 => "01010100",5807 => "00101010",5808 => "11000001",5809 => "11111100",5810 => "11101001",5811 => "00101010",5812 => "01001000",5813 => "10110110",5814 => "01111010",5815 => "11101101",5816 => "11111001",5817 => "01111011",5818 => "10111111",5819 => "01011000",5820 => "01101100",5821 => "01111010",5822 => "11100011",5823 => "11110010",5824 => "10111110",5825 => "11011000",5826 => "01011001",5827 => "10001011",5828 => "11101101",5829 => "11011011",5830 => "11011011",5831 => "11100101",5832 => "00001011",5833 => "01101010",5834 => "01110111",5835 => "00111000",5836 => "00110010",5837 => "01001101",5838 => "10011000",5839 => "01011000",5840 => "11110100",5841 => "01100100",5842 => "10001101",5843 => "00101010",5844 => "11110000",5845 => "11110111",5846 => "10110001",5847 => "10001000",5848 => "11110011",5849 => "10110111",5850 => "11100001",5851 => "01001110",5852 => "00111101",5853 => "10010011",5854 => "10001100",5855 => "10001000",5856 => "11001011",5857 => "01111001",5858 => "10100001",5859 => "11001100",5860 => "11000110",5861 => "01100110",5862 => "10011110",5863 => "11011100",5864 => "01111111",5865 => "00011000",5866 => "00010000",5867 => "00100001",5868 => "10100111",5869 => "01100011",5870 => "01111001",5871 => "01100110",5872 => "00000000",5873 => "01101111",5874 => "01110011",5875 => "01001001",5876 => "00011110",5877 => "00000010",5878 => "01000110",5879 => "10000100",5880 => "00111101",5881 => "10101101",5882 => "10000011",5883 => "11010011",5884 => "00110101",5885 => "01011000",5886 => "00110010",5887 => "00100011",5888 => "01000110",5889 => "00000111",5890 => "11101100",5891 => "00110000",5892 => "11100110",5893 => "01101101",5894 => "01111010",5895 => "01000111",5896 => "10110101",5897 => "00011101",5898 => "10010110",5899 => "00100010",5900 => "00011011",5901 => "01100000",5902 => "01100101",5903 => "10111010",5904 => "10101101",5905 => "01110101",5906 => "11110010",5907 => "00011001",5908 => "11110010",5909 => "00110011",5910 => "10111010",5911 => "11001101",5912 => "01011110",5913 => "01000001",5914 => "11010000",5915 => "11110010",5916 => "10100010",5917 => "10011001",5918 => "00011000",5919 => "10001110",5920 => "01110001",5921 => "10011000",5922 => "01101110",5923 => "11101001",5924 => "11101001",5925 => "00001101",5926 => "01001110",5927 => "11110100",5928 => "01011000",5929 => "00001101",5930 => "11110001",5931 => "00000100",5932 => "10010110",5933 => "11100101",5934 => "10010011",5935 => "10011010",5936 => "10010101",5937 => "10110011",5938 => "10100001",5939 => "10010001",5940 => "01010001",5941 => "00010101",5942 => "00011111",5943 => "01110011",5944 => "01111011",5945 => "01110011",5946 => "11110010",5947 => "10000010",5948 => "10011010",5949 => "01010111",5950 => "01000010",5951 => "11001100",5952 => "00000011",5953 => "10011010",5954 => "00010000",5955 => "00011100",5956 => "11111100",5957 => "11011011",5958 => "10100011",5959 => "10010101",5960 => "00100110",5961 => "11011000",5962 => "00001101",5963 => "11111101",5964 => "10011100",5965 => "01101010",5966 => "00001111",5967 => "00001100",5968 => "01101111",5969 => "10011011",5970 => "10010110",5971 => "11101000",5972 => "10110110",5973 => "10001011",5974 => "11000011",5975 => "10011001",5976 => "00001000",5977 => "01010000",5978 => "11111000",5979 => "00011010",5980 => "11100111",5981 => "01011110",5982 => "10010000",5983 => "11101000",5984 => "10111110",5985 => "10100111",5986 => "01111111",5987 => "01010000",5988 => "00010110",5989 => "10110001",5990 => "00111111",5991 => "01000111",5992 => "00110101",5993 => "00001001",5994 => "10011111",5995 => "00000000",5996 => "11000100",5997 => "10101000",5998 => "11001010",5999 => "01000000",6000 => "10111001",6001 => "00011000",6002 => "01110010",6003 => "01001010",6004 => "01111100",6005 => "01011101",6006 => "11111101",6007 => "00101010",6008 => "10100110",6009 => "00011010",6010 => "10111000",6011 => "00100010",6012 => "10000111",6013 => "10000000",6014 => "00111111",6015 => "11010001",6016 => "01000101",6017 => "01100011",6018 => "10011010",6019 => "11001101",6020 => "00101001",6021 => "10101010",6022 => "01011010",6023 => "01110101",6024 => "11001010",6025 => "11011010",6026 => "00101111",6027 => "11010101",6028 => "01010100",6029 => "11111100",6030 => "11010001",6031 => "01101110",6032 => "11010110",6033 => "01110111",6034 => "10011010",6035 => "01110101",6036 => "11101001",6037 => "00011111",6038 => "10010010",6039 => "00101011",6040 => "11100001",6041 => "01100000",6042 => "01001110",6043 => "10111100",6044 => "01101111",6045 => "01010100",6046 => "11000110",6047 => "00010110",6048 => "10100100",6049 => "00000010",6050 => "01110010",6051 => "11100011",6052 => "11110011",6053 => "10000011",6054 => "00110100",6055 => "10011010",6056 => "11100101",6057 => "10111000",6058 => "11100001",6059 => "11001110",6060 => "00000111",6061 => "10101011",6062 => "01001001",6063 => "01101101",6064 => "01011110",6065 => "01110011",6066 => "01010100",6067 => "00100100",6068 => "10110011",6069 => "01100100",6070 => "01011011",6071 => "10101000",6072 => "11001010",6073 => "11010110",6074 => "10011100",6075 => "01110111",6076 => "11011110",6077 => "11110100",6078 => "11111111",6079 => "10000110",6080 => "01101011",6081 => "10011000",6082 => "10101100",6083 => "00100010",6084 => "00100001",6085 => "11011010",6086 => "11101010",6087 => "00111010",6088 => "01101101",6089 => "01001010",6090 => "10011100",6091 => "00011010",6092 => "01010000",6093 => "01010100",6094 => "10010101",6095 => "10111000",6096 => "10011000",6097 => "11001010",6098 => "00000000",6099 => "10101000",6100 => "11101001",6101 => "10110001",6102 => "00010110",6103 => "11100001",6104 => "00001110",6105 => "00110010",6106 => "11101101",6107 => "10010100",6108 => "11110110",6109 => "00111110",6110 => "11101101",6111 => "10010111",6112 => "01111101",6113 => "10100100",6114 => "11011000",6115 => "00000111",6116 => "00011101",6117 => "00101011",6118 => "00111000",6119 => "11011101",6120 => "11100010",6121 => "01100101",6122 => "00011100",6123 => "10111100",6124 => "11010110",6125 => "01100111",6126 => "11010100",6127 => "11000110",6128 => "00110001",6129 => "11001001",6130 => "00100010",6131 => "10001110",6132 => "00000111",6133 => "11011111",6134 => "11001001",6135 => "10110111",6136 => "01100010",6137 => "01110000",6138 => "01000001",6139 => "11000100",6140 => "10100110",6141 => "00011000",6142 => "00000000",6143 => "11101111",6144 => "00100101",6145 => "11010100",6146 => "01010111",6147 => "11111111",6148 => "01011101",6149 => "01111011",6150 => "00101100",6151 => "10101111",6152 => "10000001",6153 => "10101101",6154 => "11110001",6155 => "10010101",6156 => "00100100",6157 => "01101111",6158 => "10010011",6159 => "11011000",6160 => "10101011",6161 => "01000101",6162 => "10010000",6163 => "10000111",6164 => "00000100",6165 => "10001000",6166 => "10010010",6167 => "11011101",6168 => "10110110",6169 => "00110011",6170 => "11100001",6171 => "10000000",6172 => "00101001",6173 => "00000111",6174 => "00100010",6175 => "01010100",6176 => "10001100",6177 => "01101000",6178 => "00110100",6179 => "01101011",6180 => "10010000",6181 => "01100100",6182 => "10110000",6183 => "10101001",6184 => "11100111",6185 => "11001001",6186 => "01000011",6187 => "10101001",6188 => "01100111",6189 => "00011011",6190 => "01010111",6191 => "10011100",6192 => "11011011",6193 => "01101001",6194 => "10110101",6195 => "01101110",6196 => "00001010",6197 => "10010100",6198 => "01111100",6199 => "01001001",6200 => "00010100",6201 => "00110111",6202 => "01101111",6203 => "10000010",6204 => "11111000",6205 => "01110100",6206 => "01101011",6207 => "11101001",6208 => "00010001",6209 => "10011010",6210 => "00001110",6211 => "00101100",6212 => "01101110",6213 => "11111000",6214 => "10111101",6215 => "01001101",6216 => "01000001",6217 => "11011011",6218 => "10111111",6219 => "01000011",6220 => "00011000",6221 => "00011000",6222 => "10111011",6223 => "11011011",6224 => "11001100",6225 => "10010010",6226 => "00011010",6227 => "11110001",6228 => "00110101",6229 => "10010010",6230 => "00110001",6231 => "00100111",6232 => "00011001",6233 => "00100000",6234 => "11101010",6235 => "11100001",6236 => "10001001",6237 => "00110010",6238 => "11010011",6239 => "01101011",6240 => "00101110",6241 => "10110011",6242 => "01000001",6243 => "11110111",6244 => "11101010",6245 => "01000100",6246 => "11001110",6247 => "10001000",6248 => "11000111",6249 => "00010110",6250 => "10011001",6251 => "00011000",6252 => "00000100",6253 => "11101001",6254 => "11111110",6255 => "10110010",6256 => "01011111",6257 => "00011100",6258 => "11010010",6259 => "00000101",6260 => "01110101",6261 => "00101100",6262 => "11111001",6263 => "10110100",6264 => "00001110",6265 => "11110010",6266 => "11010011",6267 => "01001001",6268 => "01101111",6269 => "11111101",6270 => "10100000",6271 => "01100111",6272 => "10000010",6273 => "11000011",6274 => "01100110",6275 => "01111111",6276 => "10100111",6277 => "00111111",6278 => "00000010",6279 => "01010110",6280 => "00100101",6281 => "10100101",6282 => "00110100",6283 => "10010010",6284 => "01110000",6285 => "10010110",6286 => "10010100",6287 => "00000100",6288 => "11100111",6289 => "01010011",6290 => "10101100",6291 => "01000111",6292 => "11111110",6293 => "10110101",6294 => "00000010",6295 => "11110110",6296 => "01111001",6297 => "00001100",6298 => "00001000",6299 => "10000010",6300 => "00111011",6301 => "11001001",6302 => "01100010",6303 => "11010010",6304 => "10111111",6305 => "10101000",6306 => "10111110",6307 => "00010011",6308 => "11110100",6309 => "01111010",6310 => "01001001",6311 => "10001111",6312 => "11000010",6313 => "00110111",6314 => "00011000",6315 => "00010011",6316 => "10100010",6317 => "00011001",6318 => "10010110",6319 => "00101001",6320 => "11100010",6321 => "00101010",6322 => "11110010",6323 => "11001110",6324 => "01000111",6325 => "00101101",6326 => "00000100",6327 => "10101001",6328 => "10010011",6329 => "11111101",6330 => "11011111",6331 => "00000100",6332 => "11001000",6333 => "11101110",6334 => "00111100",6335 => "11001110",6336 => "00011111",6337 => "01010001",6338 => "00101100",6339 => "11010100",6340 => "00110000",6341 => "00011001",6342 => "11110111",6343 => "00100110",6344 => "10010011",6345 => "00000101",6346 => "10110010",6347 => "00100001",6348 => "11000001",6349 => "00111001",6350 => "00100100",6351 => "11010011",6352 => "11010011",6353 => "00000010",6354 => "00110011",6355 => "00110000",6356 => "00111101",6357 => "00111101",6358 => "00011111",6359 => "10110001",6360 => "01000101",6361 => "11010111",6362 => "00111101",6363 => "11010101",6364 => "10101100",6365 => "11011011",6366 => "10100010",6367 => "01101110",6368 => "11101001",6369 => "10110011",6370 => "01011001",6371 => "01110100",6372 => "10111100",6373 => "01000110",6374 => "00101010",6375 => "11011101",6376 => "10000001",6377 => "10100000",6378 => "00001000",6379 => "01101110",6380 => "11001001",6381 => "11010111",6382 => "11001000",6383 => "00111011",6384 => "11000001",6385 => "01101001",6386 => "00000001",6387 => "01101010",6388 => "11000101",6389 => "01110001",6390 => "11110111",6391 => "00101011",6392 => "10011100",6393 => "10111100",6394 => "10011110",6395 => "11001001",6396 => "00001001",6397 => "11101111",6398 => "10100001",6399 => "00110111",6400 => "01000001",6401 => "11000001",6402 => "11100110",6403 => "01110110",6404 => "01000110",6405 => "00001100",6406 => "10011110",6407 => "11000101",6408 => "01000001",6409 => "01001001",6410 => "10001101",6411 => "10011000",6412 => "10001001",6413 => "01010001",6414 => "10000010",6415 => "10110101",6416 => "01000001",6417 => "00111010",6418 => "00000000",6419 => "00110010",6420 => "01010000",6421 => "01011111",6422 => "00101111",6423 => "10111000",6424 => "01100110",6425 => "10111001",6426 => "10001011",6427 => "01111110",6428 => "10110000",6429 => "10101000",6430 => "10100000",6431 => "10100000",6432 => "01111011",6433 => "01010011",6434 => "10011101",6435 => "01101001",6436 => "01011000",6437 => "00101111",6438 => "11011101",6439 => "00001000",6440 => "00010101",6441 => "00100011",6442 => "00101100",6443 => "11001111",6444 => "11011000",6445 => "00101010",6446 => "11000110",6447 => "00010110",6448 => "00011000",6449 => "10101100",6450 => "11101100",6451 => "00010111",6452 => "11101000",6453 => "00001110",6454 => "00100101",6455 => "00001100",6456 => "00100100",6457 => "01111011",6458 => "10001001",6459 => "10111111",6460 => "10100110",6461 => "11000101",6462 => "00100000",6463 => "11100010",6464 => "00000101",6465 => "00000111",6466 => "11011000",6467 => "10100000",6468 => "10001100",6469 => "01100011",6470 => "01000011",6471 => "11110011",6472 => "11001100",6473 => "01001010",6474 => "11011001",6475 => "11110000",6476 => "01001101",6477 => "11001101",6478 => "01100100",6479 => "11001110",6480 => "00000111",6481 => "11011001",6482 => "10111001",6483 => "01000010",6484 => "01101011",6485 => "01110001",6486 => "01001000",6487 => "01001001",6488 => "00001100",6489 => "00001011",6490 => "11000100",6491 => "11000110",6492 => "01111111",6493 => "11110110",6494 => "00011010",6495 => "11111011",6496 => "10010100",6497 => "11011100",6498 => "01111011",6499 => "10101101",6500 => "00111010",6501 => "01000010",6502 => "11001011",6503 => "00010000",6504 => "00111101",6505 => "10010001",6506 => "11100011",6507 => "10110001",6508 => "00001111",6509 => "11111111",6510 => "01111111",6511 => "01101001",6512 => "01110010",6513 => "11011110",6514 => "00111110",6515 => "00111011",6516 => "00001110",6517 => "00101111",6518 => "10001011",6519 => "01010000",6520 => "00000111",6521 => "00000110",6522 => "01011011",6523 => "01101110",6524 => "00011000",6525 => "10010000",6526 => "01011100",6527 => "00111001",6528 => "00011100",6529 => "00011000",6530 => "10100100",6531 => "00010101",6532 => "01111100",6533 => "10111001",6534 => "10101110",6535 => "11101000",6536 => "10111100",6537 => "10101000",6538 => "11000000",6539 => "01110000",6540 => "10111001",6541 => "01010001",6542 => "10010010",6543 => "11100100",6544 => "11101001",6545 => "10100100",6546 => "00100101",6547 => "11101110",6548 => "00101101",6549 => "00001111",6550 => "00111101",6551 => "11010010",6552 => "11110001",6553 => "10110000",6554 => "11000001",6555 => "01001111",6556 => "00011101",6557 => "01011011",6558 => "10101101",6559 => "10111000",6560 => "00010100",6561 => "10000011",6562 => "11110001",6563 => "01110001",6564 => "00000101",6565 => "11100101",6566 => "10010110",6567 => "01000110",6568 => "10011111",6569 => "01111100",6570 => "10001001",6571 => "11000110",6572 => "01001100",6573 => "10100000",6574 => "00010111",6575 => "10000100",6576 => "10101000",6577 => "10000000",6578 => "10001100",6579 => "00011110",6580 => "01100011",6581 => "01000111",6582 => "00111111",6583 => "11101000",6584 => "01101001",6585 => "11001010",6586 => "10100000",6587 => "01011000",6588 => "00101010",6589 => "01111111",6590 => "10010010",6591 => "10100001",6592 => "10011110",6593 => "01000010",6594 => "10111000",6595 => "00000111",6596 => "11111100",6597 => "00001010",6598 => "01010100",6599 => "11101110",6600 => "10101001",6601 => "11011010",6602 => "01101010",6603 => "10101111",6604 => "10100000",6605 => "00110010",6606 => "11000011",6607 => "00000101",6608 => "10010000",6609 => "00100110",6610 => "01110100",6611 => "11111010",6612 => "10111100",6613 => "01010100",6614 => "00101110",6615 => "00010111",6616 => "11000000",6617 => "10101101",6618 => "00000111",6619 => "10100000",6620 => "10010010",6621 => "00000010",6622 => "11110010",6623 => "01101100",6624 => "10000100",6625 => "11011001",6626 => "10000111",6627 => "00010101",6628 => "01011010",6629 => "00011000",6630 => "10100011",6631 => "10001101",6632 => "10100111",6633 => "00010000",6634 => "01010000",6635 => "11001101",6636 => "11001100",6637 => "10100111",6638 => "01101100",6639 => "11011100",6640 => "10100110",6641 => "00001011",6642 => "10000011",6643 => "00001001",6644 => "10001101",6645 => "01100111",6646 => "00001010",6647 => "01101101",6648 => "01011101",6649 => "01000011",6650 => "11010111",6651 => "10101111",6652 => "10110010",6653 => "11111110",6654 => "10111010",6655 => "01000110",6656 => "10001001",6657 => "11101100",6658 => "10001110",6659 => "10101000",6660 => "11111000",6661 => "10100110",6662 => "00000101",6663 => "00000111",6664 => "11101010",6665 => "10100011",6666 => "11101101",6667 => "10110100",6668 => "01000011",6669 => "10000110",6670 => "01110111",6671 => "01101010",6672 => "11011010",6673 => "00111011",6674 => "00111101",6675 => "00101101",6676 => "10101100",6677 => "01100011",6678 => "11001010",6679 => "10001110",6680 => "10110100",6681 => "10110101",6682 => "00010100",6683 => "01111111",6684 => "11000001",6685 => "11001111",6686 => "11001011",6687 => "00011011",6688 => "00101101",6689 => "00010101",6690 => "01101101",6691 => "10000011",6692 => "01100101",6693 => "01101101",6694 => "01010111",6695 => "10111011",6696 => "11110101",6697 => "11110111",6698 => "01100011",6699 => "10100110",6700 => "11100001",6701 => "11100100",6702 => "10110110",6703 => "10011000",6704 => "00110101",6705 => "01110000",6706 => "11011111",6707 => "11001111",6708 => "00100010",6709 => "00011101",6710 => "00110011",6711 => "01000100",6712 => "01110000",6713 => "01110011",6714 => "11110111",6715 => "00100110",6716 => "11011011",6717 => "10111111",6718 => "00001010",6719 => "10100111",6720 => "01111000",6721 => "10001000",6722 => "00010100",6723 => "11101100",6724 => "10010101",6725 => "01110011",6726 => "00010011",6727 => "10011100",6728 => "11010100",6729 => "10010001",6730 => "01110011",6731 => "01100010",6732 => "11100101",6733 => "10010010",6734 => "01000000",6735 => "00010110",6736 => "11100000",6737 => "01010011",6738 => "00101111",6739 => "00011101",6740 => "10000000",6741 => "11101111",6742 => "10010100",6743 => "11011101",6744 => "11110000",6745 => "11100111",6746 => "10111101",6747 => "11101110",6748 => "11011011",6749 => "01011001",6750 => "11100010",6751 => "00110001",6752 => "11001000",6753 => "01001001",6754 => "10111100",6755 => "10000011",6756 => "11010000",6757 => "01000011",6758 => "10111001",6759 => "11001000",6760 => "01000011",6761 => "10001110",6762 => "10100011",6763 => "00001011",6764 => "11110110",6765 => "01000001",6766 => "01100110",6767 => "01001110",6768 => "01101111",6769 => "01010110",6770 => "00100001",6771 => "11011110",6772 => "11100000",6773 => "00001000",6774 => "00000111",6775 => "01101101",6776 => "00111101",6777 => "11100010",6778 => "10101001",6779 => "00110111",6780 => "11010111",6781 => "00110010",6782 => "01001101",6783 => "00000111",6784 => "10111000",6785 => "11011010",6786 => "00011100",6787 => "01110000",6788 => "00011111",6789 => "00010001",6790 => "00000001",6791 => "00000111",6792 => "00101111",6793 => "01110101",6794 => "00000110",6795 => "01111010",6796 => "10000001",6797 => "00111001",6798 => "01101100",6799 => "00000011",6800 => "00101011",6801 => "00100110",6802 => "11001001",6803 => "00101111",6804 => "00101001",6805 => "01001110",6806 => "11001101",6807 => "00001110",6808 => "01010000",6809 => "11100100",6810 => "01110001",6811 => "10011111",6812 => "10010101",6813 => "00000111",6814 => "01001110",6815 => "11010010",6816 => "11000000",6817 => "11000011",6818 => "01011011",6819 => "11111001",6820 => "10001110",6821 => "11100000",6822 => "00111000",6823 => "10111001",6824 => "11001110",6825 => "00000011",6826 => "01011001",6827 => "11110011",6828 => "01001101",6829 => "00000001",6830 => "10110000",6831 => "00111000",6832 => "01011001",6833 => "01000001",6834 => "11111010",6835 => "10010110",6836 => "11011001",6837 => "10100010",6838 => "00001000",6839 => "01100111",6840 => "00101111",6841 => "10011011",6842 => "00100101",6843 => "11010100",6844 => "00110010",6845 => "00000011",6846 => "10110110",6847 => "00001101",6848 => "11011010",6849 => "00100010",6850 => "01110110",6851 => "11000010",6852 => "00100110",6853 => "01010001",6854 => "00011111",6855 => "10100101",6856 => "10001101",6857 => "11100000",6858 => "00011001",6859 => "00010001",6860 => "11101001",6861 => "10011011",6862 => "10001110",6863 => "10000111",6864 => "00101001",6865 => "11001011",6866 => "01110100",6867 => "10001010",6868 => "11101000",6869 => "10100001",6870 => "11110011",6871 => "00010000",6872 => "11010000",6873 => "10010001",6874 => "01101111",6875 => "10110110",6876 => "01110101",6877 => "11000101",6878 => "00000111",6879 => "10010001",6880 => "01001101",6881 => "11000110",6882 => "10111000",6883 => "11011110",6884 => "01101110",6885 => "10000100",6886 => "01111111",6887 => "01110010",6888 => "10011001",6889 => "01111000",6890 => "01110101",6891 => "00011110",6892 => "01111110",6893 => "01001011",6894 => "01101010",6895 => "11110110",6896 => "00010111",6897 => "01001000",6898 => "10001011",6899 => "11001101",6900 => "00100011",6901 => "11011010",6902 => "00011011",6903 => "11100101",6904 => "11101100",6905 => "01100001",6906 => "11000110",6907 => "01111000",6908 => "00001000",6909 => "01011100",6910 => "00101111",6911 => "10110111",6912 => "00100101",6913 => "01101001",6914 => "10110101",6915 => "11111100",6916 => "11100101",6917 => "00111100",6918 => "11101001",6919 => "00001101",6920 => "01100101",6921 => "00011111",6922 => "00100001",6923 => "11011101",6924 => "00100000",6925 => "01011111",6926 => "11011100",6927 => "11011101",6928 => "00111100",6929 => "00011100",6930 => "10011111",6931 => "11011100",6932 => "10000110",6933 => "01100111",6934 => "00001001",6935 => "11001110",6936 => "01111010",6937 => "11011010",6938 => "10001111",6939 => "10011111",6940 => "11111111",6941 => "01101011",6942 => "01101000",6943 => "10111110",6944 => "01000001",6945 => "00101100",6946 => "10111110",6947 => "00010011",6948 => "10110000",6949 => "10101011",6950 => "10100111",6951 => "11111101",6952 => "10010111",6953 => "01101101",6954 => "10011110",6955 => "11101110",6956 => "11100100",6957 => "11111100",6958 => "01010001",6959 => "11000011",6960 => "01101111",6961 => "01101011",6962 => "10010111",6963 => "00101010",6964 => "11110111",6965 => "00001010",6966 => "10100010",6967 => "10100011",6968 => "11111001",6969 => "10011011",6970 => "01000010",6971 => "10011001",6972 => "01101001",6973 => "11010110",6974 => "10100110",6975 => "00101100",6976 => "01001110",6977 => "01110101",6978 => "11101000",6979 => "01101100",6980 => "00011110",6981 => "00010111",6982 => "10011000",6983 => "10100101",6984 => "11000100",6985 => "01011011",6986 => "10010010",6987 => "00101001",6988 => "10000010",6989 => "11100011",6990 => "01001001",6991 => "10001100",6992 => "11111111",6993 => "01011110",6994 => "11101000",6995 => "11001000",6996 => "10010001",6997 => "11000000",6998 => "10101111",6999 => "01100011",7000 => "01111111",7001 => "00011111",7002 => "10011010",7003 => "01111101",7004 => "10101001",7005 => "10100000",7006 => "00111100",7007 => "01011011",7008 => "11110101",7009 => "00001000",7010 => "01100011",7011 => "11110010",7012 => "01010110",7013 => "11001101",7014 => "11101101",7015 => "11000101",7016 => "00100001",7017 => "11111100",7018 => "01110011",7019 => "10001010",7020 => "01111100",7021 => "10101000",7022 => "01100000",7023 => "10001110",7024 => "11110111",7025 => "00011010",7026 => "10011111",7027 => "00110010",7028 => "10111011",7029 => "10001000",7030 => "00101111",7031 => "00010010",7032 => "00000010",7033 => "00011001",7034 => "00110110",7035 => "10111101",7036 => "11000110",7037 => "11010111",7038 => "00001000",7039 => "01101000",7040 => "11000111",7041 => "00011010",7042 => "01111000",7043 => "10101011",7044 => "11011100",7045 => "00011011",7046 => "10000011",7047 => "10001111",7048 => "10010000",7049 => "00001011",7050 => "00111001",7051 => "10011010",7052 => "10010110",7053 => "11100101",7054 => "00110111",7055 => "11000001",7056 => "11101111",7057 => "10101011",7058 => "11000011",7059 => "10000111",7060 => "11110110",7061 => "01010101",7062 => "00100011",7063 => "11110010",7064 => "11110010",7065 => "00010000",7066 => "10101110",7067 => "00000111",7068 => "01001100",7069 => "00101101",7070 => "00001011",7071 => "00010011",7072 => "00111010",7073 => "10101101",7074 => "11011101",7075 => "00101011",7076 => "01110111",7077 => "10000001",7078 => "01010000",7079 => "00001100",7080 => "10110101",7081 => "00011000",7082 => "01001011",7083 => "01110100",7084 => "00111001",7085 => "00111001",7086 => "01100101",7087 => "01011010",7088 => "11111000",7089 => "11111101",7090 => "11010111",7091 => "11001000",7092 => "00101010",7093 => "01001000",7094 => "10000001",7095 => "01011111",7096 => "00001010",7097 => "10110111",7098 => "10010101",7099 => "10100011",7100 => "11111101",7101 => "11101110",7102 => "10010111",7103 => "10100000",7104 => "01100010",7105 => "10101001",7106 => "10101110",7107 => "00011001",7108 => "10011011",7109 => "11100110",7110 => "00100101",7111 => "10000001",7112 => "01000110",7113 => "01110001",7114 => "00100000",7115 => "00001100",7116 => "11011100",7117 => "10111100",7118 => "00011001",7119 => "01101100",7120 => "01010011",7121 => "00111100",7122 => "11001100",7123 => "10010110",7124 => "10100100",7125 => "00111110",7126 => "01001101",7127 => "00010111",7128 => "01110110",7129 => "00101010",7130 => "11000000",7131 => "01100001",7132 => "11100101",7133 => "01001000",7134 => "00000001",7135 => "01011011",7136 => "01101110",7137 => "00000101",7138 => "10010100",7139 => "00011010",7140 => "01110010",7141 => "01010111",7142 => "11101100",7143 => "00100111",7144 => "10000100",7145 => "00000101",7146 => "11111111",7147 => "10000111",7148 => "01010000",7149 => "00000010",7150 => "00101010",7151 => "11110101",7152 => "01010100",7153 => "00101000",7154 => "00100001",7155 => "11001000",7156 => "00010100",7157 => "11101110",7158 => "11010000",7159 => "10010110",7160 => "10001111",7161 => "01111101",7162 => "00100110",7163 => "01001110",7164 => "11110000",7165 => "01111001",7166 => "01010000",7167 => "00011000",7168 => "01010001",7169 => "00000101",7170 => "01100100",7171 => "01110010",7172 => "00100011",7173 => "11101110",7174 => "01110011",7175 => "00110101",7176 => "01000000",7177 => "01111101",7178 => "01110111",7179 => "11000000",7180 => "00010101",7181 => "00111111",7182 => "01011111",7183 => "10001011",7184 => "00100010",7185 => "11110010",7186 => "01100011",7187 => "00110101",7188 => "01010010",7189 => "00001011",7190 => "10000000",7191 => "00100000",7192 => "10110001",7193 => "10011001",7194 => "11010000",7195 => "01101100",7196 => "01111001",7197 => "10100011",7198 => "11001111",7199 => "11100101",7200 => "11010001",7201 => "01010110",7202 => "10000110",7203 => "01001110",7204 => "10110100",7205 => "10000111",7206 => "00000010",7207 => "01101011",7208 => "11001000",7209 => "11110100",7210 => "11100110",7211 => "11011001",7212 => "01110000",7213 => "00001011",7214 => "10110111",7215 => "01101011",7216 => "11101110",7217 => "01111111",7218 => "01001101",7219 => "10001000",7220 => "01010000",7221 => "01011001",7222 => "01101000",7223 => "10110100",7224 => "10010010",7225 => "00010100",7226 => "01011000",7227 => "00000111",7228 => "00111111",7229 => "10001000",7230 => "00001100",7231 => "00100001",7232 => "10101001",7233 => "01111001",7234 => "01011110",7235 => "01100101",7236 => "00111111",7237 => "01110101",7238 => "00000001",7239 => "00000000",7240 => "11101100",7241 => "00101110",7242 => "01110100",7243 => "10001110",7244 => "11000011",7245 => "10000000",7246 => "10001100",7247 => "10001101",7248 => "00100010",7249 => "00001100",7250 => "10011010",7251 => "11110110",7252 => "01100011",7253 => "10101100",7254 => "00000110",7255 => "01100111",7256 => "11010101",7257 => "10000100",7258 => "10100001",7259 => "01111101",7260 => "10000110",7261 => "10101010",7262 => "11111000",7263 => "10111111",7264 => "11101010",7265 => "01110100",7266 => "11101100",7267 => "11101011",7268 => "00101011",7269 => "01000101",7270 => "00001001",7271 => "11001100",7272 => "11110000",7273 => "00001100",7274 => "01101111",7275 => "10011001",7276 => "11111110",7277 => "00010010",7278 => "11100101",7279 => "01100101",7280 => "10000010",7281 => "11111111",7282 => "10111010",7283 => "10001100",7284 => "10010011",7285 => "11110001",7286 => "00000011",7287 => "10101101",7288 => "11101101",7289 => "00000101",7290 => "10010001",7291 => "11001100",7292 => "11001101",7293 => "10101000",7294 => "10100111",7295 => "11000111",7296 => "11011010",7297 => "11000111",7298 => "10000001",7299 => "00001101",7300 => "01001010",7301 => "10111111",7302 => "01010001",7303 => "01010111",7304 => "11000010",7305 => "00010110",7306 => "00111101",7307 => "01110010",7308 => "10011100",7309 => "01000010",7310 => "00011111",7311 => "01111101",7312 => "00011011",7313 => "01000010",7314 => "10101101",7315 => "01010001",7316 => "01010010",7317 => "01011010",7318 => "01010100",7319 => "00001011",7320 => "11010010",7321 => "11111011",7322 => "11000011",7323 => "10001101",7324 => "10111001",7325 => "01110010",7326 => "10111011",7327 => "01001001",7328 => "10100110",7329 => "01111010",7330 => "01011101",7331 => "10000111",7332 => "01100101",7333 => "01000001",7334 => "10000111",7335 => "11111010",7336 => "11110100",7337 => "11101000",7338 => "10010010",7339 => "00101100",7340 => "11100010",7341 => "01111101",7342 => "01100001",7343 => "10101010",7344 => "11101010",7345 => "10110010",7346 => "11000001",7347 => "01011011",7348 => "10110011",7349 => "10111111",7350 => "11101110",7351 => "01000010",7352 => "00111100",7353 => "10011101",7354 => "10010101",7355 => "11110101",7356 => "11010000",7357 => "00100110",7358 => "00101010",7359 => "00011101",7360 => "11011110",7361 => "01111100",7362 => "01001101",7363 => "10010000",7364 => "00100010",7365 => "01101100",7366 => "01000011",7367 => "00101000",7368 => "10100101",7369 => "11111100",7370 => "01110011",7371 => "00110000",7372 => "10111101",7373 => "00011100",7374 => "01011100",7375 => "01010110",7376 => "01110010",7377 => "10001111",7378 => "11010011",7379 => "10111110",7380 => "00011101",7381 => "11011100",7382 => "11101001",7383 => "11101010",7384 => "10011001",7385 => "11011100",7386 => "00000001",7387 => "00011110",7388 => "01011000",7389 => "10101010",7390 => "11100100",7391 => "01110100",7392 => "10101011",7393 => "11010111",7394 => "10001000",7395 => "11011010",7396 => "00000011",7397 => "11001111",7398 => "11000111",7399 => "00111000",7400 => "01010001",7401 => "01100010",7402 => "10100100",7403 => "10000001",7404 => "11111100",7405 => "10111010",7406 => "10010110",7407 => "10010010",7408 => "00011110",7409 => "11011100",7410 => "01100011",7411 => "10000101",7412 => "01011010",7413 => "01000010",7414 => "01010010",7415 => "11100101",7416 => "10110010",7417 => "10011011",7418 => "01101101",7419 => "00100000",7420 => "10001100",7421 => "01111011",7422 => "11110010",7423 => "11000000",7424 => "11011110",7425 => "01011101",7426 => "11011110",7427 => "11010111",7428 => "11011000",7429 => "00111110",7430 => "10101001",7431 => "11100110",7432 => "00010001",7433 => "01101111",7434 => "11001000",7435 => "01011111",7436 => "11011101",7437 => "11011100",7438 => "10010101",7439 => "11011110",7440 => "00110111",7441 => "11100000",7442 => "10101000",7443 => "00101000",7444 => "01000000",7445 => "11101011",7446 => "10111101",7447 => "10110000",7448 => "01110011",7449 => "01010001",7450 => "01001101",7451 => "11010101",7452 => "10001001",7453 => "00001001",7454 => "11110011",7455 => "11110011",7456 => "01000110",7457 => "10111011",7458 => "11110000",7459 => "01101000",7460 => "11111101",7461 => "00111000",7462 => "00001001",7463 => "10000101",7464 => "00010111",7465 => "11010111",7466 => "00110011",7467 => "11010100",7468 => "10010111",7469 => "00000100",7470 => "01010001",7471 => "10000100",7472 => "00111000",7473 => "01000101",7474 => "00000100",7475 => "00001111",7476 => "11010100",7477 => "01110100",7478 => "10110111",7479 => "10110011",7480 => "00101000",7481 => "10110111",7482 => "00000001",7483 => "00100001",7484 => "01011111",7485 => "00110110",7486 => "11101101",7487 => "10011000",7488 => "11111110",7489 => "10100011",7490 => "11010000",7491 => "10100110",7492 => "00001111",7493 => "11001011",7494 => "10010011",7495 => "10111101",7496 => "11011110",7497 => "01000010",7498 => "01110100",7499 => "01110111",7500 => "11110100",7501 => "10001001",7502 => "01111010",7503 => "10110000",7504 => "11001000",7505 => "00010000",7506 => "11111011",7507 => "01101101",7508 => "11110000",7509 => "10110101",7510 => "00101011",7511 => "00001000",7512 => "00001100",7513 => "00000101",7514 => "11100100",7515 => "11010000",7516 => "00010101",7517 => "11101111",7518 => "10011111",7519 => "01011011",7520 => "11101010",7521 => "01101010",7522 => "11000010",7523 => "01000110",7524 => "00001011",7525 => "01111101",7526 => "11010001",7527 => "00000110",7528 => "01110101",7529 => "10000010",7530 => "10110010",7531 => "11110000",7532 => "01100110",7533 => "11101001",7534 => "10110010",7535 => "01111111",7536 => "01110010",7537 => "01000111",7538 => "00010110",7539 => "00111111",7540 => "00001111",7541 => "00110010",7542 => "00110010",7543 => "10000010",7544 => "00000011",7545 => "00111011",7546 => "01101111",7547 => "00001100",7548 => "01100001",7549 => "01010001",7550 => "01011010",7551 => "11101101",7552 => "11000101",7553 => "10000100",7554 => "11111100",7555 => "11101100",7556 => "11001000",7557 => "01001101",7558 => "00011100",7559 => "01100010",7560 => "00010001",7561 => "01010111",7562 => "00000101",7563 => "00011000",7564 => "10001100",7565 => "01100010",7566 => "10001111",7567 => "01110101",7568 => "10011100",7569 => "01100111",7570 => "01100000",7571 => "01110101",7572 => "11010011",7573 => "00101001",7574 => "01101111",7575 => "10010011",7576 => "10110111",7577 => "01100001",7578 => "00100100",7579 => "11110011",7580 => "01111101",7581 => "10100110",7582 => "11000001",7583 => "00101000",7584 => "00101010",7585 => "01111100",7586 => "11010000",7587 => "10010110",7588 => "00000001",7589 => "11110000",7590 => "10100100",7591 => "00000101",7592 => "10001011",7593 => "10111111",7594 => "01111110",7595 => "11100101",7596 => "01101101",7597 => "10101011",7598 => "01101110",7599 => "00011110",7600 => "10111110",7601 => "01101110",7602 => "11101000",7603 => "10011110",7604 => "00100001",7605 => "10101010",7606 => "11110100",7607 => "10111000",7608 => "11001111",7609 => "10010100",7610 => "00000111",7611 => "10001101",7612 => "01111101",7613 => "01010010",7614 => "00110101",7615 => "01100011",7616 => "01111101",7617 => "00110101",7618 => "10010110",7619 => "00000000",7620 => "10111001",7621 => "11101001",7622 => "01110010",7623 => "10011011",7624 => "00100111",7625 => "00110011",7626 => "10100110",7627 => "11011010",7628 => "00110011",7629 => "00011000",7630 => "00001000",7631 => "11000011",7632 => "01001011",7633 => "10011010",7634 => "00010001",7635 => "00001110",7636 => "00111001",7637 => "01111111",7638 => "11111011",7639 => "00010101",7640 => "11000001",7641 => "11011000",7642 => "00010110",7643 => "10010010",7644 => "01100010",7645 => "10111010",7646 => "01001010",7647 => "10010011",7648 => "11010001",7649 => "01011110",7650 => "00110101",7651 => "11110000",7652 => "01110000",7653 => "11000000",7654 => "10010101",7655 => "11011000",7656 => "00101011",7657 => "01010101",7658 => "10110010",7659 => "10010011",7660 => "01111000",7661 => "11110011",7662 => "00111011",7663 => "11100000",7664 => "00100101",7665 => "10111011",7666 => "00110111",7667 => "10111000",7668 => "11100110",7669 => "10001110",7670 => "00101010",7671 => "01100111",7672 => "11001001",7673 => "10111010",7674 => "01110000",7675 => "10101100",7676 => "10111100",7677 => "10101100",7678 => "10011101",7679 => "10111111",7680 => "00110000",7681 => "00011100",7682 => "01000110",7683 => "01000010",7684 => "00101000",7685 => "01111010",7686 => "01011100",7687 => "01011001",7688 => "10101111",7689 => "00011101",7690 => "00100010",7691 => "01011011",7692 => "11010010",7693 => "01110100",7694 => "10011011",7695 => "01001101",7696 => "00000110",7697 => "01010000",7698 => "10011101",7699 => "01011010",7700 => "01000010",7701 => "11000101",7702 => "10111000",7703 => "01000111",7704 => "11011100",7705 => "00010111",7706 => "01000100",7707 => "11110110",7708 => "00110111",7709 => "10100010",7710 => "10001000",7711 => "00010110",7712 => "00110000",7713 => "01001101",7714 => "11100011",7715 => "11101100",7716 => "10011111",7717 => "10010110",7718 => "11010100",7719 => "10011001",7720 => "01110010",7721 => "00010110",7722 => "11001110",7723 => "00001001",7724 => "10010011",7725 => "10001001",7726 => "11011101",7727 => "11110000",7728 => "01011010",7729 => "01000000",7730 => "00111010",7731 => "01010010",7732 => "00100010",7733 => "00100110",7734 => "11111000",7735 => "10101101",7736 => "00000011",7737 => "00111111",7738 => "10100100",7739 => "00111001",7740 => "00000010",7741 => "01000011",7742 => "10010100",7743 => "00011011",7744 => "00000100",7745 => "00000001",7746 => "01100101",7747 => "11001100",7748 => "11110001",7749 => "10010011",7750 => "01110101",7751 => "10000101",7752 => "10100100",7753 => "10000000",7754 => "10010010",7755 => "00000011",7756 => "01100011",7757 => "10110100",7758 => "11011001",7759 => "10100011",7760 => "01101100",7761 => "10100010",7762 => "01000111",7763 => "10110001",7764 => "10011111",7765 => "00110011",7766 => "11100100",7767 => "01101000",7768 => "10111100",7769 => "01110100",7770 => "00001010",7771 => "00010010",7772 => "01111100",7773 => "10101010",7774 => "10000010",7775 => "01010111",7776 => "00000011",7777 => "11100001",7778 => "01001001",7779 => "11010010",7780 => "00100101",7781 => "00010000",7782 => "01010110",7783 => "00001111",7784 => "00010011",7785 => "01100101",7786 => "01100101",7787 => "00010001",7788 => "00011100",7789 => "11000111",7790 => "01111000",7791 => "11010000",7792 => "01001001",7793 => "10000110",7794 => "11011011",7795 => "11001100",7796 => "10001100",7797 => "11001101",7798 => "10110101",7799 => "11010101",7800 => "00100110",7801 => "11100000",7802 => "00001000",7803 => "11110001",7804 => "00101001",7805 => "10110001",7806 => "10100100",7807 => "00110011",7808 => "11000101",7809 => "00101011",7810 => "10001000",7811 => "01100110",7812 => "00001111",7813 => "10110100",7814 => "11110010",7815 => "11000001",7816 => "11110100",7817 => "01010100",7818 => "10001111",7819 => "01101010",7820 => "10001100",7821 => "00111010",7822 => "01001110",7823 => "00011100",7824 => "10101101",7825 => "01010001",7826 => "01001001",7827 => "01000110",7828 => "01111110",7829 => "10111101",7830 => "11000001",7831 => "11010001",7832 => "10001010",7833 => "01110101",7834 => "11011010",7835 => "00100010",7836 => "00100000",7837 => "01000110",7838 => "01010111",7839 => "01100101",7840 => "01011001",7841 => "10000110",7842 => "01111010",7843 => "11010011",7844 => "00011010",7845 => "00011000",7846 => "11000110",7847 => "10000010",7848 => "10101000",7849 => "00010110",7850 => "00001111",7851 => "00110100",7852 => "11010111",7853 => "10110110",7854 => "01100001",7855 => "11100011",7856 => "01101010",7857 => "00000100",7858 => "00110101",7859 => "01101110",7860 => "11100001",7861 => "10010100",7862 => "10111000",7863 => "10101100",7864 => "00101100",7865 => "11010111",7866 => "10100010",7867 => "11110010",7868 => "00000011",7869 => "10100000",7870 => "00001001",7871 => "10010011",7872 => "00111111",7873 => "10010110",7874 => "10100110",7875 => "01000010",7876 => "11101110",7877 => "10100111",7878 => "10010011",7879 => "00100011",7880 => "00110111",7881 => "00010111",7882 => "11000100",7883 => "00110110",7884 => "11011101",7885 => "00100101",7886 => "11001010",7887 => "10110111",7888 => "10001101",7889 => "00010100",7890 => "01010011",7891 => "00001100",7892 => "00011111",7893 => "11010011",7894 => "11100000",7895 => "10000000",7896 => "00101110",7897 => "00100111",7898 => "00000100",7899 => "01010011",7900 => "00111001",7901 => "01111001",7902 => "00111001",7903 => "10100100",7904 => "10100100",7905 => "11000100",7906 => "11101000",7907 => "11010100",7908 => "01001011",7909 => "10111100",7910 => "01000011",7911 => "00100000",7912 => "00000110",7913 => "11101101",7914 => "11101001",7915 => "01101001",7916 => "11001011",7917 => "11010011",7918 => "01001111",7919 => "10010001",7920 => "11010100",7921 => "01011101",7922 => "11011000",7923 => "01111011",7924 => "10111011",7925 => "11000111",7926 => "01100010",7927 => "11101000",7928 => "11101011",7929 => "10001000",7930 => "10000110",7931 => "11101110",7932 => "10000001",7933 => "00111011",7934 => "11000011",7935 => "11100010",7936 => "11010010",7937 => "00101001",7938 => "11100001",7939 => "11001001",7940 => "11000010",7941 => "10100101",7942 => "11100000",7943 => "10101010",7944 => "01101000",7945 => "11100011",7946 => "01001000",7947 => "11000101",7948 => "11111101",7949 => "10111010",7950 => "10011100",7951 => "10010011",7952 => "10011110",7953 => "11111001",7954 => "11001011",7955 => "10011000",7956 => "00100011",7957 => "00110000",7958 => "00101111",7959 => "01010011",7960 => "10011101",7961 => "10011111",7962 => "11000111",7963 => "11011111",7964 => "10011100",7965 => "01100101",7966 => "00100001",7967 => "10101100",7968 => "10100011",7969 => "11001010",7970 => "00100101",7971 => "10000110",7972 => "11101101",7973 => "11001000",7974 => "01111110",7975 => "01010010",7976 => "01010100",7977 => "01111100",7978 => "00110101",7979 => "11101000",7980 => "10010001",7981 => "11000000",7982 => "10000100",7983 => "01010011",7984 => "01101110",7985 => "11111010",7986 => "01010000",7987 => "10110001",7988 => "11000011",7989 => "00111011",7990 => "10101011",7991 => "01000111",7992 => "00111010",7993 => "00011000",7994 => "10011001",7995 => "00111100",7996 => "01100001",7997 => "01001000",7998 => "00001101",7999 => "00110100",8000 => "01001101",8001 => "00011011",8002 => "11110001",8003 => "00101001",8004 => "10001110",8005 => "01111100",8006 => "00010001",8007 => "01111011",8008 => "10000110",8009 => "11001010",8010 => "00011101",8011 => "00111101",8012 => "10110001",8013 => "00001000",8014 => "00110010",8015 => "00100110",8016 => "01100001",8017 => "00000100",8018 => "01001101",8019 => "11100001",8020 => "10100011",8021 => "01111011",8022 => "01111110",8023 => "10100100",8024 => "10001101",8025 => "10100101",8026 => "00111110",8027 => "11011001",8028 => "10011100",8029 => "00110100",8030 => "10111110",8031 => "10111000",8032 => "01010000",8033 => "00011101",8034 => "11011010",8035 => "01100101",8036 => "01100000",8037 => "11000000",8038 => "11111100",8039 => "01111010",8040 => "10101000",8041 => "01110110",8042 => "11001000",8043 => "10100110",8044 => "11100010",8045 => "00111110",8046 => "00110010",8047 => "01101000",8048 => "01000101",8049 => "01010111",8050 => "10010111",8051 => "11001101",8052 => "10010011",8053 => "11100010",8054 => "10011001",8055 => "10011111",8056 => "10001110",8057 => "10110000",8058 => "11110100",8059 => "01101110",8060 => "00100000",8061 => "00010110",8062 => "01000011",8063 => "01101011",8064 => "10111111",8065 => "11100000",8066 => "11110100",8067 => "01101101",8068 => "01111011",8069 => "00101100",8070 => "11100010",8071 => "11010000",8072 => "11000011",8073 => "01111000",8074 => "01000001",8075 => "10101001",8076 => "10010010",8077 => "11110001",8078 => "10010111",8079 => "01110110",8080 => "10110101",8081 => "01000110",8082 => "01111001",8083 => "01110000",8084 => "11001100",8085 => "00110000",8086 => "10010110",8087 => "01001110",8088 => "01001000",8089 => "01010001",8090 => "00100011",8091 => "10010001",8092 => "01110011",8093 => "11000110",8094 => "10100010",8095 => "11101001",8096 => "11011101",8097 => "00111101",8098 => "11110010",8099 => "00000100",8100 => "00000101",8101 => "11101011",8102 => "11001010",8103 => "00111110",8104 => "01101000",8105 => "01111110",8106 => "01011111",8107 => "00111111",8108 => "01110100",8109 => "00010110",8110 => "00010011",8111 => "10001000",8112 => "11100010",8113 => "10111100",8114 => "10111011",8115 => "01011001",8116 => "00111010",8117 => "11011011",8118 => "11000100",8119 => "10001000",8120 => "10011010",8121 => "10010110",8122 => "01111001",8123 => "10000101",8124 => "01101111",8125 => "00011000",8126 => "11011100",8127 => "10001111",8128 => "11110110",8129 => "10111000",8130 => "00101010",8131 => "01111100",8132 => "01001011",8133 => "00110110",8134 => "11111011",8135 => "00001010",8136 => "11110001",8137 => "00111010",8138 => "00101111",8139 => "01011100",8140 => "10001110",8141 => "00101110",8142 => "10100010",8143 => "00111111",8144 => "11001001",8145 => "10100010",8146 => "11000110",8147 => "11101011",8148 => "00110110",8149 => "01000000",8150 => "11001110",8151 => "10011101",8152 => "11101011",8153 => "00101110",8154 => "00000111",8155 => "00100100",8156 => "01101000",8157 => "11110001",8158 => "01000110",8159 => "01110101",8160 => "01101111",8161 => "10111000",8162 => "01001001",8163 => "10110110",8164 => "10000100",8165 => "11100100",8166 => "11111010",8167 => "11101110",8168 => "10000111",8169 => "00110011",8170 => "01111111",8171 => "01111000",8172 => "00010011",8173 => "00010010",8174 => "01100000",8175 => "01110110",8176 => "00001100",8177 => "00001010",8178 => "00011101",8179 => "00110101",8180 => "00100000",8181 => "01001101",8182 => "11001001",8183 => "01010001",8184 => "10100111",8185 => "11010001",8186 => "00010001",8187 => "11110011",8188 => "11001010",8189 => "00110011",8190 => "11010000",8191 => "10001111",8192 => "10010111",8193 => "11101110",8194 => "11100101",8195 => "00101101",8196 => "11011111",8197 => "00001100",8198 => "01100011",8199 => "01000110",8200 => "00111100",8201 => "01101100",8202 => "00001001",8203 => "00001110",8204 => "00010010",8205 => "10111000",8206 => "11110011",8207 => "00000101",8208 => "01101001",8209 => "11110101",8210 => "00111011",8211 => "10101011",8212 => "01001100",8213 => "11110001",8214 => "10111011",8215 => "10010101",8216 => "00100100",8217 => "10001111",8218 => "01111110",8219 => "11001101",8220 => "11001011",8221 => "11111000",8222 => "01001110",8223 => "00111110",8224 => "11110010",8225 => "00001110",8226 => "11111001",8227 => "10110010",8228 => "01011010",8229 => "00110100",8230 => "01001011",8231 => "10000110",8232 => "10011011",8233 => "10010001",8234 => "10001111",8235 => "00011011",8236 => "11101011",8237 => "01000100",8238 => "01111110",8239 => "11100010",8240 => "11010100",8241 => "10011111",8242 => "10110101",8243 => "11101100",8244 => "11010011",8245 => "01101010",8246 => "01010101",8247 => "00000111",8248 => "01011011",8249 => "00000100",8250 => "10011001",8251 => "11100100",8252 => "11001011",8253 => "00000100",8254 => "11101011",8255 => "01010101",8256 => "01101100",8257 => "00110100",8258 => "11101101",8259 => "10111011",8260 => "10001000",8261 => "00101110",8262 => "00101000",8263 => "11101000",8264 => "01110101",8265 => "01110101",8266 => "10000000",8267 => "11001111",8268 => "11110001",8269 => "01100111",8270 => "00111001",8271 => "10101101",8272 => "00111011",8273 => "00001111",8274 => "11111110",8275 => "10110110",8276 => "11100001",8277 => "11101000",8278 => "10000011",8279 => "01000101",8280 => "01000010",8281 => "01101111",8282 => "00001001",8283 => "00001011",8284 => "11000111",8285 => "01010110",8286 => "01111001",8287 => "10001110",8288 => "10010101",8289 => "11111100",8290 => "01000111",8291 => "01001110",8292 => "00110011",8293 => "11000000",8294 => "11011101",8295 => "11110001",8296 => "11001100",8297 => "01011010",8298 => "10000001",8299 => "10101001",8300 => "11001100",8301 => "01001110",8302 => "10110100",8303 => "01000101",8304 => "00110111",8305 => "00100000",8306 => "00100000",8307 => "00010010",8308 => "10100111",8309 => "00111011",8310 => "01100001",8311 => "10010000",8312 => "11101001",8313 => "01111111",8314 => "10101000",8315 => "11110011",8316 => "11110101",8317 => "00001110",8318 => "11000100",8319 => "01011100",8320 => "11000000",8321 => "11001111",8322 => "00000110",8323 => "10111111",8324 => "01001001",8325 => "10101000",8326 => "00110001",8327 => "11101001",8328 => "00111001",8329 => "01101100",8330 => "10100101",8331 => "00111100",8332 => "11100110",8333 => "01000101",8334 => "11000001",8335 => "01010101",8336 => "10011100",8337 => "01010010",8338 => "01001011",8339 => "00000111",8340 => "00110110",8341 => "00001001",8342 => "10101001",8343 => "10010001",8344 => "11011100",8345 => "00100010",8346 => "00110010",8347 => "10111011",8348 => "10101101",8349 => "00000000",8350 => "01001100",8351 => "00111100",8352 => "00001111",8353 => "01100101",8354 => "11000001",8355 => "10000000",8356 => "11111010",8357 => "00110001",8358 => "11000101",8359 => "10001110",8360 => "10110010",8361 => "11010000",8362 => "01010011",8363 => "01110100",8364 => "11100001",8365 => "00011000",8366 => "10001110",8367 => "10101001",8368 => "11000101",8369 => "00110011",8370 => "10101111",8371 => "01101010",8372 => "01110111",8373 => "00000100",8374 => "01110101",8375 => "00011000",8376 => "01111101",8377 => "11101101",8378 => "11101001",8379 => "11110011",8380 => "00001001",8381 => "10101010",8382 => "11000000",8383 => "00011011",8384 => "00100100",8385 => "00011000",8386 => "00010000",8387 => "01110010",8388 => "11110000",8389 => "00101010",8390 => "01110011",8391 => "11011000",8392 => "01111101",8393 => "10100111",8394 => "10110111",8395 => "11000000",8396 => "01110010",8397 => "11110001",8398 => "10011110",8399 => "00101110",8400 => "00011101",8401 => "01100101",8402 => "00010000",8403 => "10100111",8404 => "01011001",8405 => "11000001",8406 => "00111001",8407 => "00101111",8408 => "01100110",8409 => "00000000",8410 => "11111100",8411 => "01011011",8412 => "10111000",8413 => "00111111",8414 => "00011011",8415 => "10000110",8416 => "10101011",8417 => "01010110",8418 => "00111011",8419 => "01101010",8420 => "10011011",8421 => "00011000",8422 => "11011011",8423 => "11111011",8424 => "00010011",8425 => "11101100",8426 => "11001001",8427 => "11101011",8428 => "01000111",8429 => "00100001",8430 => "10100010",8431 => "10010110",8432 => "01100110",8433 => "10011110",8434 => "10011000",8435 => "10110101",8436 => "10010001",8437 => "01000110",8438 => "10110010",8439 => "10000001",8440 => "11110100",8441 => "01101110",8442 => "00010111",8443 => "11010000",8444 => "00100011",8445 => "01100001",8446 => "10100100",8447 => "11100100",8448 => "10110011",8449 => "10101100",8450 => "01011000",8451 => "10000110",8452 => "11110101",8453 => "11011100",8454 => "10000111",8455 => "01010100",8456 => "00010101",8457 => "11010001",8458 => "01001011",8459 => "00000111",8460 => "01011111",8461 => "11100010",8462 => "00001010",8463 => "11101101",8464 => "00001101",8465 => "00101100",8466 => "10000011",8467 => "10110101",8468 => "00111000",8469 => "10111010",8470 => "01001100",8471 => "01001011",8472 => "01010101",8473 => "11101010",8474 => "00101110",8475 => "00111000",8476 => "10000001",8477 => "01000100",8478 => "01001010",8479 => "10101110",8480 => "01011110",8481 => "01111010",8482 => "00101100",8483 => "10000001",8484 => "11101100",8485 => "11011100",8486 => "10111111",8487 => "01101111",8488 => "01110000",8489 => "10110011",8490 => "01100111",8491 => "01100111",8492 => "01010010",8493 => "01100101",8494 => "00010111",8495 => "00101111",8496 => "11001010",8497 => "10001110",8498 => "10110100",8499 => "00110100",8500 => "11010000",8501 => "11100010",8502 => "00001011",8503 => "00010110",8504 => "01011111",8505 => "00111000",8506 => "10001000",8507 => "10110001",8508 => "10011100",8509 => "01001110",8510 => "01100100",8511 => "11001000",8512 => "11111011",8513 => "01101000",8514 => "11110001",8515 => "01100001",8516 => "11101111",8517 => "00100110",8518 => "11000100",8519 => "01111101",8520 => "01011100",8521 => "11000101",8522 => "01110011",8523 => "00110010",8524 => "11010000",8525 => "11111101",8526 => "00110110",8527 => "11111001",8528 => "01000010",8529 => "00111011",8530 => "11000110",8531 => "00111110",8532 => "00000110",8533 => "01000001",8534 => "01010110",8535 => "00111011",8536 => "01010110",8537 => "10011001",8538 => "00111111",8539 => "00011011",8540 => "10111011",8541 => "11101000",8542 => "01101010",8543 => "11101110",8544 => "11110000",8545 => "11010001",8546 => "11010010",8547 => "10011001",8548 => "11100001",8549 => "01001000",8550 => "10110101",8551 => "11000000",8552 => "10011010",8553 => "11000101",8554 => "01110100",8555 => "11110001",8556 => "01100011",8557 => "01001001",8558 => "00111111",8559 => "01100011",8560 => "11101000",8561 => "00000110",8562 => "00010001",8563 => "01110001",8564 => "10101110",8565 => "01000000",8566 => "01001101",8567 => "11001011",8568 => "00111111",8569 => "10101110",8570 => "10111001",8571 => "00101110",8572 => "01011000",8573 => "00110111",8574 => "01010010",8575 => "00001100",8576 => "00101100",8577 => "00100111",8578 => "10001111",8579 => "01010001",8580 => "01110110",8581 => "11011111",8582 => "00011111",8583 => "11101101",8584 => "00111010",8585 => "01110001",8586 => "01011000",8587 => "01000000",8588 => "01101000",8589 => "11001001",8590 => "11001000",8591 => "00000001",8592 => "00000110",8593 => "00110011",8594 => "11010111",8595 => "10000110",8596 => "11000010",8597 => "00100000",8598 => "00101000",8599 => "00100011",8600 => "00110011",8601 => "01000001",8602 => "11100110",8603 => "11011000",8604 => "10000010",8605 => "01101001",8606 => "01111110",8607 => "00111011",8608 => "11000111",8609 => "00001100",8610 => "11111101",8611 => "10010011",8612 => "11011001",8613 => "11111000",8614 => "00001001",8615 => "10110010",8616 => "10110000",8617 => "01111100",8618 => "01100111",8619 => "10001000",8620 => "00111111",8621 => "10011011",8622 => "10100011",8623 => "11000010",8624 => "10000110",8625 => "11100001",8626 => "01001111",8627 => "11000110",8628 => "11101011",8629 => "01111111",8630 => "00101000",8631 => "10011100",8632 => "01110011",8633 => "01000001",8634 => "01101010",8635 => "10010110",8636 => "10011101",8637 => "00110001",8638 => "10010011",8639 => "11111100",8640 => "01010100",8641 => "00110101",8642 => "10001010",8643 => "10001101",8644 => "00110010",8645 => "10101111",8646 => "01011010",8647 => "01001000",8648 => "10100101",8649 => "11101000",8650 => "01010011",8651 => "00000101",8652 => "00100011",8653 => "00001001",8654 => "10010100",8655 => "11010110",8656 => "01000001",8657 => "00011100",8658 => "11001111",8659 => "00000011",8660 => "01001001",8661 => "01111100",8662 => "01111111",8663 => "01111100",8664 => "11101000",8665 => "01010110",8666 => "00100100",8667 => "01001000",8668 => "00001001",8669 => "01010110",8670 => "10110000",8671 => "01110110",8672 => "00100000",8673 => "00111111",8674 => "00010000",8675 => "11001000",8676 => "01001111",8677 => "00001101",8678 => "00001111",8679 => "11100000",8680 => "11110010",8681 => "11111111",8682 => "00100000",8683 => "11101001",8684 => "01010100",8685 => "00100001",8686 => "10001000",8687 => "11010010",8688 => "00110000",8689 => "01101010",8690 => "00001001",8691 => "01111101",8692 => "11110001",8693 => "01001101",8694 => "01000001",8695 => "01111110",8696 => "10000000",8697 => "00100111",8698 => "10111101",8699 => "00101011",8700 => "10101001",8701 => "11111111",8702 => "01110110",8703 => "00100011",8704 => "10010111",8705 => "01010110",8706 => "11000100",8707 => "00101010",8708 => "10011001",8709 => "11000110",8710 => "11000111",8711 => "01101001",8712 => "00111111",8713 => "01000101",8714 => "11110111",8715 => "11111000",8716 => "01101001",8717 => "10111101",8718 => "10110010",8719 => "10111010",8720 => "10011101",8721 => "00101011",8722 => "01010111",8723 => "01000011",8724 => "01111111",8725 => "01001110",8726 => "00001101",8727 => "01011110",8728 => "01110001",8729 => "11010000",8730 => "10100100",8731 => "01111111",8732 => "10111111",8733 => "10000100",8734 => "01111110",8735 => "11100111",8736 => "00011100",8737 => "10010010",8738 => "01010101",8739 => "01011100",8740 => "10111111",8741 => "11001111",8742 => "11101111",8743 => "11001101",8744 => "01101110",8745 => "10101101",8746 => "11111000",8747 => "11100010",8748 => "00000010",8749 => "00011111",8750 => "11000110",8751 => "10010010",8752 => "10010100",8753 => "10010101",8754 => "01110101",8755 => "00110011",8756 => "11001111",8757 => "01010001",8758 => "11110111",8759 => "00000110",8760 => "00011101",8761 => "00000001",8762 => "00010011",8763 => "11111111",8764 => "01001001",8765 => "11100011",8766 => "10001010",8767 => "10001010",8768 => "10100111",8769 => "11001001",8770 => "01011101",8771 => "00100110",8772 => "10101010",8773 => "01100001",8774 => "01001001",8775 => "11011101",8776 => "10110100",8777 => "10111100",8778 => "01010001",8779 => "00111101",8780 => "00110110",8781 => "00000001",8782 => "01111100",8783 => "11110100",8784 => "11000011",8785 => "11000011",8786 => "00011111",8787 => "11111011",8788 => "00011100",8789 => "11110011",8790 => "10000100",8791 => "10111001",8792 => "00101000",8793 => "00111101",8794 => "00000110",8795 => "11010000",8796 => "11100010",8797 => "11110001",8798 => "01110000",8799 => "00000011",8800 => "10111101",8801 => "00111101",8802 => "11011110",8803 => "10010100",8804 => "00000001",8805 => "00001001",8806 => "10011000",8807 => "10101111",8808 => "00110111",8809 => "11111101",8810 => "00100110",8811 => "00111011",8812 => "01101101",8813 => "01011011",8814 => "11101010",8815 => "10101100",8816 => "11110100",8817 => "00011111",8818 => "11011010",8819 => "01111100",8820 => "10100100",8821 => "11001111",8822 => "10010111",8823 => "00100100",8824 => "10101111",8825 => "01000100",8826 => "11000001",8827 => "00011010",8828 => "11101000",8829 => "11100111",8830 => "01110100",8831 => "01100100",8832 => "00100001",8833 => "01011011",8834 => "01100000",8835 => "01000101",8836 => "10111110",8837 => "10011100",8838 => "00101000",8839 => "01011001",8840 => "11111100",8841 => "11111010",8842 => "01010000",8843 => "10111011",8844 => "00001010",8845 => "00011010",8846 => "01111010",8847 => "01111100",8848 => "10111100",8849 => "01110000",8850 => "00000110",8851 => "11110001",8852 => "11110101",8853 => "10100101",8854 => "00001001",8855 => "11001100",8856 => "11110101",8857 => "10010010",8858 => "00001111",8859 => "01000101",8860 => "00101110",8861 => "00110000",8862 => "10110001",8863 => "00011000",8864 => "01000011",8865 => "11001111",8866 => "10000011",8867 => "01110111",8868 => "00110101",8869 => "01101001",8870 => "00110010",8871 => "00011000",8872 => "00001001",8873 => "00010000",8874 => "11010101",8875 => "01111100",8876 => "01000100",8877 => "11000111",8878 => "11100001",8879 => "11000111",8880 => "01001011",8881 => "11011010",8882 => "00000110",8883 => "00011100",8884 => "11000000",8885 => "11001011",8886 => "00011010",8887 => "00001001",8888 => "01001111",8889 => "10011000",8890 => "11010011",8891 => "11011111",8892 => "01010100",8893 => "10101111",8894 => "00010011",8895 => "11011001",8896 => "01111001",8897 => "00011111",8898 => "11011001",8899 => "11001111",8900 => "01001001",8901 => "11111110",8902 => "11101011",8903 => "00011010",8904 => "00100101",8905 => "11000000",8906 => "01001100",8907 => "11111000",8908 => "11011110",8909 => "00001101",8910 => "11100011",8911 => "11001111",8912 => "01100101",8913 => "00100100",8914 => "10100110",8915 => "11100111",8916 => "11100100",8917 => "10100111",8918 => "00111101",8919 => "01011110",8920 => "01100101",8921 => "00011101",8922 => "00000111",8923 => "00000010",8924 => "10111000",8925 => "00101011",8926 => "11110110",8927 => "10101101",8928 => "00111101",8929 => "10100110",8930 => "00000010",8931 => "11110010",8932 => "01001000",8933 => "00110101",8934 => "11101011",8935 => "01001110",8936 => "01001101",8937 => "00101010",8938 => "10001010",8939 => "10000101",8940 => "11000011",8941 => "11001110",8942 => "11010110",8943 => "01010000",8944 => "00100001",8945 => "11100110",8946 => "10100011",8947 => "10010110",8948 => "10110110",8949 => "11101010",8950 => "11001111",8951 => "10000110",8952 => "10110101",8953 => "11000100",8954 => "10001011",8955 => "10110111",8956 => "00001010",8957 => "00101011",8958 => "01010001",8959 => "00011010",8960 => "01001101",8961 => "00000111",8962 => "01010011",8963 => "10110001",8964 => "11100011",8965 => "01000100",8966 => "00100101",8967 => "00001000",8968 => "10011010",8969 => "00000001",8970 => "10001110",8971 => "00110000",8972 => "00011001",8973 => "10010110",8974 => "01000001",8975 => "01110111",8976 => "11110001",8977 => "00110110",8978 => "11011011",8979 => "01011100",8980 => "00000100",8981 => "00000010",8982 => "11100011",8983 => "01001010",8984 => "01010101",8985 => "01011011",8986 => "00010011",8987 => "10101010",8988 => "11010100",8989 => "11010011",8990 => "10011110",8991 => "10110100",8992 => "10110101",8993 => "00011110",8994 => "00001001",8995 => "00111000",8996 => "01001110",8997 => "11110011",8998 => "01010110",8999 => "10010110",9000 => "01011011",9001 => "01010100",9002 => "10100000",9003 => "00100101",9004 => "11111101",9005 => "11111100",9006 => "01001011",9007 => "10111000",9008 => "01100100",9009 => "11110110",9010 => "10010110",9011 => "00111100",9012 => "11100100",9013 => "11111100",9014 => "01011100",9015 => "00101110",9016 => "11110101",9017 => "10100101",9018 => "00010001",9019 => "01111101",9020 => "01100110",9021 => "01111111",9022 => "11010000",9023 => "01000001",9024 => "00110101",9025 => "00111101",9026 => "01110101",9027 => "11111110",9028 => "10100010",9029 => "01010010",9030 => "10001001",9031 => "00010110",9032 => "01010111",9033 => "10000011",9034 => "00010001",9035 => "11100111",9036 => "01001000",9037 => "01100100",9038 => "01100100",9039 => "00110111",9040 => "11111100",9041 => "11000100",9042 => "01010110",9043 => "10110010",9044 => "11010010",9045 => "11011111",9046 => "01001000",9047 => "01100111",9048 => "00101100",9049 => "01000110",9050 => "01001111",9051 => "11000100",9052 => "11001011",9053 => "11011111",9054 => "01011011",9055 => "11001100",9056 => "01100110",9057 => "11111001",9058 => "00111011",9059 => "10110001",9060 => "10100000",9061 => "10100101",9062 => "00110111",9063 => "01110011",9064 => "01111100",9065 => "11110000",9066 => "11101111",9067 => "11001101",9068 => "00100001",9069 => "11010110",9070 => "10001100",9071 => "10011010",9072 => "00001110",9073 => "00010001",9074 => "01100001",9075 => "11011001",9076 => "10101110",9077 => "00100101",9078 => "00100110",9079 => "01000111",9080 => "00000110",9081 => "01100001",9082 => "01011011",9083 => "10010011",9084 => "00101101",9085 => "11011011",9086 => "10011001",9087 => "10010001",9088 => "10011111",9089 => "10000100",9090 => "10001001",9091 => "11011101",9092 => "10100101",9093 => "01110110",9094 => "01010011",9095 => "10100111",9096 => "11110111",9097 => "10101010",9098 => "00011010",9099 => "01100001",9100 => "10110011",9101 => "10111000",9102 => "10000011",9103 => "10001110",9104 => "00111010",9105 => "11001110",9106 => "11110011",9107 => "10001110",9108 => "11100100",9109 => "01100010",9110 => "01000000",9111 => "00110011",9112 => "01011100",9113 => "01000101",9114 => "11010000",9115 => "00110011",9116 => "00101110",9117 => "00110001",9118 => "00111001",9119 => "01000111",9120 => "00011000",9121 => "10110111",9122 => "00100100",9123 => "00011111",9124 => "01010000",9125 => "11101001",9126 => "10100111",9127 => "11011000",9128 => "11111101",9129 => "00111001",9130 => "10100001",9131 => "01011100",9132 => "11000100",9133 => "00000111",9134 => "01100000",9135 => "00001111",9136 => "10111111",9137 => "11111110",9138 => "01111011",9139 => "10010110",9140 => "10111001",9141 => "01010100",9142 => "01110101",9143 => "01100100",9144 => "11011111",9145 => "10010011",9146 => "00010101",9147 => "11000010",9148 => "00111110",9149 => "11101111",9150 => "11000101",9151 => "00011001",9152 => "10001111",9153 => "11001111",9154 => "10100100",9155 => "10101110",9156 => "11011110",9157 => "01000010",9158 => "01100011",9159 => "11110100",9160 => "10111001",9161 => "10111100",9162 => "10010100",9163 => "11010111",9164 => "00110101",9165 => "10011000",9166 => "11111101",9167 => "01111010",9168 => "11001000",9169 => "11110001",9170 => "10011100",9171 => "00001111",9172 => "11111111",9173 => "01100001",9174 => "01011001",9175 => "11001101",9176 => "10101000",9177 => "00011101",9178 => "11001110",9179 => "11011001",9180 => "01010101",9181 => "10011111",9182 => "11011000",9183 => "11011000",9184 => "10001011",9185 => "01101111",9186 => "00101010",9187 => "00011010",9188 => "01011011",9189 => "10010110",9190 => "11010001",9191 => "10110000",9192 => "11010001",9193 => "00010110",9194 => "10000110",9195 => "00000001",9196 => "00010110",9197 => "00111000",9198 => "11001101",9199 => "10001010",9200 => "11011101",9201 => "11011011",9202 => "00100100",9203 => "01110110",9204 => "11100110",9205 => "01101010",9206 => "01101001",9207 => "10000110",9208 => "00111110",9209 => "01010011",9210 => "10010110",9211 => "11100101",9212 => "11010011",9213 => "00010010",9214 => "10111011",9215 => "11001101",9216 => "00000000",9217 => "11001000",9218 => "11110011",9219 => "11010000",9220 => "10000001",9221 => "10111010",9222 => "00001011",9223 => "11111010",9224 => "01100110",9225 => "10111110",9226 => "00011000",9227 => "11010100",9228 => "00001011",9229 => "00100110",9230 => "01000000",9231 => "01010101",9232 => "11100000",9233 => "00000111",9234 => "11010011",9235 => "10110111",9236 => "11011001",9237 => "01011011",9238 => "11001010",9239 => "00100010",9240 => "10101100",9241 => "10011011",9242 => "01110101",9243 => "11011010",9244 => "00000100",9245 => "00110100",9246 => "00011000",9247 => "11111101",9248 => "01101011",9249 => "11110011",9250 => "11010110",9251 => "01101111",9252 => "01101110",9253 => "11011111",9254 => "00010111",9255 => "00111100",9256 => "01001000",9257 => "01100100",9258 => "10000011",9259 => "00000010",9260 => "00100111",9261 => "10001100",9262 => "00010000",9263 => "11011111",9264 => "11000011",9265 => "11001100",9266 => "10100001",9267 => "00111110",9268 => "10010111",9269 => "10111010",9270 => "10111100",9271 => "01010110",9272 => "11101000",9273 => "10101010",9274 => "11010010",9275 => "11000001",9276 => "10011001",9277 => "10110111",9278 => "00010001",9279 => "10000000",9280 => "01110101",9281 => "01111100",9282 => "01111000",9283 => "10101011",9284 => "00001111",9285 => "00100101",9286 => "10110101",9287 => "01010001",9288 => "01010001",9289 => "10110111",9290 => "00011101",9291 => "10010100",9292 => "01001010",9293 => "00000101",9294 => "00001000",9295 => "00010111",9296 => "10110100",9297 => "01101001",9298 => "10000001",9299 => "00111011",9300 => "00111110",9301 => "01100110",9302 => "01110010",9303 => "11101100",9304 => "00110101",9305 => "11100110",9306 => "01000100",9307 => "00011010",9308 => "10011101",9309 => "00101010",9310 => "10001101",9311 => "01000110",9312 => "01010010",9313 => "01100010",9314 => "10011011",9315 => "01011001",9316 => "01110011",9317 => "11111101",9318 => "10110101",9319 => "00000111",9320 => "00001011",9321 => "10011101",9322 => "01111100",9323 => "01011111",9324 => "10001110",9325 => "10111011",9326 => "00010011",9327 => "01001110",9328 => "00000011",9329 => "00011001",9330 => "11110110",9331 => "00110001",9332 => "10010011",9333 => "00110001",9334 => "11000100",9335 => "11100110",9336 => "10011000",9337 => "11000010",9338 => "00101111",9339 => "10001110",9340 => "01110011",9341 => "00100110",9342 => "10000001",9343 => "10100110",9344 => "11011000",9345 => "11010110",9346 => "10101000",9347 => "10010101",9348 => "11110101",9349 => "00101110",9350 => "00101001",9351 => "01001101",9352 => "10000000",9353 => "10010011",9354 => "11110001",9355 => "00110011",9356 => "00000000",9357 => "00011100",9358 => "00001011",9359 => "00000110",9360 => "11000011",9361 => "11000100",9362 => "01111111",9363 => "11001000",9364 => "00000111",9365 => "10101101",9366 => "11100011",9367 => "10111100",9368 => "11100001",9369 => "01010111",9370 => "10110110",9371 => "10111101",9372 => "10111101",9373 => "01101000",9374 => "01001110",9375 => "11101101",9376 => "01001110",9377 => "10011100",9378 => "01011110",9379 => "11110001",9380 => "11011101",9381 => "01011110",9382 => "11011110",9383 => "00011101",9384 => "01100011",9385 => "11101111",9386 => "10010100",9387 => "10101010",9388 => "01110100",9389 => "00001000",9390 => "00010000",9391 => "01100110",9392 => "11000111",9393 => "11000010",9394 => "11110010",9395 => "10000000",9396 => "11000011",9397 => "11110010",9398 => "01000001",9399 => "01010110",9400 => "11011000",9401 => "10000100",9402 => "01000010",9403 => "11101001",9404 => "00011010",9405 => "10001010",9406 => "01101110",9407 => "00111010",9408 => "10100111",9409 => "11100001",9410 => "11111000",9411 => "10011111",9412 => "11010100",9413 => "10011101",9414 => "00101001",9415 => "10011000",9416 => "10000101",9417 => "10000001",9418 => "00001110",9419 => "00000110",9420 => "00001000",9421 => "00000111",9422 => "00100111",9423 => "00101001",9424 => "11101111",9425 => "00110011",9426 => "01111110",9427 => "01110110",9428 => "00111000",9429 => "11000100",9430 => "00011101",9431 => "00010111",9432 => "10100010",9433 => "10101001",9434 => "01001111",9435 => "00011101",9436 => "00000100",9437 => "01111101",9438 => "11101001",9439 => "11010000",9440 => "00000001",9441 => "00100001",9442 => "00101100",9443 => "11100110",9444 => "10101010",9445 => "10000000",9446 => "10000111",9447 => "10010001",9448 => "01000001",9449 => "11000100",9450 => "11011101",9451 => "00000110",9452 => "11111111",9453 => "10101001",9454 => "10000011",9455 => "10110111",9456 => "10010110",9457 => "11000000",9458 => "11100001",9459 => "01010110",9460 => "10110011",9461 => "11011000",9462 => "01101110",9463 => "01000100",9464 => "10001000",9465 => "11000001",9466 => "10111111",9467 => "11010110",9468 => "01101101",9469 => "11011010",9470 => "11111011",9471 => "11001110",9472 => "11111100",9473 => "11010100",9474 => "00111000",9475 => "00101011",9476 => "00010110",9477 => "11001001",9478 => "10000001",9479 => "01111011",9480 => "00101011",9481 => "11010010",9482 => "11111001",9483 => "01111100",9484 => "10101110",9485 => "11001001",9486 => "11100111",9487 => "11000000",9488 => "00111110",9489 => "01111001",9490 => "10110101",9491 => "11011100",9492 => "11011010",9493 => "10100100",9494 => "00101000",9495 => "01111000",9496 => "00100100",9497 => "01101011",9498 => "00111000",9499 => "11010010",9500 => "10101110",9501 => "11110001",9502 => "11100011",9503 => "10110001",9504 => "10001011",9505 => "10111111",9506 => "01000111",9507 => "10001010",9508 => "11011010",9509 => "10011001",9510 => "00111111",9511 => "10100001",9512 => "11001110",9513 => "11000111",9514 => "10101110",9515 => "11110100",9516 => "01100010",9517 => "10011100",9518 => "11110110",9519 => "10101001",9520 => "00001101",9521 => "11111101",9522 => "10001111",9523 => "10111000",9524 => "01111000",9525 => "01010101",9526 => "11010100",9527 => "11011000",9528 => "01001111",9529 => "10000110",9530 => "11111011",9531 => "01000001",9532 => "10111110",9533 => "10001011",9534 => "11000010",9535 => "11000001",9536 => "00101010",9537 => "01011111",9538 => "01011110",9539 => "00000011",9540 => "11111001",9541 => "10101001",9542 => "11100010",9543 => "00011101",9544 => "00111101",9545 => "11000101",9546 => "00001001",9547 => "10101011",9548 => "00011101",9549 => "11001111",9550 => "01000011",9551 => "01110011",9552 => "00101000",9553 => "01101001",9554 => "01011001",9555 => "11110101",9556 => "01010001",9557 => "10101001",9558 => "01111101",9559 => "00000101",9560 => "01110000",9561 => "01100001",9562 => "10100001",9563 => "01011111",9564 => "11010010",9565 => "10001110",9566 => "00101010",9567 => "10110111",9568 => "00011001",9569 => "01001100",9570 => "11111010",9571 => "00000100",9572 => "01100011",9573 => "10101010",9574 => "11010001",9575 => "01110000",9576 => "01110100",9577 => "01001000",9578 => "01111100",9579 => "10100000",9580 => "01100000",9581 => "00111100",9582 => "01111011",9583 => "01100000",9584 => "00111001",9585 => "00010001",9586 => "11000001",9587 => "10111011",9588 => "10000010",9589 => "00111000",9590 => "01000110",9591 => "10101010",9592 => "10000110",9593 => "10010001",9594 => "10110100",9595 => "00000001",9596 => "00100110",9597 => "10011001",9598 => "01001101",9599 => "00000010",9600 => "10001011",9601 => "01000010",9602 => "11110000",9603 => "01010010",9604 => "10011111",9605 => "01010010",9606 => "10110011",9607 => "01010001",9608 => "00010011",9609 => "00001110",9610 => "01101111",9611 => "01111100",9612 => "01111010",9613 => "11110000",9614 => "11000101",9615 => "10110110",9616 => "00100100",9617 => "11110010",9618 => "00101010",9619 => "10110000",9620 => "00101000",9621 => "11100000",9622 => "10001001",9623 => "11111001",9624 => "11001101",9625 => "11000101",9626 => "10010000",9627 => "00110101",9628 => "10111110",9629 => "01001100",9630 => "00000101",9631 => "11000101",9632 => "01010011",9633 => "00100101",9634 => "11110100",9635 => "11001011",9636 => "01110101",9637 => "00111010",9638 => "11001110",9639 => "01101011",9640 => "00110101",9641 => "00011001",9642 => "11100110",9643 => "01100110",9644 => "01011111",9645 => "01001011",9646 => "00100101",9647 => "11101001",9648 => "00010010",9649 => "11101001",9650 => "11100011",9651 => "10011110",9652 => "01001111",9653 => "11011110",9654 => "11010001",9655 => "01111011",9656 => "00110110",9657 => "01010111",9658 => "11010100",9659 => "11011000",9660 => "10010101",9661 => "01011001",9662 => "00000100",9663 => "00001101",9664 => "11011001",9665 => "11011111",9666 => "00001000",9667 => "00010011",9668 => "00010001",9669 => "11011001",9670 => "01101111",9671 => "10001011",9672 => "10110111",9673 => "10011101",9674 => "11001010",9675 => "00110010",9676 => "10100001",9677 => "00110000",9678 => "01110100",9679 => "10111010",9680 => "01110000",9681 => "00011100",9682 => "00101111",9683 => "00100001",9684 => "00110000",9685 => "01111111",9686 => "00100010",9687 => "11100111",9688 => "00100000",9689 => "10010111",9690 => "11101011",9691 => "11011010",9692 => "01100101",9693 => "11001000",9694 => "10110100",9695 => "00010100",9696 => "10011101",9697 => "10000000",9698 => "00100100",9699 => "11001111",9700 => "11011110",9701 => "01111011",9702 => "00110110",9703 => "11010101",9704 => "10111111",9705 => "10101000",9706 => "00000110",9707 => "11101101",9708 => "01000001",9709 => "00111001",9710 => "10101100",9711 => "11010000",9712 => "01111001",9713 => "00011010",9714 => "11110011",9715 => "10100010",9716 => "11110011",9717 => "00011111",9718 => "10000101",9719 => "11110101",9720 => "00111101",9721 => "00111001",9722 => "01011011",9723 => "10011001",9724 => "01110010",9725 => "01000100",9726 => "11000000",9727 => "00001110",9728 => "10110000",9729 => "10101001",9730 => "11010110",9731 => "10100111",9732 => "01101010",9733 => "10110010",9734 => "00110001",9735 => "10011011",9736 => "11111110",9737 => "11101000",9738 => "01100010",9739 => "01110100",9740 => "10111111",9741 => "10110101",9742 => "01111000",9743 => "00110110",9744 => "11110011",9745 => "00111010",9746 => "11101000",9747 => "00010011",9748 => "01100010",9749 => "11001101",9750 => "11010111",9751 => "01101010",9752 => "11100111",9753 => "01111011",9754 => "10001110",9755 => "00101100",9756 => "11011011",9757 => "01010100",9758 => "01101110",9759 => "01010110",9760 => "10001000",9761 => "01010100",9762 => "01101101",9763 => "10100000",9764 => "10010101",9765 => "10011110",9766 => "01111011",9767 => "01000010",9768 => "11000110",9769 => "01001001",9770 => "01101001",9771 => "01101100",9772 => "11010011",9773 => "00111101",9774 => "10110100",9775 => "11010100",9776 => "10000110",9777 => "00001011",9778 => "01110111",9779 => "11101111",9780 => "10000101",9781 => "11000011",9782 => "00110011",9783 => "11100001",9784 => "00111101",9785 => "10100001",9786 => "01110000",9787 => "11111001",9788 => "11110110",9789 => "10110011",9790 => "10111010",9791 => "10011110",9792 => "00101110",9793 => "00110010",9794 => "11110000",9795 => "00011110",9796 => "00001111",9797 => "11010011",9798 => "01011111",9799 => "01000101",9800 => "01101110",9801 => "11110001",9802 => "01111000",9803 => "10010101",9804 => "01111011",9805 => "01010110",9806 => "11011001",9807 => "00010101",9808 => "00100001",9809 => "01010111",9810 => "10010001",9811 => "11010011",9812 => "01111101",9813 => "10101110",9814 => "11010100",9815 => "11001001",9816 => "00110000",9817 => "00010001",9818 => "10110101",9819 => "01101001",9820 => "00001011",9821 => "11010001",9822 => "11110001",9823 => "01101010",9824 => "11001101",9825 => "00110011",9826 => "01010000",9827 => "00000111",9828 => "10110011",9829 => "01010001",9830 => "00010000",9831 => "01101110",9832 => "00110111",9833 => "00001111",9834 => "10011111",9835 => "00111001",9836 => "01101001",9837 => "11100111",9838 => "01001110",9839 => "11101101",9840 => "10010001",9841 => "00100000",9842 => "00001101",9843 => "10110100",9844 => "00110100",9845 => "00010000",9846 => "11000100",9847 => "00011110",9848 => "10011010",9849 => "10101010",9850 => "00011111",9851 => "00100100",9852 => "00110101",9853 => "00111110",9854 => "10100010",9855 => "11010011",9856 => "00001100",9857 => "01001010",9858 => "10100111",9859 => "01100000",9860 => "01101110",9861 => "10100100",9862 => "00111011",9863 => "01001001",9864 => "11111011",9865 => "00111110",9866 => "01101111",9867 => "10001111",9868 => "01111010",9869 => "00010101",9870 => "10111001",9871 => "00000001",9872 => "11000000",9873 => "10000101",9874 => "00010010",9875 => "01101101",9876 => "11001010",9877 => "10111101",9878 => "10110010",9879 => "11001100",9880 => "10101100",9881 => "11000010",9882 => "11100000",9883 => "10011010",9884 => "10111110",9885 => "01111010",9886 => "10011001",9887 => "01001101",9888 => "11010101",9889 => "11100101",9890 => "10010100",9891 => "11000001",9892 => "00110001",9893 => "11101111",9894 => "11001111",9895 => "00000110",9896 => "01100101",9897 => "01001000",9898 => "01100010",9899 => "11000000",9900 => "11000001",9901 => "01011111",9902 => "11001111",9903 => "11001000",9904 => "00100110",9905 => "00001111",9906 => "11110111",9907 => "11111110",9908 => "01111110",9909 => "10010000",9910 => "01110110",9911 => "00011111",9912 => "10110111",9913 => "01101001",9914 => "01101010",9915 => "11000111",9916 => "10011000",9917 => "01101101",9918 => "11110110",9919 => "01010001",9920 => "01001001",9921 => "00110010",9922 => "10011100",9923 => "00101101",9924 => "11010001",9925 => "01111110",9926 => "11001001",9927 => "00010000",9928 => "11001101",9929 => "10000010",9930 => "00010000",9931 => "01011001",9932 => "11100100",9933 => "10001000",9934 => "10010100",9935 => "10000110",9936 => "10110111",9937 => "11111011",9938 => "00000100",9939 => "00001011",9940 => "00110001",9941 => "10000100",9942 => "01001101",9943 => "00111100",9944 => "11101111",9945 => "10001010",9946 => "01101000",9947 => "11001101",9948 => "10001001",9949 => "00100111",9950 => "00000110",9951 => "10000100",9952 => "01000001",9953 => "11100000",9954 => "00000010",9955 => "01010110",9956 => "10111000",9957 => "10100010",9958 => "10111101",9959 => "10000111",9960 => "00000110",9961 => "00111001",9962 => "00111100",9963 => "11011100",9964 => "10010001",9965 => "11101000",9966 => "11111101",9967 => "11000001",9968 => "01010111",9969 => "11110101",9970 => "01000000",9971 => "10111011",9972 => "01100010",9973 => "01100011",9974 => "11111101",9975 => "01111111",9976 => "10111101",9977 => "00000111",9978 => "00110101",9979 => "01011010",9980 => "11101101",9981 => "01110000",9982 => "11100011",9983 => "11010001",9984 => "00000110",9985 => "11000110",9986 => "00100001",9987 => "10000010",9988 => "10100010",9989 => "01000100",9990 => "01110000",9991 => "11001010",9992 => "11111101",9993 => "01100111",9994 => "10000111",9995 => "00101010",9996 => "10111000",9997 => "10010010",9998 => "00010111",9999 => "10000000",10000 => "01111100",10001 => "11001011",10002 => "10110010",10003 => "00001110",10004 => "11101101",10005 => "10110011",10006 => "10100110",10007 => "00000010",10008 => "11011001",10009 => "11011101",10010 => "11111100",10011 => "10001010",10012 => "10100001",10013 => "10100110",10014 => "01000010",10015 => "11100001",10016 => "01010000",10017 => "11111110",10018 => "01011000",10019 => "10111001",10020 => "10010001",10021 => "00001000",10022 => "01110010",10023 => "00101001",10024 => "11010101",10025 => "10110010",10026 => "10011110",10027 => "10001101",10028 => "10010000",10029 => "00010001",10030 => "11011111",10031 => "11101110",10032 => "00010011",10033 => "10101000",10034 => "00011001",10035 => "00101001",10036 => "01101000",10037 => "01010101",10038 => "10011010",10039 => "00010000",10040 => "10110011",10041 => "11101111",10042 => "11000110",10043 => "01000111",10044 => "00100011",10045 => "11101110",10046 => "11110000",10047 => "11000000",10048 => "10001110",10049 => "01101000",10050 => "10011111",10051 => "00101101",10052 => "11011011",10053 => "01100111",10054 => "00011000",10055 => "11001001",10056 => "11000001",10057 => "00100101",10058 => "11011011",10059 => "11101010",10060 => "11111011",10061 => "10010000",10062 => "01000111",10063 => "01001010",10064 => "11100010",10065 => "10110111",10066 => "10000101",10067 => "10110100",10068 => "10010111",10069 => "00000011",10070 => "01011011",10071 => "00111010",10072 => "11100111",10073 => "00110011",10074 => "00000000",10075 => "11000111",10076 => "11110101",10077 => "00110010",10078 => "11111011",10079 => "01101011",10080 => "00010011",10081 => "10000011",10082 => "11001001",10083 => "11110001",10084 => "11000111",10085 => "10010111",10086 => "01110101",10087 => "01101101",10088 => "10010011",10089 => "00101001",10090 => "01100010",10091 => "00110011",10092 => "10001110",10093 => "01111100",10094 => "01000100",10095 => "10011010",10096 => "00011101",10097 => "00000010",10098 => "00111000",10099 => "01101010",10100 => "10111000",10101 => "01111000",10102 => "00100001",10103 => "11010001",10104 => "10110000",10105 => "11100110",10106 => "11100110",10107 => "00111001",10108 => "10100000",10109 => "11011001",10110 => "10111000",10111 => "01010110",10112 => "11110010",10113 => "01001110",10114 => "00101100",10115 => "10011100",10116 => "11111001",10117 => "00011011",10118 => "11000111",10119 => "01101111",10120 => "00111010",10121 => "11101011",10122 => "01111100",10123 => "11011001",10124 => "11100010",10125 => "01001101",10126 => "11111111",10127 => "10010010",10128 => "11000111",10129 => "11101001",10130 => "00100111",10131 => "10110000",10132 => "11010110",10133 => "00011101",10134 => "01010001",10135 => "10110000",10136 => "10010110",10137 => "11111011",10138 => "00001101",10139 => "11100110",10140 => "11000011",10141 => "10100010",10142 => "00110101",10143 => "01010110",10144 => "10011000",10145 => "10101110",10146 => "00011101",10147 => "10001000",10148 => "01011101",10149 => "01100011",10150 => "00000000",10151 => "00111000",10152 => "11010100",10153 => "01101101",10154 => "10001011",10155 => "11110010",10156 => "01010000",10157 => "11000000",10158 => "11111100",10159 => "00101101",10160 => "00001011",10161 => "11111110",10162 => "11100001",10163 => "01110011",10164 => "11101001",10165 => "01010001",10166 => "11100110",10167 => "10010111",10168 => "11001100",10169 => "10001001",10170 => "10010100",10171 => "10100000",10172 => "11000001",10173 => "01110110",10174 => "10000101",10175 => "10110011",10176 => "10001110",10177 => "01010110",10178 => "10001101",10179 => "00000110",10180 => "10110110",10181 => "10001101",10182 => "00111011",10183 => "10110000",10184 => "01110000",10185 => "11010010",10186 => "01001011",10187 => "00001111",10188 => "10101010",10189 => "01101111",10190 => "11010001",10191 => "01100011",10192 => "11100000",10193 => "11100101",10194 => "11000010",10195 => "11000111",10196 => "10000100",10197 => "10000011",10198 => "00111001",10199 => "10110101",10200 => "10111000",10201 => "01010101",10202 => "11100001",10203 => "11000100",10204 => "11000011",10205 => "01110010",10206 => "11011001",10207 => "01101100",10208 => "11111010",10209 => "01111011",10210 => "11010110",10211 => "01111011",10212 => "11100100",10213 => "10110111",10214 => "11100010",10215 => "00111011",10216 => "01110001",10217 => "11101110",10218 => "11101000",10219 => "10111100",10220 => "00010100",10221 => "11101001",10222 => "10000100",10223 => "00100101",10224 => "01101100",10225 => "00011010",10226 => "11000010",10227 => "01011101",10228 => "11000000",10229 => "01110101",10230 => "11000111",10231 => "00001011",10232 => "11010011",10233 => "11100111",10234 => "01110100",10235 => "11001010",10236 => "00111111",10237 => "10110110",10238 => "00110011",10239 => "00010010",10240 => "01111101",10241 => "11011011",10242 => "10011100",10243 => "00001110",10244 => "10001101",10245 => "11101000",10246 => "01100010",10247 => "11100111",10248 => "11010001",10249 => "11010001",10250 => "01011011",10251 => "00111010",10252 => "11101000",10253 => "00111010",10254 => "00100001",10255 => "11011110",10256 => "01000110",10257 => "00011000",10258 => "11100010",10259 => "10101011",10260 => "01111001",10261 => "11010100",10262 => "00011110",10263 => "11010110",10264 => "10110111",10265 => "00000111",10266 => "11001011",10267 => "10010101",10268 => "11101111",10269 => "00110001",10270 => "00000111",10271 => "10000101",10272 => "10001001",10273 => "11101101",10274 => "10100111",10275 => "01100100",10276 => "11000101",10277 => "00110110",10278 => "01011111",10279 => "01100100",10280 => "00010101",10281 => "11110000",10282 => "10011111",10283 => "10111101",10284 => "00111100",10285 => "00111111",10286 => "00101100",10287 => "01010100",10288 => "10001010",10289 => "01011111",10290 => "00100111",10291 => "11010110",10292 => "10110101",10293 => "01001101",10294 => "10101001",10295 => "00001100",10296 => "01111011",10297 => "10110110",10298 => "00001010",10299 => "01101100",10300 => "11001111",10301 => "01101000",10302 => "11100111",10303 => "00110110",10304 => "10010010",10305 => "00100011",10306 => "00001010",10307 => "00111100",10308 => "01001100",10309 => "00100011",10310 => "00111010",10311 => "10110100",10312 => "10011011",10313 => "10001111",10314 => "11011011",10315 => "01010111",10316 => "00111101",10317 => "01011011",10318 => "00000110",10319 => "11011111",10320 => "10001010",10321 => "10111111",10322 => "01100100",10323 => "01001001",10324 => "00111001",10325 => "10100111",10326 => "11010100",10327 => "10011111",10328 => "01010010",10329 => "10111010",10330 => "01111111",10331 => "01001111",10332 => "01001001",10333 => "00100010",10334 => "10101011",10335 => "10011111",10336 => "00001011",10337 => "11101001",10338 => "11000100",10339 => "10110001",10340 => "10101110",10341 => "01101010",10342 => "01100110",10343 => "00111111",10344 => "01111001",10345 => "10001111",10346 => "10010111",10347 => "00011100",10348 => "11100001",10349 => "10110111",10350 => "11011001",10351 => "10100000",10352 => "00011110",10353 => "10101111",10354 => "01011110",10355 => "10100110",10356 => "11010100",10357 => "10111001",10358 => "11110101",10359 => "00001001",10360 => "10100110",10361 => "00000010",10362 => "11110000",10363 => "10111100",10364 => "01110111",10365 => "11111100",10366 => "10000010",10367 => "10010011",10368 => "01101110",10369 => "00011000",10370 => "10010100",10371 => "01100011",10372 => "10100011",10373 => "11110011",10374 => "01100010",10375 => "01011000",10376 => "01100111",10377 => "11110011",10378 => "00000110",10379 => "10010100",10380 => "01111111",10381 => "10001010",10382 => "01011000",10383 => "00011010",10384 => "00101111",10385 => "01110001",10386 => "11100011",10387 => "00111111",10388 => "00001110",10389 => "10010110",10390 => "01010100",10391 => "01111110",10392 => "00000110",10393 => "00110011",10394 => "00100101",10395 => "01011101",10396 => "10011101",10397 => "00111110",10398 => "00100000",10399 => "00101101",10400 => "10010100",10401 => "10000001",10402 => "01011010",10403 => "00000100",10404 => "11000000",10405 => "11111101",10406 => "00101000",10407 => "10111001",10408 => "10101111",10409 => "10100100",10410 => "00110111",10411 => "00111001",10412 => "00011010",10413 => "01101101",10414 => "01100010",10415 => "10011010",10416 => "11110010",10417 => "10010100",10418 => "10100011",10419 => "10111101",10420 => "11111110",10421 => "11101110",10422 => "11101101",10423 => "01111011",10424 => "00000100",10425 => "11011000",10426 => "11100011",10427 => "10010101",10428 => "01000000",10429 => "01100000",10430 => "00111110",10431 => "00000010",10432 => "11001110",10433 => "10000111",10434 => "01000001",10435 => "01011011",10436 => "00000000",10437 => "00101110",10438 => "01001010",10439 => "00101110",10440 => "00100011",10441 => "00101010",10442 => "01101101",10443 => "10001011",10444 => "10000110",10445 => "00100000",10446 => "11010100",10447 => "10111000",10448 => "01111011",10449 => "10011010",10450 => "11000000",10451 => "01010100",10452 => "11001000",10453 => "01111010",10454 => "00100010",10455 => "01100011",10456 => "01011101",10457 => "00101000",10458 => "10010101",10459 => "00100000",10460 => "00011100",10461 => "11001110",10462 => "00100000",10463 => "10110011",10464 => "00001111",10465 => "10110010",10466 => "10101110",10467 => "01010000",10468 => "00100101",10469 => "00111010",10470 => "11000100",10471 => "11100111",10472 => "00001100",10473 => "10000010",10474 => "10111110",10475 => "11111110",10476 => "00100010",10477 => "00110010",10478 => "11001100",10479 => "00001100",10480 => "01100110",10481 => "10100001",10482 => "11110000",10483 => "00111001",10484 => "10011111",10485 => "00010011",10486 => "00111101",10487 => "01100010",10488 => "01111001",10489 => "11110101",10490 => "10011000",10491 => "10110100",10492 => "00111111",10493 => "11000000",10494 => "11011001",10495 => "00110000",10496 => "11110011",10497 => "10100000",10498 => "10001001",10499 => "10100001",10500 => "01010011",10501 => "01001100",10502 => "00111110",10503 => "11001101",10504 => "01101101",10505 => "11100001",10506 => "10110000",10507 => "11011111",10508 => "11110011",10509 => "01101101",10510 => "11011011",10511 => "01100000",10512 => "01000010",10513 => "11011101",10514 => "10111111",10515 => "10111100",10516 => "01110011",10517 => "00110100",10518 => "11001101",10519 => "10111110",10520 => "11110110",10521 => "01100011",10522 => "10001100",10523 => "01111001",10524 => "10010110",10525 => "10001111",10526 => "10100101",10527 => "11011111",10528 => "00110010",10529 => "10111001",10530 => "11001111",10531 => "10011111",10532 => "01010101",10533 => "10000111",10534 => "11011110",10535 => "10110001",10536 => "01101100",10537 => "01010100",10538 => "00101001",10539 => "11111010",10540 => "10010011",10541 => "01101110",10542 => "01001111",10543 => "01001000",10544 => "11011100",10545 => "10101111",10546 => "00101000",10547 => "01010111",10548 => "11001001",10549 => "01010011",10550 => "11101110",10551 => "10110110",10552 => "10111100",10553 => "01001011",10554 => "01101111",10555 => "11111101",10556 => "01100000",10557 => "10000001",10558 => "01100011",10559 => "00010111",10560 => "11000010",10561 => "11001000",10562 => "11000100",10563 => "00111100",10564 => "01010011",10565 => "11100110",10566 => "11101011",10567 => "00111111",10568 => "10000101",10569 => "10100111",10570 => "01110111",10571 => "00110100",10572 => "00010110",10573 => "00101000",10574 => "01111000",10575 => "00010000",10576 => "11011111",10577 => "10111110",10578 => "10111011",10579 => "01001100",10580 => "10001100",10581 => "10010000",10582 => "10010110",10583 => "11011010",10584 => "01101111",10585 => "10110100",10586 => "10100101",10587 => "11110110",10588 => "01010000",10589 => "00111001",10590 => "00001000",10591 => "11000001",10592 => "01101011",10593 => "00110111",10594 => "00011010",10595 => "11010001",10596 => "11011000",10597 => "10001101",10598 => "00101000",10599 => "00101100",10600 => "11011001",10601 => "00101100",10602 => "11010100",10603 => "10001110",10604 => "00100101",10605 => "01000111",10606 => "11110010",10607 => "00100100",10608 => "01101110",10609 => "10010110",10610 => "00100100",10611 => "01101001",10612 => "00111101",10613 => "00000101",10614 => "11011100",10615 => "11001100",10616 => "00110011",10617 => "00010011",10618 => "01011010",10619 => "01101111",10620 => "01001101",10621 => "10000110",10622 => "11101011",10623 => "00100000",10624 => "11110111",10625 => "11000110",10626 => "01010111",10627 => "01010110",10628 => "10011111",10629 => "00110000",10630 => "10000000",10631 => "01011100",10632 => "01100001",10633 => "11110011",10634 => "01100010",10635 => "11000100",10636 => "10100000",10637 => "00000101",10638 => "01101100",10639 => "10110110",10640 => "11110110",10641 => "10111011",10642 => "10110110",10643 => "00100101",10644 => "11101011",10645 => "01011100",10646 => "11101000",10647 => "00011001",10648 => "01101010",10649 => "01110011",10650 => "01001111",10651 => "01000111",10652 => "01110110",10653 => "10010010",10654 => "10110000",10655 => "00101001",10656 => "01110100",10657 => "10001010",10658 => "00111100",10659 => "11100000",10660 => "10111011",10661 => "10101010",10662 => "11110111",10663 => "10110000",10664 => "11011100",10665 => "11001101",10666 => "01010110",10667 => "00111110",10668 => "00110101",10669 => "10011011",10670 => "00000011",10671 => "01110011",10672 => "00101101",10673 => "01000001",10674 => "00001000",10675 => "11000111",10676 => "00110000",10677 => "10101100",10678 => "10011101",10679 => "00010000",10680 => "00010011",10681 => "00110111",10682 => "11001110",10683 => "10100000",10684 => "11101111",10685 => "11111101",10686 => "00100100",10687 => "01000010",10688 => "00111011",10689 => "10111011",10690 => "10001101",10691 => "01001001",10692 => "11101000",10693 => "00100100",10694 => "10000011",10695 => "10111010",10696 => "00010000",10697 => "00001110",10698 => "00101011",10699 => "11001100",10700 => "01001110",10701 => "10101011",10702 => "01111010",10703 => "10110101",10704 => "10111111",10705 => "01100100",10706 => "10010010",10707 => "01010010",10708 => "00001101",10709 => "11111000",10710 => "01100101",10711 => "10000010",10712 => "10101101",10713 => "01000100",10714 => "11111111",10715 => "11000100",10716 => "01010000",10717 => "10000001",10718 => "00000101",10719 => "00010111",10720 => "11000000",10721 => "01110110",10722 => "10000110",10723 => "01110111",10724 => "00100011",10725 => "10100100",10726 => "00101101",10727 => "10001011",10728 => "01101001",10729 => "01001011",10730 => "11011100",10731 => "11101110",10732 => "11001011",10733 => "01111011",10734 => "11000000",10735 => "10011111",10736 => "00000111",10737 => "00110010",10738 => "10000101",10739 => "11100001",10740 => "10010010",10741 => "11011011",10742 => "10000001",10743 => "11111011",10744 => "10101000",10745 => "11110000",10746 => "10110111",10747 => "10000011",10748 => "10001111",10749 => "10010010",10750 => "01001110",10751 => "11010011",10752 => "11000110",10753 => "10101000",10754 => "00001001",10755 => "00101101",10756 => "11011101",10757 => "10010111",10758 => "10110010",10759 => "11011000",10760 => "11001011",10761 => "10101100",10762 => "00100001",10763 => "10110111",10764 => "00000010",10765 => "01011101",10766 => "10011101",10767 => "00110001",10768 => "11010001",10769 => "01000011",10770 => "10101110",10771 => "00111111",10772 => "01001010",10773 => "11001001",10774 => "00001001",10775 => "01011111",10776 => "10001110",10777 => "11100110",10778 => "01101011",10779 => "00100010",10780 => "11011110",10781 => "00111101",10782 => "11100101",10783 => "10110101",10784 => "00011101",10785 => "10111101",10786 => "10110100",10787 => "01101010",10788 => "01010011",10789 => "11100000",10790 => "01010110",10791 => "00111011",10792 => "01001100",10793 => "11111100",10794 => "00001111",10795 => "00011111",10796 => "10101111",10797 => "10001010",10798 => "11111100",10799 => "11101110",10800 => "10100001",10801 => "11001000",10802 => "01100001",10803 => "00100101",10804 => "00101110",10805 => "01100110",10806 => "00001011",10807 => "10100001",10808 => "01001011",10809 => "11101011",10810 => "00000011",10811 => "00010100",10812 => "00111100",10813 => "00100011",10814 => "01111001",10815 => "00010100",10816 => "11111001",10817 => "01111101",10818 => "10011010",10819 => "11010000",10820 => "00111010",10821 => "00011011",10822 => "11011001",10823 => "01110100",10824 => "00101101",10825 => "00001001",10826 => "01110101",10827 => "00101111",10828 => "00011110",10829 => "11010110",10830 => "11001100",10831 => "10110000",10832 => "01111011",10833 => "11010000",10834 => "11100101",10835 => "01001111",10836 => "00111100",10837 => "00011111",10838 => "01100111",10839 => "01010110",10840 => "00010100",10841 => "11001001",10842 => "11011011",10843 => "01011110",10844 => "00000011",10845 => "10011100",10846 => "11110010",10847 => "10100011",10848 => "11100111",10849 => "00110100",10850 => "10001010",10851 => "01000110",10852 => "11000000",10853 => "00011101",10854 => "01100011",10855 => "10000001",10856 => "00101111",10857 => "00011001",10858 => "00100011",10859 => "10011001",10860 => "11110110",10861 => "10001001",10862 => "10100101",10863 => "10000000",10864 => "11001110",10865 => "11111010",10866 => "11011011",10867 => "11011100",10868 => "10110110",10869 => "01111010",10870 => "10000001",10871 => "10000100",10872 => "11001111",10873 => "01000011",10874 => "00101010",10875 => "10000011",10876 => "01100011",10877 => "10110110",10878 => "01111001",10879 => "00010001",10880 => "11000001",10881 => "00000110",10882 => "00110001",10883 => "00100000",10884 => "11000111",10885 => "01100011",10886 => "00011001",10887 => "01101000",10888 => "01001011",10889 => "10011111",10890 => "00000101",10891 => "10101100",10892 => "01100110",10893 => "01111111",10894 => "11000101",10895 => "10100001",10896 => "00001111",10897 => "01001111",10898 => "10001011",10899 => "00000111",10900 => "11100010",10901 => "00111111",10902 => "10101111",10903 => "11011101",10904 => "10100011",10905 => "01110101",10906 => "11000110",10907 => "01100111",10908 => "10011000",10909 => "00001000",10910 => "00101011",10911 => "00001010",10912 => "10111001",10913 => "01100101",10914 => "01101011",10915 => "00011111",10916 => "10011111",10917 => "10110100",10918 => "10000111",10919 => "11100111",10920 => "01110000",10921 => "11101000",10922 => "11110010",10923 => "00000001",10924 => "01010011",10925 => "01001101",10926 => "00101000",10927 => "10001101",10928 => "10000101",10929 => "00110010",10930 => "00101011",10931 => "00100110",10932 => "11110111",10933 => "10111011",10934 => "11000011",10935 => "00111111",10936 => "00011110",10937 => "10100011",10938 => "10001001",10939 => "00000101",10940 => "01111101",10941 => "00111111",10942 => "01001001",10943 => "01000111",10944 => "10101100",10945 => "01101111",10946 => "11001111",10947 => "01011110",10948 => "00000100",10949 => "10110110",10950 => "00100101",10951 => "01100111",10952 => "11000100",10953 => "11010111",10954 => "01101010",10955 => "11011000",10956 => "11000000",10957 => "00011000",10958 => "11111111",10959 => "00111110",10960 => "10101001",10961 => "11011110",10962 => "11001010",10963 => "10010011",10964 => "10101011",10965 => "10001000",10966 => "11010101",10967 => "00011000",10968 => "11100010",10969 => "10101000",10970 => "11110000",10971 => "00010111",10972 => "11111001",10973 => "01110100",10974 => "11011010",10975 => "01101000",10976 => "01100010",10977 => "01101001",10978 => "10101111",10979 => "10001011",10980 => "10100110",10981 => "01101011",10982 => "00011111",10983 => "01101110",10984 => "01100111",10985 => "11001001",10986 => "10110111",10987 => "10111111",10988 => "11100010",10989 => "01011110",10990 => "11011101",10991 => "10111001",10992 => "11110011",10993 => "01000110",10994 => "00011011",10995 => "10100111",10996 => "01001111",10997 => "00000101",10998 => "00101111",10999 => "00011111",11000 => "00111001",11001 => "11001001",11002 => "01111101",11003 => "11001010",11004 => "10011010",11005 => "11111100",11006 => "11011010",11007 => "00010001",11008 => "00011011",11009 => "11101101",11010 => "11100010",11011 => "11100000",11012 => "11001011",11013 => "00101111",11014 => "01100010",11015 => "10000010",11016 => "10111001",11017 => "01100111",11018 => "00101001",11019 => "10111011",11020 => "11110100",11021 => "11110101",11022 => "00110011",11023 => "01110010",11024 => "01111000",11025 => "01001010",11026 => "01000111",11027 => "00100010",11028 => "01100000",11029 => "11000010",11030 => "00001111",11031 => "10011011",11032 => "00011111",11033 => "01110010",11034 => "01101011",11035 => "11111111",11036 => "00011001",11037 => "10001010",11038 => "11100111",11039 => "01110000",11040 => "01010100",11041 => "11010100",11042 => "10000001",11043 => "11111000",11044 => "01110001",11045 => "11001011",11046 => "11011010",11047 => "00010100",11048 => "11101010",11049 => "00100001",11050 => "10111001",11051 => "00111111",11052 => "01001111",11053 => "00111100",11054 => "00100100",11055 => "00111011",11056 => "00001011",11057 => "01111100",11058 => "00111000",11059 => "00010011",11060 => "01010110",11061 => "00101011",11062 => "01110111",11063 => "10001101",11064 => "10000101",11065 => "00010111",11066 => "11000001",11067 => "11110001",11068 => "11100100",11069 => "00010111",11070 => "11110000",11071 => "11011011",11072 => "10111000",11073 => "00001100",11074 => "00101111",11075 => "11000011",11076 => "10110100",11077 => "11001010",11078 => "10010100",11079 => "11110101",11080 => "00000000",11081 => "01111001",11082 => "10010101",11083 => "00000100",11084 => "00100101",11085 => "01100101",11086 => "00010100",11087 => "11010101",11088 => "11101000",11089 => "11101010",11090 => "11100110",11091 => "11010000",11092 => "10011010",11093 => "00010110",11094 => "00111000",11095 => "10101011",11096 => "10001000",11097 => "00111010",11098 => "00011011",11099 => "01011000",11100 => "01001110",11101 => "10010110",11102 => "11010110",11103 => "11000110",11104 => "10010011",11105 => "00011001",11106 => "10010010",11107 => "10001010",11108 => "01010100",11109 => "10011010",11110 => "11000100",11111 => "11011110",11112 => "10000001",11113 => "10101100",11114 => "01111011",11115 => "00101110",11116 => "11111110",11117 => "00011111",11118 => "01010100",11119 => "01000101",11120 => "11101101",11121 => "01111110",11122 => "01111000",11123 => "10001101",11124 => "00110011",11125 => "00000010",11126 => "10111110",11127 => "10010110",11128 => "10011111",11129 => "10101101",11130 => "00111011",11131 => "01000101",11132 => "00000100",11133 => "01011101",11134 => "01111111",11135 => "10001010",11136 => "11011010",11137 => "11111100",11138 => "10101101",11139 => "01001001",11140 => "00111101",11141 => "11001011",11142 => "00101000",11143 => "01100001",11144 => "10110011",11145 => "11001001",11146 => "01100110",11147 => "11000010",11148 => "00101101",11149 => "01110101",11150 => "11101011",11151 => "01100001",11152 => "11010111",11153 => "01000011",11154 => "10111001",11155 => "11100110",11156 => "00000001",11157 => "10101111",11158 => "01110000",11159 => "01010000",11160 => "11001001",11161 => "01000010",11162 => "11010100",11163 => "01100010",11164 => "11010000",11165 => "10110100",11166 => "11000011",11167 => "11110110",11168 => "01111000",11169 => "00101110",11170 => "00010100",11171 => "11110111",11172 => "10101001",11173 => "01011111",11174 => "11010010",11175 => "01011110",11176 => "11110110",11177 => "01111000",11178 => "01011101",11179 => "10111011",11180 => "11000010",11181 => "10101111",11182 => "01000000",11183 => "10111101",11184 => "00001101",11185 => "01111000",11186 => "00010001",11187 => "00010100",11188 => "11001011",11189 => "00111111",11190 => "11111000",11191 => "11010101",11192 => "11010100",11193 => "10001110",11194 => "00010110",11195 => "01010110",11196 => "00110100",11197 => "00110001",11198 => "10010111",11199 => "00010101",11200 => "10010001",11201 => "10100011",11202 => "01111101",11203 => "10110001",11204 => "00000001",11205 => "00101100",11206 => "11000001",11207 => "00101110",11208 => "11001110",11209 => "00110010",11210 => "11110000",11211 => "10100111",11212 => "10010001",11213 => "00100001",11214 => "01000010",11215 => "10111110",11216 => "11101001",11217 => "00010011",11218 => "11110110",11219 => "00111000",11220 => "11010011",11221 => "10101010",11222 => "10111110",11223 => "01001100",11224 => "11011100",11225 => "01010001",11226 => "10011011",11227 => "11101101",11228 => "01010001",11229 => "11011001",11230 => "10100101",11231 => "11010001",11232 => "11111100",11233 => "11100110",11234 => "10011001",11235 => "00111010",11236 => "11111001",11237 => "00110001",11238 => "10001101",11239 => "10010001",11240 => "11110011",11241 => "01010100",11242 => "11101101",11243 => "00001001",11244 => "11111001",11245 => "00111000",11246 => "10011011",11247 => "11011100",11248 => "00011110",11249 => "10111100",11250 => "00010101",11251 => "10101100",11252 => "01000011",11253 => "00000011",11254 => "10010000",11255 => "10011101",11256 => "01010111",11257 => "00111010",11258 => "10111100",11259 => "00111100",11260 => "11000001",11261 => "01010111",11262 => "10010001",11263 => "11010110",11264 => "01101100",11265 => "01011110",11266 => "01100110",11267 => "11111101",11268 => "11001001",11269 => "11101110",11270 => "00000111",11271 => "01010111",11272 => "00010010",11273 => "01100101",11274 => "00010010",11275 => "10100100",11276 => "11100111",11277 => "10110100",11278 => "11010100",11279 => "00101011",11280 => "00000001",11281 => "00000011",11282 => "11001011",11283 => "00000110",11284 => "01100111",11285 => "01001001",11286 => "11000011",11287 => "01001010",11288 => "11100010",11289 => "11111010",11290 => "01000111",11291 => "10011011",11292 => "10110000",11293 => "10100001",11294 => "11101000",11295 => "11111010",11296 => "00101101",11297 => "01101101",11298 => "10000110",11299 => "10101101",11300 => "00111101",11301 => "10000110",11302 => "00000010",11303 => "11010011",11304 => "10010111",11305 => "01010010",11306 => "00001000",11307 => "00011011",11308 => "01000001",11309 => "11110100",11310 => "11001011",11311 => "10000100",11312 => "11111011",11313 => "00000111",11314 => "01111110",11315 => "11000010",11316 => "01010111",11317 => "10000110",11318 => "11100111",11319 => "11001110",11320 => "01101001",11321 => "10111100",11322 => "01100011",11323 => "01001100",11324 => "10010111",11325 => "00100001",11326 => "01111011",11327 => "00101101",11328 => "10111100",11329 => "00110100",11330 => "00000101",11331 => "00101000",11332 => "01101001",11333 => "00111011",11334 => "01100110",11335 => "00101001",11336 => "00010111",11337 => "01000111",11338 => "11011000",11339 => "00110010",11340 => "00100100",11341 => "11000111",11342 => "10100010",11343 => "01100111",11344 => "01111001",11345 => "10011100",11346 => "01011000",11347 => "11011010",11348 => "11111101",11349 => "01111100",11350 => "00100011",11351 => "00010001",11352 => "01101110",11353 => "01011000",11354 => "01001110",11355 => "11110010",11356 => "01011100",11357 => "01000110",11358 => "10011011",11359 => "01111000",11360 => "10101011",11361 => "00011101",11362 => "00000000",11363 => "00110011",11364 => "01100110",11365 => "11110100",11366 => "01010000",11367 => "01100010",11368 => "11000011",11369 => "11000011",11370 => "10011111",11371 => "00000000",11372 => "10011010",11373 => "00101010",11374 => "00001101",11375 => "10000101",11376 => "00110111",11377 => "00001101",11378 => "11001011",11379 => "11100101",11380 => "10001111",11381 => "10001000",11382 => "01011000",11383 => "10000101",11384 => "11111010",11385 => "10111110",11386 => "01000111",11387 => "00110001",11388 => "10011010",11389 => "00011001",11390 => "11110000",11391 => "00100010",11392 => "01110101",11393 => "00000001",11394 => "01111100",11395 => "01111111",11396 => "01010111",11397 => "00000001",11398 => "01110111",11399 => "01010011",11400 => "00010000",11401 => "00000001",11402 => "00101010",11403 => "01111111",11404 => "01100111",11405 => "00001011",11406 => "11010110",11407 => "10000111",11408 => "11001000",11409 => "10001101",11410 => "00011010",11411 => "01110001",11412 => "11111111",11413 => "00100000",11414 => "11010100",11415 => "11010011",11416 => "00101110",11417 => "01010000",11418 => "00100111",11419 => "01101100",11420 => "10001010",11421 => "00011111",11422 => "01001111",11423 => "11110101",11424 => "01110110",11425 => "00110000",11426 => "01110111",11427 => "00100001",11428 => "11011110",11429 => "10000100",11430 => "00011010",11431 => "01100101",11432 => "11000101",11433 => "11111110",11434 => "00000000",11435 => "10010101",11436 => "10011100",11437 => "10001001",11438 => "01001111",11439 => "00000100",11440 => "00100001",11441 => "00101110",11442 => "10100000",11443 => "01110110",11444 => "10001001",11445 => "00011010",11446 => "11100100",11447 => "00100001",11448 => "01011110",11449 => "00110010",11450 => "10001000",11451 => "00111100",11452 => "10101011",11453 => "10011001",11454 => "00010101",11455 => "01011000",11456 => "01110010",11457 => "01111001",11458 => "10101100",11459 => "11001011",11460 => "01011100",11461 => "01110100",11462 => "00100100",11463 => "10010111",11464 => "10011111",11465 => "10000111",11466 => "00001010",11467 => "11010010",11468 => "10100011",11469 => "11000111",11470 => "11111101",11471 => "01000010",11472 => "11010010",11473 => "11011101",11474 => "01100001",11475 => "01010111",11476 => "11001111",11477 => "00111101",11478 => "01011110",11479 => "01011010",11480 => "11110000",11481 => "01011000",11482 => "10101100",11483 => "00001111",11484 => "01111111",11485 => "10010011",11486 => "01111101",11487 => "01101101",11488 => "11110011",11489 => "00010101",11490 => "01010111",11491 => "01101001",11492 => "00100000",11493 => "10100110",11494 => "00010100",11495 => "00011011",11496 => "01000000",11497 => "10000110",11498 => "00110111",11499 => "10001011",11500 => "01110100",11501 => "00100101",11502 => "10110010",11503 => "00110100",11504 => "10011000",11505 => "10001100",11506 => "01111111",11507 => "10011010",11508 => "00010010",11509 => "00001100",11510 => "00001111",11511 => "01110111",11512 => "10101100",11513 => "00100001",11514 => "10001111",11515 => "10001110",11516 => "11010001",11517 => "01111001",11518 => "01010110",11519 => "10101111",11520 => "10011001",11521 => "11110011",11522 => "00001001",11523 => "01001010",11524 => "10100110",11525 => "10100000",11526 => "11010001",11527 => "01110011",11528 => "10101111",11529 => "11100111",11530 => "01010011",11531 => "11010100",11532 => "11011110",11533 => "10001001",11534 => "11011010",11535 => "01111100",11536 => "11100000",11537 => "11101001",11538 => "00100111",11539 => "11111011",11540 => "11001010",11541 => "00011101",11542 => "10001000",11543 => "00111011",11544 => "10100000",11545 => "11111010",11546 => "10101010",11547 => "11101000",11548 => "00001000",11549 => "01111011",11550 => "11110100",11551 => "01000001",11552 => "11011001",11553 => "10001111",11554 => "00001111",11555 => "00000101",11556 => "01000111",11557 => "10010001",11558 => "11110100",11559 => "11101100",11560 => "11100110",11561 => "00011100",11562 => "00100110",11563 => "10000010",11564 => "11010001",11565 => "01001010",11566 => "00110110",11567 => "01100100",11568 => "01110100",11569 => "10000100",11570 => "01100010",11571 => "10000011",11572 => "00110110",11573 => "01001101",11574 => "00001011",11575 => "00000101",11576 => "01011111",11577 => "11000100",11578 => "10000100",11579 => "11001010",11580 => "00010101",11581 => "10110001",11582 => "11000110",11583 => "10111110",11584 => "11011010",11585 => "00001111",11586 => "01111011",11587 => "01001001",11588 => "00101110",11589 => "11111111",11590 => "11101000",11591 => "01010110",11592 => "01010111",11593 => "00100011",11594 => "10101001",11595 => "01100011",11596 => "00010001",11597 => "01110110",11598 => "10111011",11599 => "10011000",11600 => "00000110",11601 => "00100011",11602 => "01000011",11603 => "00101001",11604 => "00110010",11605 => "01101010",11606 => "01011101",11607 => "11111100",11608 => "01100000",11609 => "00110001",11610 => "10100011",11611 => "01011110",11612 => "11110011",11613 => "00110001",11614 => "11111010",11615 => "00011100",11616 => "01110000",11617 => "10111001",11618 => "01000111",11619 => "10011000",11620 => "11010010",11621 => "10101111",11622 => "00001110",11623 => "00110011",11624 => "00010011",11625 => "10100011",11626 => "01110100",11627 => "01010101",11628 => "01000110",11629 => "10011110",11630 => "01100011",11631 => "01000100",11632 => "11001000",11633 => "10110001",11634 => "10110001",11635 => "11101010",11636 => "10011111",11637 => "10110000",11638 => "01100110",11639 => "11100101",11640 => "00100100",11641 => "10011100",11642 => "00010010",11643 => "00001010",11644 => "11010100",11645 => "10011111",11646 => "10000110",11647 => "10010011",11648 => "11011101",11649 => "10001100",11650 => "10100111",11651 => "00110001",11652 => "11000010",11653 => "00010001",11654 => "01101100",11655 => "11000100",11656 => "00011100",11657 => "01010001",11658 => "00011101",11659 => "10100100",11660 => "00000001",11661 => "10000100",11662 => "10111000",11663 => "00100111",11664 => "00011101",11665 => "10111000",11666 => "10110011",11667 => "10110101",11668 => "10010100",11669 => "01010010",11670 => "01011011",11671 => "00011010",11672 => "00110110",11673 => "01010100",11674 => "00110000",11675 => "10010010",11676 => "00110110",11677 => "00111010",11678 => "10110000",11679 => "01110001",11680 => "11100101",11681 => "00100111",11682 => "01100010",11683 => "01000010",11684 => "00010000",11685 => "10110000",11686 => "10001101",11687 => "00111010",11688 => "00001011",11689 => "10101111",11690 => "11000010",11691 => "01011010",11692 => "11010010",11693 => "10101100",11694 => "00000100",11695 => "01101101",11696 => "01001001",11697 => "10101111",11698 => "01111101",11699 => "10001001",11700 => "11101110",11701 => "10010001",11702 => "00000110",11703 => "00010100",11704 => "10010111",11705 => "11101010",11706 => "10001110",11707 => "00011111",11708 => "11111011",11709 => "11010110",11710 => "01011110",11711 => "10110010",11712 => "11000001",11713 => "10000000",11714 => "00011110",11715 => "11001001",11716 => "10010000",11717 => "00001110",11718 => "00011100",11719 => "11110110",11720 => "10011111",11721 => "11100111",11722 => "11011011",11723 => "01100100",11724 => "00011101",11725 => "11000111",11726 => "11100000",11727 => "11100001",11728 => "01101100",11729 => "11111111",11730 => "00100111",11731 => "10110111",11732 => "01101111",11733 => "00101110",11734 => "01011111",11735 => "00010100",11736 => "00010111",11737 => "10010001",11738 => "11010101",11739 => "00110000",11740 => "00101011",11741 => "11101100",11742 => "00110101",11743 => "10001010",11744 => "10100000",11745 => "10010001",11746 => "00001000",11747 => "00001100",11748 => "00100101",11749 => "01100000",11750 => "00011111",11751 => "11111001",11752 => "10010111",11753 => "11010110",11754 => "11100011",11755 => "00101011",11756 => "00111010",11757 => "00101011",11758 => "11011100",11759 => "01110000",11760 => "00110001",11761 => "00101000",11762 => "01001001",11763 => "01011011",11764 => "00011111",11765 => "01011111",11766 => "10100100",11767 => "00100010",11768 => "01110011",11769 => "11101101",11770 => "01101010",11771 => "11011110",11772 => "10110110",11773 => "11000011",11774 => "01011011",11775 => "11101011",11776 => "11001100",11777 => "00101001",11778 => "10011101",11779 => "01010101",11780 => "11111101",11781 => "00010010",11782 => "01110110",11783 => "11011101",11784 => "01011110",11785 => "10010011",11786 => "11010101",11787 => "01011101",11788 => "10101110",11789 => "10001110",11790 => "01101001",11791 => "10111001",11792 => "00011110",11793 => "00111010",11794 => "00000001",11795 => "11001010",11796 => "01110000",11797 => "01010011",11798 => "10101010",11799 => "01011000",11800 => "01100011",11801 => "10101010",11802 => "11010101",11803 => "10010001",11804 => "01010000",11805 => "00111000",11806 => "01010001",11807 => "10000000",11808 => "01001011",11809 => "00011110",11810 => "00000101",11811 => "00111101",11812 => "11010110",11813 => "00110110",11814 => "01010100",11815 => "10101011",11816 => "10001011",11817 => "10001010",11818 => "11010010",11819 => "01100000",11820 => "10110010",11821 => "00000000",11822 => "01000001",11823 => "01001010",11824 => "10001100",11825 => "10010101",11826 => "10000100",11827 => "01101111",11828 => "00101000",11829 => "00101110",11830 => "10000100",11831 => "01011000",11832 => "01000000",11833 => "01000110",11834 => "00001100",11835 => "11100101",11836 => "10001010",11837 => "11111111",11838 => "11010100",11839 => "11110000",11840 => "00111010",11841 => "01111111",11842 => "01000100",11843 => "00010101",11844 => "00100111",11845 => "00011011",11846 => "01110010",11847 => "10101111",11848 => "00001111",11849 => "01101100",11850 => "10000101",11851 => "00000000",11852 => "11110010",11853 => "01010010",11854 => "01011111",11855 => "10000111",11856 => "11101010",11857 => "00010100",11858 => "10011011",11859 => "10100000",11860 => "11100100",11861 => "01101001",11862 => "00000101",11863 => "11000001",11864 => "01010100",11865 => "10100001",11866 => "00001110",11867 => "00001000",11868 => "01010011",11869 => "00010100",11870 => "10110100",11871 => "11101001",11872 => "00111110",11873 => "01101110",11874 => "10000000",11875 => "00110110",11876 => "01000011",11877 => "00101011",11878 => "00011010",11879 => "10001011",11880 => "10110001",11881 => "00100001",11882 => "11110000",11883 => "01001111",11884 => "11110100",11885 => "10101001",11886 => "01100111",11887 => "00101010",11888 => "00001111",11889 => "00011100",11890 => "10110010",11891 => "10000101",11892 => "11101001",11893 => "00111101",11894 => "10011110",11895 => "10011101",11896 => "11111001",11897 => "00001101",11898 => "11010000",11899 => "00111010",11900 => "01100001",11901 => "10101001",11902 => "11111111",11903 => "10000110",11904 => "11001001",11905 => "01011001",11906 => "00010011",11907 => "10110011",11908 => "11000000",11909 => "10111001",11910 => "00100101",11911 => "11111101",11912 => "01101010",11913 => "01001000",11914 => "11001000",11915 => "01100001",11916 => "00011010",11917 => "11111010",11918 => "11001011",11919 => "00100100",11920 => "11100000",11921 => "01010010",11922 => "00100111",11923 => "10011001",11924 => "01011001",11925 => "11010000",11926 => "10010000",11927 => "11111111",11928 => "11111111",11929 => "00011100",11930 => "11110000",11931 => "01101100",11932 => "01000101",11933 => "01100100",11934 => "11001011",11935 => "01011100",11936 => "00000110",11937 => "00100111",11938 => "01011111",11939 => "00010100",11940 => "01000110",11941 => "11010001",11942 => "11001100",11943 => "01001000",11944 => "00111011",11945 => "11010111",11946 => "11011101",11947 => "10110100",11948 => "00010000",11949 => "00101101",11950 => "00100110",11951 => "00001010",11952 => "11111100",11953 => "00111101",11954 => "11111100",11955 => "11100000",11956 => "11110000",11957 => "10101111",11958 => "11010010",11959 => "10011000",11960 => "11110001",11961 => "11011001",11962 => "10100001",11963 => "10001000",11964 => "00010011",11965 => "11111000",11966 => "01010100",11967 => "11110111",11968 => "01001010",11969 => "11011101",11970 => "00010111",11971 => "01110100",11972 => "00001100",11973 => "00000001",11974 => "10101111",11975 => "00110110",11976 => "11101101",11977 => "10001001",11978 => "01101110",11979 => "01100100",11980 => "11110101",11981 => "00101001",11982 => "11101010",11983 => "00011010",11984 => "10000000",11985 => "00001010",11986 => "10000010",11987 => "10111100",11988 => "11011111",11989 => "10111011",11990 => "00011000",11991 => "11000011",11992 => "11001001",11993 => "01001000",11994 => "11100101",11995 => "11101001",11996 => "10110100",11997 => "00110000",11998 => "00100110",11999 => "10011001",12000 => "10011100",12001 => "00110010",12002 => "10010001",12003 => "11011101",12004 => "10000001",12005 => "10100101",12006 => "10000110",12007 => "01001111",12008 => "01011001",12009 => "10100110",12010 => "01000101",12011 => "01010100",12012 => "00011100",12013 => "11100101",12014 => "10110010",12015 => "01101010",12016 => "00101110",12017 => "00100111",12018 => "10001010",12019 => "00101000",12020 => "10100110",12021 => "10110000",12022 => "10010010",12023 => "10001001",12024 => "11110000",12025 => "00011111",12026 => "01011101",12027 => "11000101",12028 => "01000000",12029 => "01011100",12030 => "01001111",12031 => "10000000",12032 => "10011100",12033 => "01101001",12034 => "00010011",12035 => "01000100",12036 => "00011101",12037 => "10100001",12038 => "11100101",12039 => "10010100",12040 => "01010001",12041 => "01111111",12042 => "00100001",12043 => "01111000",12044 => "11010100",12045 => "11100011",12046 => "11000010",12047 => "10111101",12048 => "10010110",12049 => "11110010",12050 => "10101000",12051 => "01000010",12052 => "01111110",12053 => "01111110",12054 => "01000110",12055 => "11011010",12056 => "01010010",12057 => "10100001",12058 => "10001100",12059 => "01100101",12060 => "11100011",12061 => "01100100",12062 => "00100011",12063 => "01000110",12064 => "01001110",12065 => "01100011",12066 => "00110000",12067 => "00111101",12068 => "10001100",12069 => "10001001",12070 => "01101011",12071 => "01000011",12072 => "10000001",12073 => "00110001",12074 => "01101100",12075 => "00110001",12076 => "01100000",12077 => "11011011",12078 => "10110010",12079 => "00011100",12080 => "11001110",12081 => "11101000",12082 => "10001101",12083 => "01100111",12084 => "01110001",12085 => "01101111",12086 => "11001111",12087 => "01101010",12088 => "01110101",12089 => "10011011",12090 => "01100111",12091 => "00001011",12092 => "10100101",12093 => "11000000",12094 => "00101001",12095 => "11000000",12096 => "10101011",12097 => "00000100",12098 => "10001100",12099 => "00101010",12100 => "11100111",12101 => "10100111",12102 => "00011110",12103 => "10110011",12104 => "01011001",12105 => "10010011",12106 => "00001011",12107 => "11001101",12108 => "10010100",12109 => "01001101",12110 => "10110100",12111 => "01011101",12112 => "10100101",12113 => "01101011",12114 => "01100110",12115 => "00001111",12116 => "00111010",12117 => "11101010",12118 => "10101011",12119 => "01000101",12120 => "01000000",12121 => "10000011",12122 => "10000010",12123 => "01101001",12124 => "01000011",12125 => "10010100",12126 => "10000010",12127 => "01110100",12128 => "01111111",12129 => "11100101",12130 => "01100000",12131 => "10101111",12132 => "01110000",12133 => "01100110",12134 => "11001101",12135 => "10110110",12136 => "11001111",12137 => "10110011",12138 => "01110100",12139 => "11011111",12140 => "01001110",12141 => "01000010",12142 => "01101000",12143 => "11101111",12144 => "01101010",12145 => "10100100",12146 => "11011011",12147 => "01111100",12148 => "01100001",12149 => "10100011",12150 => "00011111",12151 => "10001110",12152 => "00111010",12153 => "00011101",12154 => "10010100",12155 => "01010100",12156 => "11011101",12157 => "10110001",12158 => "10101101",12159 => "11100111",12160 => "00011110",12161 => "00010011",12162 => "01110010",12163 => "10110010",12164 => "00111011",12165 => "00001010",12166 => "00001111",12167 => "00011100",12168 => "11110001",12169 => "00111010",12170 => "00001011",12171 => "11101000",12172 => "10111100",12173 => "00011101",12174 => "10010100",12175 => "11001011",12176 => "11110111",12177 => "11001000",12178 => "10110111",12179 => "11000000",12180 => "11000010",12181 => "10011010",12182 => "01100101",12183 => "01010101",12184 => "11000010",12185 => "00001111",12186 => "00001100",12187 => "01001111",12188 => "11110110",12189 => "01000011",12190 => "10001110",12191 => "11101100",12192 => "00010000",12193 => "01101000",12194 => "00000100",12195 => "11000000",12196 => "11000111",12197 => "11010011",12198 => "11001011",12199 => "10001011",12200 => "01000111",12201 => "11011101",12202 => "00110011",12203 => "00001011",12204 => "01011100",12205 => "11101101",12206 => "01111111",12207 => "10001011",12208 => "01000110",12209 => "10101101",12210 => "10110001",12211 => "00010011",12212 => "00101110",12213 => "10011111",12214 => "01111000",12215 => "01011011",12216 => "01111011",12217 => "11001101",12218 => "11110100",12219 => "10101010",12220 => "11000100",12221 => "11101110",12222 => "11000101",12223 => "01011100",12224 => "10000101",12225 => "11111101",12226 => "01111010",12227 => "11101101",12228 => "00011001",12229 => "10110000",12230 => "01001010",12231 => "00101000",12232 => "01101011",12233 => "10010000",12234 => "11110000",12235 => "00110101",12236 => "11000111",12237 => "10110001",12238 => "00010100",12239 => "01100101",12240 => "11000010",12241 => "10110011",12242 => "11100100",12243 => "10100011",12244 => "01011101",12245 => "00010010",12246 => "11000101",12247 => "10100111",12248 => "10100010",12249 => "10111001",12250 => "01111110",12251 => "00010110",12252 => "10001000",12253 => "11000110",12254 => "11001111",12255 => "10001011",12256 => "01010000",12257 => "11110111",12258 => "00111111",12259 => "01000000",12260 => "11000000",12261 => "00000010",12262 => "01100100",12263 => "01011001",12264 => "01101001",12265 => "00011000",12266 => "11110100",12267 => "10110111",12268 => "10001010",12269 => "01100000",12270 => "01111010",12271 => "00010100",12272 => "10110111",12273 => "11000010",12274 => "11101110",12275 => "10001011",12276 => "11101100",12277 => "10000100",12278 => "01100001",12279 => "10001111",12280 => "01100100",12281 => "10111000",12282 => "00110000",12283 => "00111000",12284 => "00001011",12285 => "00001001",12286 => "11011011",12287 => "01100001",12288 => "00000101",12289 => "11100010",12290 => "01101101",12291 => "11010000",12292 => "01000100",12293 => "01111111",12294 => "10110010",12295 => "01111001",12296 => "00101111",12297 => "00001110",12298 => "00100000",12299 => "10011110",12300 => "01001001",12301 => "01010010",12302 => "11100111",12303 => "10000001",12304 => "00100011",12305 => "00000110",12306 => "10100011",12307 => "01111010",12308 => "10100100",12309 => "10001001",12310 => "00110111",12311 => "01000011",12312 => "11100000",12313 => "01010010",12314 => "10100011",12315 => "00101100",12316 => "10011001",12317 => "10000001",12318 => "11100101",12319 => "10001111",12320 => "00000100",12321 => "11000010",12322 => "10100110",12323 => "01110000",12324 => "11000010",12325 => "10000101",12326 => "10100010",12327 => "01000110",12328 => "00110010",12329 => "10111101",12330 => "10111101",12331 => "11010101",12332 => "11111011",12333 => "01100110",12334 => "10101100",12335 => "01111001",12336 => "11110101",12337 => "00011111",12338 => "00010100",12339 => "10010010",12340 => "00001001",12341 => "10111000",12342 => "10101011",12343 => "11000111",12344 => "11111000",12345 => "00101000",12346 => "01010100",12347 => "11001101",12348 => "00100111",12349 => "11001100",12350 => "01111110",12351 => "00101001",12352 => "00100110",12353 => "00111100",12354 => "10100111",12355 => "00100010",12356 => "10010010",12357 => "00010111",12358 => "01100101",12359 => "10001010",12360 => "01101011",12361 => "01100011",12362 => "10111110",12363 => "10100011",12364 => "01011000",12365 => "11101110",12366 => "01000101",12367 => "00100000",12368 => "01111101",12369 => "11010011",12370 => "00100100",12371 => "01001110",12372 => "00010011",12373 => "00000010",12374 => "10111111",12375 => "11100001",12376 => "10010011",12377 => "11111000",12378 => "10110101",12379 => "00010000",12380 => "10101110",12381 => "01101011",12382 => "01000001",12383 => "10000110",12384 => "00110010",12385 => "10000000",12386 => "10000110",12387 => "10101000",12388 => "11011011",12389 => "00000100",12390 => "11011001",12391 => "11010011",12392 => "10101010",12393 => "01110100",12394 => "00110100",12395 => "11001001",12396 => "01111111",12397 => "11100001",12398 => "01101000",12399 => "00010101",12400 => "01000010",12401 => "10011011",12402 => "10100100",12403 => "01010100",12404 => "10101101",12405 => "00001000",12406 => "11011001",12407 => "00110001",12408 => "01101100",12409 => "01010101",12410 => "00110000",12411 => "10100000",12412 => "10000111",12413 => "10011011",12414 => "00100000",12415 => "10000010",12416 => "10011100",12417 => "11000001",12418 => "01100111",12419 => "11001111",12420 => "01101011",12421 => "01100011",12422 => "00000001",12423 => "01011001",12424 => "00101110",12425 => "00110010",12426 => "10010100",12427 => "11101010",12428 => "01010010",12429 => "11001100",12430 => "01010100",12431 => "01011010",12432 => "11100000",12433 => "00000111",12434 => "00100001",12435 => "00010010",12436 => "01110110",12437 => "10011000",12438 => "01010100",12439 => "11111011",12440 => "11111100",12441 => "01101110",12442 => "10010000",12443 => "01101101",12444 => "01010111",12445 => "01001110",12446 => "00100100",12447 => "00101011",12448 => "00001100",12449 => "00010111",12450 => "00001010",12451 => "11010010",12452 => "00001101",12453 => "00010010",12454 => "11110110",12455 => "10101000",12456 => "00100110",12457 => "11011110",12458 => "01100101",12459 => "10000100",12460 => "01110011",12461 => "11100111",12462 => "00000111",12463 => "11011110",12464 => "11101000",12465 => "01110011",12466 => "10000001",12467 => "01010000",12468 => "11011100",12469 => "10110101",12470 => "01010010",12471 => "11101100",12472 => "01011000",12473 => "11010011",12474 => "11011011",12475 => "01000010",12476 => "11101111",12477 => "10000101",12478 => "10100100",12479 => "01000001",12480 => "00111111",12481 => "00011010",12482 => "01101101",12483 => "10010000",12484 => "11010110",12485 => "10000111",12486 => "01101111",12487 => "10101000",12488 => "10100000",12489 => "10011101",12490 => "01101010",12491 => "10111101",12492 => "10110111",12493 => "10001000",12494 => "01101000",12495 => "10110011",12496 => "00100000",12497 => "10000011",12498 => "11100110",12499 => "10111010",12500 => "01100111",12501 => "00000110",12502 => "00110011",12503 => "10100011",12504 => "01110001",12505 => "01100100",12506 => "11110000",12507 => "10010100",12508 => "00100100",12509 => "00011101",12510 => "00100010",12511 => "10100101",12512 => "10101011",12513 => "11001001",12514 => "11100100",12515 => "11001111",12516 => "11010011",12517 => "11010011",12518 => "11101011",12519 => "01010111",12520 => "00000011",12521 => "00001011",12522 => "00010111",12523 => "10001100",12524 => "01100110",12525 => "01111100",12526 => "00110110",12527 => "10010011",12528 => "00100010",12529 => "11001000",12530 => "10110010",12531 => "10010000",12532 => "11000011",12533 => "00010111",12534 => "01010010",12535 => "11101001",12536 => "11100001",12537 => "11011111",12538 => "00101010",12539 => "01100100",12540 => "00111000",12541 => "00111100",12542 => "00000000",12543 => "01010101",12544 => "11100111",12545 => "11110000",12546 => "01111100",12547 => "01001010",12548 => "01000010",12549 => "00011000",12550 => "10110011",12551 => "11001111",12552 => "10000100",12553 => "10111101",12554 => "01000101",12555 => "00000000",12556 => "00111111",12557 => "01010011",12558 => "01101001",12559 => "00100101",12560 => "00001111",12561 => "00110100",12562 => "11010100",12563 => "00011000",12564 => "10011111",12565 => "11000101",12566 => "01001100",12567 => "11100100",12568 => "11001101",12569 => "11010001",12570 => "00011010",12571 => "10111111",12572 => "00010100",12573 => "11111010",12574 => "00101011",12575 => "11101100",12576 => "11001100",12577 => "01111111",12578 => "01110010",12579 => "00000010",12580 => "10011110",12581 => "00110110",12582 => "10111110",12583 => "00011010",12584 => "11001110",12585 => "11010000",12586 => "10011010",12587 => "00001001",12588 => "01011101",12589 => "01110111",12590 => "01101010",12591 => "00110101",12592 => "10110100",12593 => "10101010",12594 => "00111010",12595 => "01111001",12596 => "11101111",12597 => "00111010",12598 => "10111001",12599 => "01000100",12600 => "01010001",12601 => "11110111",12602 => "01011100",12603 => "00001001",12604 => "10010000",12605 => "10111111",12606 => "11110000",12607 => "01100010",12608 => "11011100",12609 => "01100110",12610 => "01101000",12611 => "01000111",12612 => "10000110",12613 => "00110111",12614 => "01110000",12615 => "11111100",12616 => "01011010",12617 => "10000100",12618 => "11111101",12619 => "00001111",12620 => "10001100",12621 => "10011101",12622 => "00011000",12623 => "10100111",12624 => "01000111",12625 => "00010101",12626 => "00111000",12627 => "01100001",12628 => "10101000",12629 => "11111011",12630 => "10110010",12631 => "10000000",12632 => "00100010",12633 => "11010011",12634 => "01001101",12635 => "00111101",12636 => "01110011",12637 => "01001110",12638 => "00111000",12639 => "11100111",12640 => "00110100",12641 => "11101111",12642 => "10101110",12643 => "01010001",12644 => "00010100",12645 => "00110110",12646 => "00001100",12647 => "10101101",12648 => "00111011",12649 => "00110011",12650 => "10110101",12651 => "11100010",12652 => "10110101",12653 => "10010111",12654 => "01100000",12655 => "10000100",12656 => "00001100",12657 => "00111010",12658 => "11110010",12659 => "00001101",12660 => "00011010",12661 => "00110011",12662 => "01011011",12663 => "00001100",12664 => "10101001",12665 => "10101100",12666 => "01000111",12667 => "00001100",12668 => "01010100",12669 => "01111010",12670 => "00011000",12671 => "10000101",12672 => "11111111",12673 => "10010111",12674 => "00011001",12675 => "01110010",12676 => "10101101",12677 => "00100000",12678 => "00011101",12679 => "01100101",12680 => "00001010",12681 => "10000110",12682 => "11110010",12683 => "00100011",12684 => "00010011",12685 => "11000010",12686 => "01011111",12687 => "00101100",12688 => "00001101",12689 => "10110100",12690 => "10100000",12691 => "00101011",12692 => "11111101",12693 => "00111010",12694 => "01010110",12695 => "01101001",12696 => "00000010",12697 => "11011101",12698 => "00110101",12699 => "11101000",12700 => "10110001",12701 => "10000101",12702 => "11000001",12703 => "11010001",12704 => "00100011",12705 => "01010111",12706 => "11001011",12707 => "10010101",12708 => "10111011",12709 => "10101110",12710 => "00101111",12711 => "01111101",12712 => "10100011",12713 => "01011111",12714 => "11101110",12715 => "10110111",12716 => "10111011",12717 => "00001010",12718 => "10111111",12719 => "01010101",12720 => "10110010",12721 => "11101110",12722 => "11111000",12723 => "01000001",12724 => "11011001",12725 => "01100101",12726 => "00101010",12727 => "01111001",12728 => "10101001",12729 => "11010100",12730 => "11011000",12731 => "00011101",12732 => "11101111",12733 => "01011100",12734 => "11101111",12735 => "10100010",12736 => "11110101",12737 => "10101111",12738 => "01001011",12739 => "10111111",12740 => "01111110",12741 => "11001000",12742 => "10010100",12743 => "01010011",12744 => "00111101",12745 => "10110001",12746 => "00101001",12747 => "01100000",12748 => "11111110",12749 => "00111010",12750 => "11000000",12751 => "10100111",12752 => "10001100",12753 => "10111000",12754 => "10100000",12755 => "00101100",12756 => "00101000",12757 => "00001010",12758 => "00000010",12759 => "00010111",12760 => "10110010",12761 => "10100100",12762 => "00100000",12763 => "10101100",12764 => "11101100",12765 => "00101000",12766 => "01100001",12767 => "01001010",12768 => "01111111",12769 => "10101011",12770 => "00010001",12771 => "01100100",12772 => "11011000",12773 => "11101110",12774 => "01111100",12775 => "11001110",12776 => "11001100",12777 => "00110010",12778 => "00111011",12779 => "00100010",12780 => "11011111",12781 => "10011001",12782 => "11011001",12783 => "10000101",12784 => "10001011",12785 => "01110111",12786 => "00110111",12787 => "01101001",12788 => "10000011",12789 => "10011100",12790 => "00101011",12791 => "01101111",12792 => "11000011",12793 => "10100111",12794 => "11010010",12795 => "00111101",12796 => "01111100",12797 => "11111110",12798 => "11000111",12799 => "10010110",12800 => "01010010",12801 => "00101111",12802 => "10110100",12803 => "10010101",12804 => "00000001",12805 => "10101011",12806 => "00000001",12807 => "01110111",12808 => "11011100",12809 => "10101100",12810 => "11100111",12811 => "11011101",12812 => "01110001",12813 => "11001011",12814 => "01111000",12815 => "10111001",12816 => "10101010",12817 => "00100100",12818 => "01101010",12819 => "01100110",12820 => "10010110",12821 => "10101111",12822 => "01110111",12823 => "00011101",12824 => "01111000",12825 => "10101011",12826 => "00000101",12827 => "10000110",12828 => "11011000",12829 => "10100101",12830 => "11011011",12831 => "01110011",12832 => "10010000",12833 => "00100010",12834 => "10000010",12835 => "11111000",12836 => "11001000",12837 => "01011000",12838 => "00000111",12839 => "11010100",12840 => "10000011",12841 => "10001001",12842 => "11110111",12843 => "01000100",12844 => "00010100",12845 => "00011010",12846 => "00110000",12847 => "00011000",12848 => "10110010",12849 => "01111100",12850 => "11100111",12851 => "11101011",12852 => "00010100",12853 => "11110000",12854 => "11111100",12855 => "11111111",12856 => "11001010",12857 => "01001110",12858 => "00110110",12859 => "10010011",12860 => "11101100",12861 => "01001101",12862 => "01010010",12863 => "10011011",12864 => "00000110",12865 => "00111010",12866 => "00111110",12867 => "11111000",12868 => "10011111",12869 => "01100101",12870 => "01000010",12871 => "10110100",12872 => "10111110",12873 => "00011100",12874 => "11011010",12875 => "11110110",12876 => "10001101",12877 => "01010111",12878 => "11011001",12879 => "01001010",12880 => "00000110",12881 => "01001011",12882 => "00000011",12883 => "00110110",12884 => "01110111",12885 => "10010000",12886 => "01001001",12887 => "11011111",12888 => "11100100",12889 => "00011000",12890 => "10000100",12891 => "00100100",12892 => "11011000",12893 => "00011110",12894 => "10000110",12895 => "01000110",12896 => "00001011",12897 => "00111110",12898 => "00000110",12899 => "01010001",12900 => "01100110",12901 => "01111111",12902 => "00001010",12903 => "10100001",12904 => "11110010",12905 => "11111001",12906 => "00101100",12907 => "11000010",12908 => "00111100",12909 => "10010001",12910 => "10000101",12911 => "00011001",12912 => "11000000",12913 => "01010001",12914 => "01000110",12915 => "10011011",12916 => "00010011",12917 => "10100101",12918 => "10001111",12919 => "11100100",12920 => "10000110",12921 => "11010110",12922 => "10000100",12923 => "01000000",12924 => "11010100",12925 => "01101010",12926 => "10111101",12927 => "11111010",12928 => "11011001",12929 => "11100010",12930 => "11100111",12931 => "01100101",12932 => "10010101",12933 => "00101011",12934 => "01011110",12935 => "00001100",12936 => "00000010",12937 => "01011001",12938 => "00011100",12939 => "00010100",12940 => "11000110",12941 => "01010101",12942 => "00110000",12943 => "00100111",12944 => "10111000",12945 => "00001011",12946 => "01010110",12947 => "01000101",12948 => "01101001",12949 => "10110111",12950 => "11011011",12951 => "11101010",12952 => "01000100",12953 => "11100011",12954 => "10110011",12955 => "11100011",12956 => "00110001",12957 => "11010110",12958 => "00001111",12959 => "11100011",12960 => "00110111",12961 => "11011011",12962 => "00000111",12963 => "11011100",12964 => "11100100",12965 => "01001011",12966 => "00001101",12967 => "00001000",12968 => "10110100",12969 => "11001001",12970 => "00001110",12971 => "00100110",12972 => "01110011",12973 => "01110100",12974 => "01110111",12975 => "10100010",12976 => "11101010",12977 => "01101010",12978 => "00010111",12979 => "10010100",12980 => "01100001",12981 => "01010111",12982 => "10010010",12983 => "00011101",12984 => "01001110",12985 => "11000100",12986 => "10101111",12987 => "11011010",12988 => "10000011",12989 => "00010010",12990 => "11111100",12991 => "10011011",12992 => "11100000",12993 => "10111101",12994 => "01011001",12995 => "01010110",12996 => "11011101",12997 => "10011100",12998 => "11101000",12999 => "00011011",13000 => "01101101",13001 => "11101001",13002 => "11001011",13003 => "01001100",13004 => "00011110",13005 => "01110011",13006 => "10010000",13007 => "11001000",13008 => "01100110",13009 => "10111001",13010 => "11001001",13011 => "10001010",13012 => "10100000",13013 => "00001101",13014 => "10010101",13015 => "01101100",13016 => "00000111",13017 => "00111000",13018 => "00000010",13019 => "11000011",13020 => "01101010",13021 => "10101110",13022 => "11000110",13023 => "10100110",13024 => "00010011",13025 => "11100111",13026 => "00101011",13027 => "10000101",13028 => "10100000",13029 => "11010011",13030 => "01001100",13031 => "00011101",13032 => "10000100",13033 => "01010101",13034 => "11101011",13035 => "01010011",13036 => "01101111",13037 => "00001110",13038 => "00011101",13039 => "10111010",13040 => "00000110",13041 => "10010110",13042 => "11100110",13043 => "11010001",13044 => "11011010",13045 => "11111000",13046 => "01001101",13047 => "00100010",13048 => "11101111",13049 => "00011110",13050 => "00111001",13051 => "11011110",13052 => "10001111",13053 => "00000111",13054 => "01001000",13055 => "10110101",13056 => "10010010",13057 => "01011000",13058 => "01110001",13059 => "01110101",13060 => "00100100",13061 => "11110110",13062 => "01010001",13063 => "11010100",13064 => "10111010",13065 => "10111110",13066 => "00110010",13067 => "00111100",13068 => "00011000",13069 => "10001111",13070 => "11111101",13071 => "11011011",13072 => "11100101",13073 => "00011010",13074 => "01010010",13075 => "01011011",13076 => "01101010",13077 => "10111011",13078 => "00101101",13079 => "00111100",13080 => "11111001",13081 => "00110001",13082 => "10000100",13083 => "00110011",13084 => "11001101",13085 => "00100101",13086 => "11000001",13087 => "10110101",13088 => "01101011",13089 => "11010000",13090 => "11010001",13091 => "00111101",13092 => "11100101",13093 => "01110101",13094 => "10010000",13095 => "01110101",13096 => "00000111",13097 => "10011010",13098 => "01111110",13099 => "01010001",13100 => "10100000",13101 => "11001110",13102 => "00100001",13103 => "10100010",13104 => "10011011",13105 => "00100110",13106 => "11001100",13107 => "00101110",13108 => "11001011",13109 => "01011100",13110 => "01010101",13111 => "10101100",13112 => "00000101",13113 => "10111000",13114 => "01110101",13115 => "10110001",13116 => "01100001",13117 => "11110101",13118 => "11101000",13119 => "10101000",13120 => "10111100",13121 => "11110100",13122 => "01000110",13123 => "00110101",13124 => "00001110",13125 => "01100000",13126 => "01110100",13127 => "10001000",13128 => "10110111",13129 => "01111110",13130 => "00011101",13131 => "01001000",13132 => "01110101",13133 => "11111010",13134 => "10101001",13135 => "00010111",13136 => "00101001",13137 => "01111111",13138 => "11000100",13139 => "11001101",13140 => "10111011",13141 => "11101100",13142 => "11001000",13143 => "01111101",13144 => "01000110",13145 => "10101001",13146 => "00011100",13147 => "00111010",13148 => "10111000",13149 => "11111111",13150 => "00101110",13151 => "10010110",13152 => "10000000",13153 => "01111001",13154 => "11011001",13155 => "11000101",13156 => "10101010",13157 => "10001010",13158 => "11011000",13159 => "00100100",13160 => "10010110",13161 => "00000111",13162 => "11111011",13163 => "00100101",13164 => "10111100",13165 => "00000010",13166 => "01010111",13167 => "00001100",13168 => "01110000",13169 => "11110000",13170 => "00010010",13171 => "10110111",13172 => "11110010",13173 => "01111001",13174 => "10100111",13175 => "10001011",13176 => "10000110",13177 => "00110100",13178 => "10111011",13179 => "00001110",13180 => "01111000",13181 => "01000100",13182 => "01100011",13183 => "00100101",13184 => "11111001",13185 => "11101010",13186 => "11101011",13187 => "11100100",13188 => "10010010",13189 => "11000110",13190 => "01000000",13191 => "10100010",13192 => "01000011",13193 => "01100110",13194 => "11111101",13195 => "01001001",13196 => "11001100",13197 => "01101000",13198 => "11011010",13199 => "01001101",13200 => "10000110",13201 => "01110100",13202 => "10100111",13203 => "10011001",13204 => "00000001",13205 => "11100101",13206 => "11111001",13207 => "11111010",13208 => "01110001",13209 => "10101110",13210 => "10111011",13211 => "01100100",13212 => "00101010",13213 => "10110000",13214 => "10111010",13215 => "01101100",13216 => "01111101",13217 => "10010101",13218 => "10011111",13219 => "11001111",13220 => "11101001",13221 => "00111100",13222 => "11110110",13223 => "10100111",13224 => "10110111",13225 => "00000011",13226 => "00011110",13227 => "01000111",13228 => "11101000",13229 => "01111010",13230 => "11110111",13231 => "11100111",13232 => "11100110",13233 => "00001100",13234 => "11001011",13235 => "00010110",13236 => "01101110",13237 => "10001100",13238 => "11101011",13239 => "11010110",13240 => "11100001",13241 => "00110111",13242 => "11001101",13243 => "00001100",13244 => "10100111",13245 => "01100101",13246 => "11000010",13247 => "00100011",13248 => "10010011",13249 => "11101101",13250 => "11001101",13251 => "11111001",13252 => "00110110",13253 => "00111001",13254 => "00100101",13255 => "00111101",13256 => "11001001",13257 => "00010100",13258 => "10111100",13259 => "10000111",13260 => "01011010",13261 => "10010100",13262 => "01110110",13263 => "11100110",13264 => "10000011",13265 => "01100001",13266 => "01101011",13267 => "10101010",13268 => "10001100",13269 => "10001001",13270 => "00100111",13271 => "10101011",13272 => "11111000",13273 => "10110111",13274 => "10000110",13275 => "10110011",13276 => "11100000",13277 => "00111101",13278 => "11111110",13279 => "10011000",13280 => "10110000",13281 => "01100010",13282 => "11000001",13283 => "00100010",13284 => "11001011",13285 => "00010000",13286 => "10101101",13287 => "00010000",13288 => "00010110",13289 => "10001101",13290 => "01010100",13291 => "11010100",13292 => "11100111",13293 => "00110100",13294 => "01000101",13295 => "00110110",13296 => "11000000",13297 => "11110110",13298 => "01011010",13299 => "10010010",13300 => "00011101",13301 => "11001000",13302 => "01100011",13303 => "01001111",13304 => "01011010",13305 => "10101111",13306 => "01111110",13307 => "01001010",13308 => "00010100",13309 => "00000001",13310 => "01001011",13311 => "00110010",13312 => "00100011",13313 => "10001011",13314 => "11100000",13315 => "00101100",13316 => "01111011",13317 => "00111111",13318 => "01111111",13319 => "10001001",13320 => "00001001",13321 => "10010000",13322 => "11100011",13323 => "10110100",13324 => "10100000",13325 => "11111011",13326 => "11010110",13327 => "11000111",13328 => "11100010",13329 => "11111110",13330 => "00011111",13331 => "11111001",13332 => "10110000",13333 => "00110111",13334 => "01011010",13335 => "00111111",13336 => "11011110",13337 => "00000110",13338 => "10110010",13339 => "00100001",13340 => "01101010",13341 => "01011010",13342 => "01000010",13343 => "11011100",13344 => "01101011",13345 => "00010111",13346 => "10000011",13347 => "01011110",13348 => "11010010",13349 => "00000000",13350 => "11010101",13351 => "01011011",13352 => "00011010",13353 => "01010110",13354 => "00111100",13355 => "01011010",13356 => "11001001",13357 => "00101101",13358 => "11011100",13359 => "00011011",13360 => "10100111",13361 => "00111011",13362 => "01001010",13363 => "01110011",13364 => "00101010",13365 => "10001111",13366 => "00111110",13367 => "00110000",13368 => "01111011",13369 => "00100101",13370 => "10011101",13371 => "10101100",13372 => "10000111",13373 => "00110111",13374 => "01010110",13375 => "00010111",13376 => "00010100",13377 => "11010010",13378 => "01001100",13379 => "11110100",13380 => "00111101",13381 => "00001101",13382 => "10011111",13383 => "00001001",13384 => "01110000",13385 => "11010100",13386 => "10101101",13387 => "01011000",13388 => "11010111",13389 => "01010111",13390 => "00011010",13391 => "01000000",13392 => "00001101",13393 => "00111011",13394 => "01111010",13395 => "11010011",13396 => "00111001",13397 => "00001011",13398 => "01000101",13399 => "00101011",13400 => "01101110",13401 => "00110011",13402 => "01110111",13403 => "01110100",13404 => "00010011",13405 => "11100110",13406 => "01011000",13407 => "10110000",13408 => "11110010",13409 => "01001001",13410 => "11100010",13411 => "10100010",13412 => "10110001",13413 => "11000010",13414 => "10010000",13415 => "01010100",13416 => "11000100",13417 => "11001001",13418 => "01101111",13419 => "00001001",13420 => "00011011",13421 => "01011000",13422 => "01101111",13423 => "11101010",13424 => "10111100",13425 => "11000110",13426 => "10101111",13427 => "00011100",13428 => "11011001",13429 => "11110110",13430 => "10000000",13431 => "10011001",13432 => "01101011",13433 => "01010100",13434 => "10001010",13435 => "00001100",13436 => "01110010",13437 => "10111011",13438 => "10010011",13439 => "01111101",13440 => "10001001",13441 => "00100101",13442 => "11010011",13443 => "10010010",13444 => "11010100",13445 => "10101001",13446 => "00010011",13447 => "10110001",13448 => "10110010",13449 => "11011010",13450 => "10101100",13451 => "11011101",13452 => "00000001",13453 => "01010101",13454 => "10111001",13455 => "11111001",13456 => "01010001",13457 => "11101110",13458 => "10110110",13459 => "11110011",13460 => "10111010",13461 => "11011111",13462 => "11100011",13463 => "01011110",13464 => "00111001",13465 => "10100001",13466 => "00100010",13467 => "11110111",13468 => "11111101",13469 => "01101110",13470 => "01111111",13471 => "10000100",13472 => "00100000",13473 => "11111101",13474 => "11011111",13475 => "00100110",13476 => "10111100",13477 => "01010101",13478 => "00101100",13479 => "10010111",13480 => "10110001",13481 => "10001011",13482 => "10110001",13483 => "10101110",13484 => "11111011",13485 => "01110011",13486 => "00100000",13487 => "00100100",13488 => "00011011",13489 => "00001001",13490 => "00001110",13491 => "10111111",13492 => "00010011",13493 => "00000011",13494 => "10001100",13495 => "11001010",13496 => "10101100",13497 => "10011101",13498 => "01110110",13499 => "01000000",13500 => "01010101",13501 => "01011100",13502 => "10000010",13503 => "00111100",13504 => "11011101",13505 => "10100011",13506 => "01010111",13507 => "01011100",13508 => "10110000",13509 => "00011000",13510 => "11111000",13511 => "11110010",13512 => "11000010",13513 => "11111110",13514 => "01001101",13515 => "11111011",13516 => "10110001",13517 => "00001011",13518 => "00000101",13519 => "10110010",13520 => "10000101",13521 => "10000000",13522 => "01001000",13523 => "10011010",13524 => "01000100",13525 => "10100110",13526 => "10001111",13527 => "01100010",13528 => "11101000",13529 => "10101011",13530 => "01010000",13531 => "11101000",13532 => "00100111",13533 => "10111011",13534 => "01101100",13535 => "11111100",13536 => "11101110",13537 => "00010111",13538 => "10011001",13539 => "10101010",13540 => "00110010",13541 => "10110101",13542 => "00111101",13543 => "00011100",13544 => "00101010",13545 => "01000000",13546 => "01101110",13547 => "10011100",13548 => "00100001",13549 => "11001010",13550 => "01000111",13551 => "11001111",13552 => "11001000",13553 => "11000111",13554 => "11111110",13555 => "00011010",13556 => "00111101",13557 => "11101110",13558 => "10011010",13559 => "10010001",13560 => "01010101",13561 => "01000111",13562 => "01001011",13563 => "10000111",13564 => "00001101",13565 => "11010001",13566 => "10011000",13567 => "10011011",13568 => "11011101",13569 => "10111100",13570 => "01000001",13571 => "00110111",13572 => "10011010",13573 => "01001011",13574 => "01000101",13575 => "11001010",13576 => "00011010",13577 => "01101010",13578 => "01001011",13579 => "00011011",13580 => "10100111",13581 => "00001011",13582 => "10001110",13583 => "10010101",13584 => "10101000",13585 => "00001010",13586 => "10101100",13587 => "00001011",13588 => "10010101",13589 => "11001001",13590 => "10111101",13591 => "11001001",13592 => "11001000",13593 => "00111101",13594 => "11110000",13595 => "11110100",13596 => "01000011",13597 => "00001000",13598 => "10111010",13599 => "10001001",13600 => "01000101",13601 => "00010011",13602 => "11011111",13603 => "01001001",13604 => "00000010",13605 => "01001101",13606 => "00101100",13607 => "00011001",13608 => "01010101",13609 => "00011010",13610 => "00011110",13611 => "11101011",13612 => "00100001",13613 => "10100011",13614 => "10110011",13615 => "01110001",13616 => "01000001",13617 => "10101100",13618 => "11010100",13619 => "00011011",13620 => "11101010",13621 => "11111100",13622 => "00110111",13623 => "10001100",13624 => "01110111",13625 => "01001010",13626 => "11101010",13627 => "11001100",13628 => "01101101",13629 => "01000101",13630 => "00110011",13631 => "11100001",13632 => "00011000",13633 => "10001100",13634 => "10011011",13635 => "11101100",13636 => "10011111",13637 => "10110001",13638 => "11011110",13639 => "10110011",13640 => "10111110",13641 => "00100101",13642 => "00110000",13643 => "10011011",13644 => "10000001",13645 => "11011000",13646 => "11110110",13647 => "00100101",13648 => "01010101",13649 => "00101101",13650 => "00001000",13651 => "10110010",13652 => "00001100",13653 => "01000001",13654 => "10110111",13655 => "10100100",13656 => "10010101",13657 => "01001010",13658 => "00010001",13659 => "01000111",13660 => "10010111",13661 => "01110111",13662 => "00000110",13663 => "01100101",13664 => "00010001",13665 => "10100101",13666 => "01011001",13667 => "00000101",13668 => "00111111",13669 => "11101100",13670 => "10101101",13671 => "11000001",13672 => "00001011",13673 => "00011011",13674 => "00001101",13675 => "11111101",13676 => "10001101",13677 => "01101100",13678 => "11000010",13679 => "11001011",13680 => "00001001",13681 => "01101100",13682 => "11111001",13683 => "00101010",13684 => "10001000",13685 => "11110000",13686 => "10100001",13687 => "10000001",13688 => "01000101",13689 => "00101010",13690 => "01101010",13691 => "01011101",13692 => "10011111",13693 => "01101100",13694 => "00110011",13695 => "01101010",13696 => "01000000",13697 => "00101110",13698 => "01101111",13699 => "10110100",13700 => "10000110",13701 => "10101110",13702 => "00101011",13703 => "00100010",13704 => "01100111",13705 => "00001100",13706 => "11011110",13707 => "00010010",13708 => "11110110",13709 => "01110101",13710 => "11010111",13711 => "10001010",13712 => "01001101",13713 => "11001011",13714 => "10111001",13715 => "01010001",13716 => "11011001",13717 => "11000000",13718 => "00101011",13719 => "10011001",13720 => "01010111",13721 => "11001011",13722 => "01111000",13723 => "11101000",13724 => "11000100",13725 => "11110011",13726 => "11110100",13727 => "01101100",13728 => "10000011",13729 => "00110011",13730 => "11111011",13731 => "00101001",13732 => "00101010",13733 => "01010101",13734 => "01110100",13735 => "00000101",13736 => "00100100",13737 => "00001001",13738 => "11010011",13739 => "01001000",13740 => "10001010",13741 => "00000101",13742 => "01000000",13743 => "00111110",13744 => "10000001",13745 => "00011001",13746 => "10110011",13747 => "10111111",13748 => "00001110",13749 => "11101110",13750 => "01111000",13751 => "11001010",13752 => "11011111",13753 => "01011010",13754 => "10010010",13755 => "10111000",13756 => "00000111",13757 => "01110111",13758 => "00111100",13759 => "01110000",13760 => "10100110",13761 => "11000110",13762 => "10011111",13763 => "11011010",13764 => "11111111",13765 => "00111101",13766 => "00000011",13767 => "10000101",13768 => "11001011",13769 => "11000011",13770 => "11011110",13771 => "11000011",13772 => "01010010",13773 => "01000111",13774 => "10001011",13775 => "01110110",13776 => "10001000",13777 => "01000110",13778 => "11000011",13779 => "11010100",13780 => "01110001",13781 => "10011110",13782 => "00111010",13783 => "00111000",13784 => "11011110",13785 => "00000010",13786 => "11010101",13787 => "00101111",13788 => "00010011",13789 => "11101001",13790 => "11011011",13791 => "10000000",13792 => "11011010",13793 => "10000001",13794 => "01001101",13795 => "00001101",13796 => "10001110",13797 => "10110110",13798 => "00000101",13799 => "01110111",13800 => "00011110",13801 => "00010101",13802 => "10111010",13803 => "01011001",13804 => "00110000",13805 => "01010100",13806 => "01010100",13807 => "00101111",13808 => "01011011",13809 => "01110100",13810 => "10011001",13811 => "00010111",13812 => "00100011",13813 => "01110111",13814 => "00011010",13815 => "10011010",13816 => "01101010",13817 => "10011101",13818 => "10001110",13819 => "11111101",13820 => "00001011",13821 => "11011000",13822 => "10100000",13823 => "10110101",13824 => "11011010",13825 => "10000011",13826 => "10101000",13827 => "01100000",13828 => "10101100",13829 => "10110001",13830 => "00111001",13831 => "10011111",13832 => "11111101",13833 => "11110010",13834 => "11110011",13835 => "00011010",13836 => "00111111",13837 => "11111001",13838 => "10111100",13839 => "10100000",13840 => "10100011",13841 => "11101101",13842 => "11011110",13843 => "01010100",13844 => "01001001",13845 => "01010011",13846 => "00010101",13847 => "10100110",13848 => "00000100",13849 => "11111111",13850 => "00111101",13851 => "00100011",13852 => "10110110",13853 => "01001010",13854 => "01010011",13855 => "00011010",13856 => "10001101",13857 => "11111011",13858 => "10001110",13859 => "00100001",13860 => "11001101",13861 => "11110110",13862 => "00101101",13863 => "00011111",13864 => "11100111",13865 => "01111000",13866 => "10101101",13867 => "00000100",13868 => "10000011",13869 => "01101001",13870 => "11111000",13871 => "01010100",13872 => "01110001",13873 => "01101111",13874 => "11010110",13875 => "10101011",13876 => "11111000",13877 => "01011111",13878 => "01010001",13879 => "10100000",13880 => "00110011",13881 => "11111001",13882 => "11111100",13883 => "11101111",13884 => "10100101",13885 => "00101000",13886 => "00110001",13887 => "10001011",13888 => "10000101",13889 => "10100000",13890 => "00100010",13891 => "00011000",13892 => "00111111",13893 => "00110000",13894 => "01101001",13895 => "10000011",13896 => "01010100",13897 => "01100000",13898 => "00100000",13899 => "10101100",13900 => "11011011",13901 => "11101011",13902 => "11010101",13903 => "11001000",13904 => "00111111",13905 => "11001001",13906 => "00101111",13907 => "11011111",13908 => "00001011",13909 => "01011100",13910 => "00100010",13911 => "01100101",13912 => "01011110",13913 => "11101100",13914 => "10001000",13915 => "10111010",13916 => "01100000",13917 => "01111010",13918 => "10010011",13919 => "00110111",13920 => "10000110",13921 => "11111011",13922 => "10110011",13923 => "10011011",13924 => "10111010",13925 => "00100101",13926 => "11100011",13927 => "10101000",13928 => "00000001",13929 => "00100000",13930 => "00101111",13931 => "10011111",13932 => "00111011",13933 => "00110111",13934 => "10101101",13935 => "10100011",13936 => "00001101",13937 => "11110110",13938 => "00110001",13939 => "11000010",13940 => "11011100",13941 => "00001001",13942 => "00011101",13943 => "01001000",13944 => "11001011",13945 => "11000101",13946 => "11101000",13947 => "10001111",13948 => "10100001",13949 => "00111100",13950 => "00011110",13951 => "00000010",13952 => "10100010",13953 => "10111010",13954 => "10001000",13955 => "10010010",13956 => "00001111",13957 => "11110111",13958 => "11110100",13959 => "00011001",13960 => "11010101",13961 => "00011101",13962 => "00011100",13963 => "01001110",13964 => "11100000",13965 => "01101000",13966 => "10001010",13967 => "10001110",13968 => "00000001",13969 => "10010000",13970 => "11100101",13971 => "00101000",13972 => "00010111",13973 => "00001001",13974 => "00111111",13975 => "01101111",13976 => "11010011",13977 => "11111101",13978 => "10101011",13979 => "00100101",13980 => "00111110",13981 => "00001100",13982 => "11100110",13983 => "11001000",13984 => "10101000",13985 => "11100010",13986 => "10100001",13987 => "01100001",13988 => "11110110",13989 => "11010000",13990 => "01000110",13991 => "11100101",13992 => "00000100",13993 => "11110011",13994 => "11001000",13995 => "01011100",13996 => "00010011",13997 => "10110010",13998 => "01010100",13999 => "00111001",14000 => "00100111",14001 => "10101000",14002 => "01010010",14003 => "00110110",14004 => "11011111",14005 => "11001110",14006 => "00010111",14007 => "11010101",14008 => "10100101",14009 => "00001000",14010 => "00100011",14011 => "11000001",14012 => "10010000",14013 => "01111001",14014 => "00110010",14015 => "10000111",14016 => "01011100",14017 => "00100100",14018 => "00101011",14019 => "00111001",14020 => "10100101",14021 => "11010010",14022 => "01100101",14023 => "11110100",14024 => "10111010",14025 => "00100001",14026 => "00101001",14027 => "11000101",14028 => "01110110",14029 => "01001001",14030 => "11001110",14031 => "00111001",14032 => "10010100",14033 => "11111000",14034 => "01010001",14035 => "00001110",14036 => "11011111",14037 => "00001110",14038 => "01110111",14039 => "10101000",14040 => "00101001",14041 => "00010101",14042 => "00001101",14043 => "00100010",14044 => "11101010",14045 => "01110101",14046 => "11111010",14047 => "10000110",14048 => "01101010",14049 => "00110110",14050 => "10001011",14051 => "00001010",14052 => "01101101",14053 => "00010101",14054 => "10110011",14055 => "00011101",14056 => "11100100",14057 => "10010101",14058 => "10001001",14059 => "01011000",14060 => "11101110",14061 => "10000110",14062 => "10100010",14063 => "00101001",14064 => "10111111",14065 => "01101100",14066 => "01111111",14067 => "11101000",14068 => "11111111",14069 => "01110101",14070 => "11110100",14071 => "10100100",14072 => "01011100",14073 => "00110100",14074 => "01111111",14075 => "00000101",14076 => "00011110",14077 => "00110001",14078 => "10010110",14079 => "11100001",14080 => "11011011",14081 => "10001000",14082 => "01111000",14083 => "10110001",14084 => "11111001",14085 => "00010001",14086 => "00110001",14087 => "01100001",14088 => "11010010",14089 => "11011010",14090 => "10000101",14091 => "11100001",14092 => "00001101",14093 => "01010110",14094 => "01010001",14095 => "11100101",14096 => "10001110",14097 => "10011010",14098 => "11111000",14099 => "10110100",14100 => "00101011",14101 => "11111110",14102 => "11111000",14103 => "01110111",14104 => "10100110",14105 => "11000010",14106 => "00101011",14107 => "01111001",14108 => "00111110",14109 => "11000011",14110 => "11110010",14111 => "00101110",14112 => "00001110",14113 => "10000011",14114 => "10011010",14115 => "10101001",14116 => "01001110",14117 => "00100001",14118 => "01101101",14119 => "11000001",14120 => "10011111",14121 => "11111001",14122 => "10110111",14123 => "00101110",14124 => "01101001",14125 => "10001101",14126 => "10101111",14127 => "01001001",14128 => "11000110",14129 => "11000010",14130 => "01101010",14131 => "10111110",14132 => "11011111",14133 => "01101100",14134 => "00111110",14135 => "11011010",14136 => "01110010",14137 => "10011111",14138 => "10111011",14139 => "11101110",14140 => "11001100",14141 => "10011111",14142 => "00011000",14143 => "00000011",14144 => "10110100",14145 => "11001010",14146 => "00010011",14147 => "00101000",14148 => "01001100",14149 => "01101010",14150 => "11011010",14151 => "10000110",14152 => "10110011",14153 => "01010100",14154 => "00001101",14155 => "10010110",14156 => "10110111",14157 => "10010110",14158 => "01011000",14159 => "10111000",14160 => "00100111",14161 => "01111010",14162 => "00110101",14163 => "01011101",14164 => "01111101",14165 => "11100000",14166 => "00101000",14167 => "11100001",14168 => "11100111",14169 => "00011000",14170 => "01110110",14171 => "11111111",14172 => "10110101",14173 => "00110000",14174 => "01000000",14175 => "00001010",14176 => "01011001",14177 => "10101110",14178 => "10111000",14179 => "00000100",14180 => "10001100",14181 => "11100000",14182 => "00011010",14183 => "10111101",14184 => "10010101",14185 => "00101111",14186 => "11100010",14187 => "10100011",14188 => "11101101",14189 => "00110111",14190 => "11100111",14191 => "01110010",14192 => "00011110",14193 => "00100010",14194 => "11100001",14195 => "11011000",14196 => "10100010",14197 => "10010001",14198 => "00111000",14199 => "11101011",14200 => "00110101",14201 => "01101000",14202 => "10111110",14203 => "01110010",14204 => "00111100",14205 => "01010110",14206 => "00011001",14207 => "11101001",14208 => "10110000",14209 => "11010010",14210 => "00010000",14211 => "01101100",14212 => "01011111",14213 => "00101101",14214 => "01101001",14215 => "00100010",14216 => "10110011",14217 => "00111100",14218 => "01000110",14219 => "00010010",14220 => "11111011",14221 => "01110100",14222 => "11001110",14223 => "11100010",14224 => "11010110",14225 => "00000110",14226 => "01100011",14227 => "11000111",14228 => "01010101",14229 => "01100011",14230 => "00011001",14231 => "11101000",14232 => "00010111",14233 => "01111001",14234 => "00001000",14235 => "11111110",14236 => "10001111",14237 => "11001100",14238 => "11110010",14239 => "10111010",14240 => "10001111",14241 => "01001101",14242 => "11010001",14243 => "01001100",14244 => "10100101",14245 => "10000000",14246 => "01010001",14247 => "00110100",14248 => "11010011",14249 => "01010101",14250 => "10011001",14251 => "11011010",14252 => "11110101",14253 => "01111010",14254 => "11010001",14255 => "10000111",14256 => "01111000",14257 => "00011001",14258 => "01011111",14259 => "10110110",14260 => "11100111",14261 => "00011011",14262 => "00101001",14263 => "00101101",14264 => "10100100",14265 => "11000111",14266 => "10001110",14267 => "01010110",14268 => "00000010",14269 => "01000101",14270 => "11001110",14271 => "10101010",14272 => "00110110",14273 => "00011100",14274 => "11000011",14275 => "10110100",14276 => "01001001",14277 => "10011110",14278 => "00110110",14279 => "00111011",14280 => "10010111",14281 => "01000100",14282 => "11001011",14283 => "01000110",14284 => "11001000",14285 => "11111101",14286 => "00101000",14287 => "01001101",14288 => "01101011",14289 => "10010101",14290 => "11000100",14291 => "10100001",14292 => "00111010",14293 => "00111011",14294 => "10010111",14295 => "10100000",14296 => "10000001",14297 => "10000000",14298 => "00110101",14299 => "01100101",14300 => "10101100",14301 => "01000100",14302 => "01101101",14303 => "00001010",14304 => "11000100",14305 => "00001011",14306 => "10100100",14307 => "00111000",14308 => "11101011",14309 => "11101001",14310 => "10001110",14311 => "11100111",14312 => "11100111",14313 => "00110011",14314 => "10101010",14315 => "10111000",14316 => "10111101",14317 => "00011111",14318 => "00100011",14319 => "11100000",14320 => "10101110",14321 => "11100100",14322 => "11011010",14323 => "01011011",14324 => "00100001",14325 => "10011111",14326 => "11000111",14327 => "01111010",14328 => "11000101",14329 => "11011001",14330 => "11111111",14331 => "01101000",14332 => "11011101",14333 => "01111010",14334 => "00111111",14335 => "00110110",14336 => "00100000",14337 => "11010001",14338 => "00010001",14339 => "00000010",14340 => "11110110",14341 => "00110001",14342 => "01010001",14343 => "10001101",14344 => "11001111",14345 => "01101011",14346 => "01011111",14347 => "11101100",14348 => "10100010",14349 => "01110111",14350 => "01100101",14351 => "11100111",14352 => "01001011",14353 => "10100001",14354 => "01000001",14355 => "11110001",14356 => "00011110",14357 => "10010111",14358 => "10101101",14359 => "11110110",14360 => "00001001",14361 => "01100100",14362 => "00111101",14363 => "00101110",14364 => "11010110",14365 => "10101111",14366 => "01000010",14367 => "00000100",14368 => "00001101",14369 => "00101101",14370 => "10101001",14371 => "10101111",14372 => "01110000",14373 => "01001100",14374 => "11100001",14375 => "11001110",14376 => "11100111",14377 => "11000000",14378 => "00110101",14379 => "01100111",14380 => "11010111",14381 => "00000100",14382 => "00000100",14383 => "01111100",14384 => "10111000",14385 => "01100000",14386 => "00110001",14387 => "10101101",14388 => "10101011",14389 => "00010010",14390 => "11111010",14391 => "00000110",14392 => "11000001",14393 => "10110111",14394 => "00000001",14395 => "10110101",14396 => "01101110",14397 => "11101001",14398 => "01101001",14399 => "11001100",14400 => "01110000",14401 => "01010001",14402 => "10001001",14403 => "01110011",14404 => "11100110",14405 => "01101101",14406 => "11010001",14407 => "10010010",14408 => "01100010",14409 => "00001011",14410 => "11000001",14411 => "00110100",14412 => "01111001",14413 => "01101110",14414 => "00100111",14415 => "00101111",14416 => "00011011",14417 => "11111000",14418 => "11010011",14419 => "11110110",14420 => "00111100",14421 => "11011011",14422 => "01101001",14423 => "10011101",14424 => "00110110",14425 => "01101101",14426 => "11100101",14427 => "00000110",14428 => "00111000",14429 => "10110010",14430 => "00110001",14431 => "11110010",14432 => "10100001",14433 => "10111100",14434 => "01000101",14435 => "01001001",14436 => "10010001",14437 => "00000001",14438 => "01100011",14439 => "11001101",14440 => "00110111",14441 => "00110101",14442 => "00111000",14443 => "10111011",14444 => "10111001",14445 => "00101110",14446 => "10111011",14447 => "01100000",14448 => "10010011",14449 => "01101111",14450 => "00111110",14451 => "10010011",14452 => "11011100",14453 => "01100011",14454 => "10011010",14455 => "01010010",14456 => "00101101",14457 => "10101101",14458 => "11100111",14459 => "10011011",14460 => "00111001",14461 => "01000100",14462 => "01110101",14463 => "01001011",14464 => "11111111",14465 => "00100110",14466 => "00001111",14467 => "01011011",14468 => "11101001",14469 => "01111101",14470 => "00111100",14471 => "01101100",14472 => "01000010",14473 => "10001100",14474 => "10101001",14475 => "11101100",14476 => "11111010",14477 => "10100000",14478 => "01011101",14479 => "01111111",14480 => "10011101",14481 => "10000010",14482 => "00101010",14483 => "10110101",14484 => "11000001",14485 => "01101000",14486 => "11111100",14487 => "00010001",14488 => "01100001",14489 => "11111101",14490 => "10110011",14491 => "01010011",14492 => "01100011",14493 => "00100111",14494 => "11000101",14495 => "01110000",14496 => "00110101",14497 => "00101101",14498 => "10111101",14499 => "00110001",14500 => "10011101",14501 => "01100001",14502 => "00000000",14503 => "11101111",14504 => "00000101",14505 => "00000100",14506 => "10100110",14507 => "11001110",14508 => "10010010",14509 => "11010010",14510 => "10000011",14511 => "10101011",14512 => "01111001",14513 => "00110101",14514 => "10110111",14515 => "00110110",14516 => "10100111",14517 => "10011010",14518 => "00110010",14519 => "10101100",14520 => "01011111",14521 => "10000110",14522 => "01100101",14523 => "10110110",14524 => "10110011",14525 => "11100001",14526 => "01100000",14527 => "01100101",14528 => "11111110",14529 => "10000000",14530 => "01010010",14531 => "11101000",14532 => "10010101",14533 => "01100001",14534 => "11011011",14535 => "10110101",14536 => "00000010",14537 => "00010100",14538 => "01100100",14539 => "11100110",14540 => "01001011",14541 => "01101000",14542 => "11011101",14543 => "00011000",14544 => "11100111",14545 => "10010000",14546 => "01101110",14547 => "11001000",14548 => "10110111",14549 => "01111100",14550 => "00100110",14551 => "10011110",14552 => "11110010",14553 => "01010111",14554 => "11110000",14555 => "01011110",14556 => "01110010",14557 => "10000010",14558 => "11011000",14559 => "01101110",14560 => "11110101",14561 => "10011111",14562 => "11111010",14563 => "10000100",14564 => "01101000",14565 => "11001101",14566 => "00110111",14567 => "01001101",14568 => "01000110",14569 => "01111110",14570 => "00100001",14571 => "10000111",14572 => "01110110",14573 => "11101111",14574 => "10101100",14575 => "11001001",14576 => "00001111",14577 => "01001001",14578 => "01110100",14579 => "10101110",14580 => "10010101",14581 => "01010110",14582 => "10110001",14583 => "00111111",14584 => "00000101",14585 => "00000101",14586 => "10101001",14587 => "00001000",14588 => "01000010",14589 => "11001110",14590 => "00100111",14591 => "01110110",14592 => "10100101",14593 => "11001111",14594 => "11001000",14595 => "10100001",14596 => "11101110",14597 => "10010111",14598 => "11001111",14599 => "01010101",14600 => "01101011",14601 => "10011111",14602 => "10111011",14603 => "01110100",14604 => "10001110",14605 => "01101111",14606 => "10110101",14607 => "00110101",14608 => "11000100",14609 => "10111010",14610 => "10000100",14611 => "11010110",14612 => "11101010",14613 => "10111011",14614 => "00111110",14615 => "10000110",14616 => "11000110",14617 => "11001010",14618 => "10011100",14619 => "10000001",14620 => "11111001",14621 => "00100000",14622 => "00100010",14623 => "10001111",14624 => "10001111",14625 => "10000011",14626 => "00001111",14627 => "10111110",14628 => "01101111",14629 => "10111100",14630 => "11000011",14631 => "00011011",14632 => "11101100",14633 => "11100101",14634 => "00010011",14635 => "11000010",14636 => "00000010",14637 => "11100000",14638 => "10100100",14639 => "10011000",14640 => "11001100",14641 => "01000100",14642 => "10111011",14643 => "01101101",14644 => "00001101",14645 => "10101001",14646 => "00101111",14647 => "11011111",14648 => "11010011",14649 => "10011110",14650 => "00000011",14651 => "11101100",14652 => "11010111",14653 => "11001100",14654 => "10100000",14655 => "10010111",14656 => "01010011",14657 => "10101101",14658 => "10000001",14659 => "01010011",14660 => "11100101",14661 => "00011000",14662 => "10101010",14663 => "11000000",14664 => "00000001",14665 => "11110010",14666 => "00110000",14667 => "11000000",14668 => "01010011",14669 => "01000111",14670 => "11110010",14671 => "11101110",14672 => "00010110",14673 => "11010111",14674 => "00111001",14675 => "11101100",14676 => "01001010",14677 => "01010101",14678 => "10111011",14679 => "11011010",14680 => "11010000",14681 => "11111111",14682 => "01110110",14683 => "10001001",14684 => "10001111",14685 => "10101001",14686 => "00000000",14687 => "01010001",14688 => "01000001",14689 => "00111010",14690 => "10000000",14691 => "01000000",14692 => "01010010",14693 => "10100100",14694 => "11111001",14695 => "11010101",14696 => "10001011",14697 => "10101110",14698 => "00001111",14699 => "10110011",14700 => "00100000",14701 => "00000101",14702 => "10000101",14703 => "10011100",14704 => "01100010",14705 => "01101101",14706 => "00111111",14707 => "00011011",14708 => "01010001",14709 => "11111011",14710 => "11110111",14711 => "10111110",14712 => "00110001",14713 => "01000010",14714 => "10111011",14715 => "00010011",14716 => "00110011",14717 => "00001110",14718 => "01000101",14719 => "11110000",14720 => "10101110",14721 => "10101110",14722 => "00111111",14723 => "00110000",14724 => "11100110",14725 => "10110101",14726 => "00010000",14727 => "11100111",14728 => "00001001",14729 => "01011111",14730 => "01011111",14731 => "01000010",14732 => "01001011",14733 => "01010110",14734 => "10111111",14735 => "00000100",14736 => "01000011",14737 => "10101011",14738 => "00100111",14739 => "11100010",14740 => "01101000",14741 => "00001011",14742 => "00111111",14743 => "00101110",14744 => "00111011",14745 => "11110001",14746 => "11101010",14747 => "00001111",14748 => "00001001",14749 => "10001100",14750 => "01011011",14751 => "00011111",14752 => "11111001",14753 => "01101010",14754 => "00101111",14755 => "10100001",14756 => "11010010",14757 => "11000110",14758 => "01110101",14759 => "01000110",14760 => "00011110",14761 => "01110001",14762 => "00101011",14763 => "11001100",14764 => "10001000",14765 => "01100101",14766 => "10001011",14767 => "10010101",14768 => "00000111",14769 => "01101111",14770 => "00101100",14771 => "10111010",14772 => "10001010",14773 => "00110101",14774 => "00111010",14775 => "01110010",14776 => "00100100",14777 => "10100001",14778 => "11010110",14779 => "01010011",14780 => "00100000",14781 => "01011111",14782 => "11010011",14783 => "01001101",14784 => "01101111",14785 => "01101101",14786 => "00000000",14787 => "11001111",14788 => "11100110",14789 => "01101000",14790 => "01110100",14791 => "10001101",14792 => "00000010",14793 => "10000011",14794 => "11110110",14795 => "10000010",14796 => "11101011",14797 => "11100001",14798 => "10111010",14799 => "00010100",14800 => "11111110",14801 => "01111000",14802 => "00101100",14803 => "11101010",14804 => "11000111",14805 => "01101101",14806 => "00100010",14807 => "11010110",14808 => "01010101",14809 => "10110101",14810 => "00101110",14811 => "10110010",14812 => "00000011",14813 => "01001010",14814 => "10000110",14815 => "10000100",14816 => "01101011",14817 => "00001010",14818 => "00100000",14819 => "10011010",14820 => "10010111",14821 => "10011101",14822 => "11000110",14823 => "10001010",14824 => "10000101",14825 => "01111000",14826 => "11100011",14827 => "01110101",14828 => "10000001",14829 => "11110000",14830 => "10011011",14831 => "01011011",14832 => "10110001",14833 => "01101011",14834 => "01111111",14835 => "11010100",14836 => "11100110",14837 => "10010010",14838 => "00110011",14839 => "10001110",14840 => "11000101",14841 => "11101100",14842 => "00000000",14843 => "11010010",14844 => "00101010",14845 => "11101100",14846 => "00101011",14847 => "11001111",14848 => "10010110",14849 => "00110100",14850 => "00100111",14851 => "10010001",14852 => "11010001",14853 => "01001100",14854 => "10001100",14855 => "10011101",14856 => "10000010",14857 => "01101011",14858 => "10100001",14859 => "00000111",14860 => "00011010",14861 => "11000001",14862 => "00000010",14863 => "00000001",14864 => "11101011",14865 => "11101000",14866 => "00111000",14867 => "00101111",14868 => "01110101",14869 => "00000011",14870 => "00111011",14871 => "00010101",14872 => "10000000",14873 => "11010111",14874 => "01001101",14875 => "10111001",14876 => "11001100",14877 => "00111010",14878 => "10010011",14879 => "00010000",14880 => "01100011",14881 => "11111011",14882 => "10100101",14883 => "00011111",14884 => "11101110",14885 => "01010011",14886 => "10010110",14887 => "10001101",14888 => "01111001",14889 => "00100011",14890 => "00010000",14891 => "10101001",14892 => "01110011",14893 => "01001101",14894 => "01010111",14895 => "10001010",14896 => "00111010",14897 => "01110111",14898 => "00000000",14899 => "01110011",14900 => "00100110",14901 => "01011001",14902 => "00001110",14903 => "10010000",14904 => "11010000",14905 => "00010011",14906 => "10011000",14907 => "01101010",14908 => "00001010",14909 => "00101000",14910 => "01010101",14911 => "11001111",14912 => "01111000",14913 => "11101111",14914 => "01100111",14915 => "11110101",14916 => "01100101",14917 => "11011110",14918 => "10001011",14919 => "00000011",14920 => "10101011",14921 => "01110111",14922 => "01001110",14923 => "00110001",14924 => "00110010",14925 => "00000111",14926 => "11110010",14927 => "10000010",14928 => "00100101",14929 => "10100101",14930 => "11001101",14931 => "10011010",14932 => "10110001",14933 => "00011000",14934 => "01101110",14935 => "11100110",14936 => "00000011",14937 => "01110110",14938 => "00101000",14939 => "10010010",14940 => "10011010",14941 => "00101000",14942 => "10101001",14943 => "11110110",14944 => "11011101",14945 => "01111011",14946 => "11100011",14947 => "01000100",14948 => "01100111",14949 => "10000000",14950 => "11001100",14951 => "00100100",14952 => "10011110",14953 => "01001100",14954 => "10000101",14955 => "11111011",14956 => "01010110",14957 => "01110111",14958 => "11100011",14959 => "01100011",14960 => "10111110",14961 => "11011111",14962 => "11111011",14963 => "10011000",14964 => "11100010",14965 => "11100001",14966 => "10100111",14967 => "01110101",14968 => "10100010",14969 => "01010011",14970 => "01010011",14971 => "11000101",14972 => "11010110",14973 => "10011000",14974 => "01010001",14975 => "01000101",14976 => "11110010",14977 => "01100100",14978 => "00010110",14979 => "11001011",14980 => "00110010",14981 => "10001101",14982 => "10111011",14983 => "01010110",14984 => "01010000",14985 => "11100110",14986 => "01000111",14987 => "01110000",14988 => "10001011",14989 => "10100000",14990 => "01001100",14991 => "11101000",14992 => "11000010",14993 => "11111000",14994 => "10011111",14995 => "11110101",14996 => "01111011",14997 => "11100111",14998 => "01110101",14999 => "10000000",15000 => "11000000",15001 => "10011111",15002 => "11011100",15003 => "10000001",15004 => "00110100",15005 => "11111101",15006 => "01001100",15007 => "00110000",15008 => "10101110",15009 => "11001001",15010 => "11000100",15011 => "11000000",15012 => "11010000",15013 => "10100001",15014 => "00110111",15015 => "11101100",15016 => "00010110",15017 => "10110111",15018 => "00000101",15019 => "11001011",15020 => "00111101",15021 => "10000011",15022 => "11000011",15023 => "11100010",15024 => "00100101",15025 => "10011111",15026 => "10011000",15027 => "01001111",15028 => "10101000",15029 => "01001101",15030 => "01010100",15031 => "00110010",15032 => "11001001",15033 => "00101111",15034 => "01110010",15035 => "01111000",15036 => "10101001",15037 => "00010100",15038 => "00001100",15039 => "10110100",15040 => "10111000",15041 => "10101111",15042 => "11110101",15043 => "10111100",15044 => "11110001",15045 => "00100001",15046 => "01010011",15047 => "01100001",15048 => "01111001",15049 => "00100011",15050 => "01000101",15051 => "10011101",15052 => "00001001",15053 => "11101000",15054 => "11011010",15055 => "00111000",15056 => "10110011",15057 => "11000000",15058 => "00011011",15059 => "11111001",15060 => "10101100",15061 => "11111100",15062 => "11011110",15063 => "01010010",15064 => "00011111",15065 => "10000101",15066 => "00001010",15067 => "11101110",15068 => "00110110",15069 => "11011110",15070 => "01000001",15071 => "11000110",15072 => "10101011",15073 => "00011101",15074 => "00010110",15075 => "10101110",15076 => "11100010",15077 => "00101011",15078 => "10011111",15079 => "11100000",15080 => "10011101",15081 => "00000110",15082 => "00010101",15083 => "00000000",15084 => "10100000",15085 => "11000100",15086 => "11110100",15087 => "10000100",15088 => "11100110",15089 => "00100011",15090 => "11110101",15091 => "01010001",15092 => "11001101",15093 => "11100101",15094 => "11010000",15095 => "11110101",15096 => "10111011",15097 => "01110000",15098 => "00001010",15099 => "01010100",15100 => "00010100",15101 => "01000000",15102 => "01011100",15103 => "11001011",15104 => "00001000",15105 => "10000110",15106 => "11110101",15107 => "10100100",15108 => "11110001",15109 => "01000110",15110 => "11010100",15111 => "00100101",15112 => "11000011",15113 => "11111000",15114 => "10010010",15115 => "11100010",15116 => "10001011",15117 => "01101011",15118 => "01000110",15119 => "01000111",15120 => "01111011",15121 => "00001100",15122 => "10111101",15123 => "01110100",15124 => "01011100",15125 => "00111111",15126 => "10100000",15127 => "10101110",15128 => "11100101",15129 => "11110000",15130 => "10001011",15131 => "00101001",15132 => "11010000",15133 => "10111000",15134 => "00100001",15135 => "00011110",15136 => "00101111",15137 => "01000111",15138 => "00110001",15139 => "01000100",15140 => "00100100",15141 => "00110000",15142 => "01111100",15143 => "10100011",15144 => "00001111",15145 => "10110100",15146 => "00000110",15147 => "11010001",15148 => "01011111",15149 => "10100010",15150 => "01011010",15151 => "00011000",15152 => "11001001",15153 => "01100010",15154 => "01010001",15155 => "01100101",15156 => "10110101",15157 => "10010100",15158 => "01001001",15159 => "01001010",15160 => "00001110",15161 => "10100001",15162 => "11010101",15163 => "11001110",15164 => "01000010",15165 => "00010111",15166 => "00101011",15167 => "11111111",15168 => "01110101",15169 => "10000000",15170 => "01011000",15171 => "11100011",15172 => "10011001",15173 => "10111001",15174 => "00100001",15175 => "11111110",15176 => "10100011",15177 => "01111001",15178 => "10101001",15179 => "10111001",15180 => "00010011",15181 => "00011100",15182 => "11010111",15183 => "10001110",15184 => "11010111",15185 => "00111111",15186 => "00011111",15187 => "01001000",15188 => "00110100",15189 => "00101111",15190 => "10111101",15191 => "01000010",15192 => "00010110",15193 => "10110101",15194 => "10110010",15195 => "01101100",15196 => "01100011",15197 => "00011011",15198 => "11111101",15199 => "00010010",15200 => "10101010",15201 => "00100001",15202 => "00110100",15203 => "00111110",15204 => "10100001",15205 => "00111011",15206 => "10010101",15207 => "00011011",15208 => "11110100",15209 => "10101111",15210 => "00010000",15211 => "01011001",15212 => "01001011",15213 => "01010110",15214 => "11101010",15215 => "10010101",15216 => "01100100",15217 => "01111010",15218 => "01010000",15219 => "01010100",15220 => "10110011",15221 => "00100111",15222 => "10010111",15223 => "01000010",15224 => "01000100",15225 => "10101011",15226 => "10000000",15227 => "10111111",15228 => "01110000",15229 => "00011100",15230 => "11010100",15231 => "00110101",15232 => "00011000",15233 => "01000101",15234 => "10010010",15235 => "01001101",15236 => "10111111",15237 => "10010110",15238 => "00010100",15239 => "01011010",15240 => "10010101",15241 => "01100001",15242 => "01101101",15243 => "00100111",15244 => "10001101",15245 => "00001100",15246 => "01010010",15247 => "00110000",15248 => "01100010",15249 => "10001001",15250 => "00011010",15251 => "01010110",15252 => "01100010",15253 => "11110100",15254 => "11100110",15255 => "00110100",15256 => "00001101",15257 => "01111001",15258 => "11001001",15259 => "11001001",15260 => "00111100",15261 => "01101010",15262 => "00000000",15263 => "00101001",15264 => "01010010",15265 => "11101101",15266 => "00000000",15267 => "11100011",15268 => "01110111",15269 => "00111011",15270 => "11000000",15271 => "00000011",15272 => "10001000",15273 => "00000100",15274 => "10101110",15275 => "01000010",15276 => "11010101",15277 => "00000000",15278 => "01101111",15279 => "00000111",15280 => "11001111",15281 => "10100000",15282 => "00010111",15283 => "10111000",15284 => "11100110",15285 => "01100011",15286 => "10011000",15287 => "10001100",15288 => "10100011",15289 => "10010001",15290 => "01011101",15291 => "01100011",15292 => "01010110",15293 => "00111010",15294 => "11111100",15295 => "11011000",15296 => "01011101",15297 => "01111100",15298 => "10111011",15299 => "11100000",15300 => "11101110",15301 => "10000111",15302 => "11001101",15303 => "00111100",15304 => "10010010",15305 => "01100110",15306 => "11001110",15307 => "11010110",15308 => "10011001",15309 => "01011000",15310 => "01000101",15311 => "00111100",15312 => "11001011",15313 => "00000111",15314 => "00101110",15315 => "11111111",15316 => "10101111",15317 => "00111100",15318 => "11010000",15319 => "00010111",15320 => "11101100",15321 => "11001011",15322 => "11100110",15323 => "01110010",15324 => "01001001",15325 => "01101011",15326 => "00111110",15327 => "01111111",15328 => "11001001",15329 => "11001100",15330 => "11100011",15331 => "11010011",15332 => "00011011",15333 => "11110110",15334 => "00010000",15335 => "11100111",15336 => "11011010",15337 => "10100001",15338 => "10000011",15339 => "00010010",15340 => "00110001",15341 => "11111101",15342 => "10010100",15343 => "10011111",15344 => "01100011",15345 => "01001011",15346 => "01101000",15347 => "01110001",15348 => "01101010",15349 => "01100011",15350 => "11011111",15351 => "00110100",15352 => "10011101",15353 => "11110011",15354 => "00100000",15355 => "10100111",15356 => "01001010",15357 => "10101110",15358 => "11100111",15359 => "11011110",15360 => "10111111",15361 => "01010000",15362 => "01101001",15363 => "11111001",15364 => "01011100",15365 => "00000101",15366 => "11001010",15367 => "01110111",15368 => "10101101",15369 => "00010110",15370 => "11100001",15371 => "01011110",15372 => "10100100",15373 => "00010101",15374 => "01011001",15375 => "11011110",15376 => "01100011",15377 => "00101100",15378 => "11101100",15379 => "00000000",15380 => "11110000",15381 => "00000010",15382 => "01011000",15383 => "01000011",15384 => "11101011",15385 => "00100100",15386 => "00110001",15387 => "01011110",15388 => "11000001",15389 => "10001101",15390 => "01000111",15391 => "11010011",15392 => "10011110",15393 => "11100000",15394 => "01110100",15395 => "00110010",15396 => "11101011",15397 => "01101111",15398 => "10101000",15399 => "11100000",15400 => "10000011",15401 => "10010101",15402 => "11011101",15403 => "01000111",15404 => "10011110",15405 => "00011101",15406 => "11110111",15407 => "00110001",15408 => "11000000",15409 => "00001001",15410 => "00010011",15411 => "10110011",15412 => "10110111",15413 => "00111110",15414 => "00010110",15415 => "00000011",15416 => "10110000",15417 => "10111111",15418 => "10001111",15419 => "00001001",15420 => "11101101",15421 => "10101111",15422 => "10000101",15423 => "00010111",15424 => "01001010",15425 => "10101011",15426 => "11101001",15427 => "10100001",15428 => "10100000",15429 => "11111111",15430 => "11101000",15431 => "10100101",15432 => "10100010",15433 => "00010011",15434 => "01011111",15435 => "11110100",15436 => "10110111",15437 => "10110100",15438 => "10110001",15439 => "11101001",15440 => "10111010",15441 => "01101101",15442 => "10110000",15443 => "00110110",15444 => "10110100",15445 => "01010010",15446 => "10111101",15447 => "10101010",15448 => "00111110",15449 => "01001111",15450 => "10111001",15451 => "01111110",15452 => "01000011",15453 => "10000000",15454 => "01011100",15455 => "00011110",15456 => "10111001",15457 => "01000000",15458 => "00100001",15459 => "01011010",15460 => "00111001",15461 => "00011110",15462 => "00100011",15463 => "00100001",15464 => "10111110",15465 => "01100100",15466 => "10111101",15467 => "11110001",15468 => "00011110",15469 => "00010000",15470 => "00110111",15471 => "11000001",15472 => "10111100",15473 => "00001001",15474 => "00011100",15475 => "01011001",15476 => "01001110",15477 => "11001100",15478 => "11111101",15479 => "01111001",15480 => "01001011",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00111100" report "FAIL high bits" severity failure;
assert RAM(0) = "01111000" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
