 library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
 
entity project_tb is
end project_tb;


architecture projecttb of project_tb is
constant c_CLOCK_PERIOD		: time := 15 ns;
signal   tb_done		: std_logic;
signal   mem_address		: std_logic_vector (15 downto 0) := (others => '0');
signal   tb_rst		    : std_logic := '0';
signal   tb_start		: std_logic := '0';
signal   tb_clk		    : std_logic := '0';
signal   mem_o_data,mem_i_data		: std_logic_vector (7 downto 0);
signal   enable_wire  		: std_logic;
signal   mem_we		: std_logic;

type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
signal RAM: ram_type := (2 => "11000101",3 => "00011100",4 => "01011111",5 => "10001001",6 => "00000000",7 => "10111111",8 => "00001111",9 => "10001010",10 => "10011101",11 => "10100001",12 => "01100100",13 => "00000100",14 => "00001101",15 => "11110001",16 => "10111101",17 => "01001111",18 => "00100100",19 => "01100000",20 => "11000111",21 => "11000011",22 => "11000001",23 => "11000110",24 => "01111001",25 => "11101100",26 => "00111111",27 => "10011101",28 => "10010101",29 => "00110111",30 => "00101110",31 => "11001100",32 => "10010010",33 => "10110010",34 => "11010001",35 => "11001000",36 => "00000010",37 => "01000111",38 => "00011010",39 => "01001101",40 => "01111001",41 => "01110001",42 => "00001001",43 => "01100010",44 => "11010001",45 => "10001111",46 => "11101000",47 => "01110010",48 => "10011011",49 => "10111101",50 => "00011000",51 => "11110000",52 => "01101001",53 => "01100011",54 => "10001101",55 => "00111000",56 => "00001101",57 => "00001111",58 => "01001000",59 => "11100101",60 => "11101100",61 => "00000010",62 => "00011001",63 => "00111110",64 => "00101000",65 => "10000110",66 => "00000001",67 => "00100010",68 => "11100010",69 => "00010000",70 => "10011100",71 => "11110000",72 => "01111110",73 => "00001111",74 => "01100011",75 => "11110010",76 => "01101000",77 => "10111011",78 => "10010101",79 => "00011110",80 => "11001111",81 => "00011110",82 => "10110100",83 => "10101100",84 => "01011110",85 => "11011111",86 => "01101011",87 => "10011011",88 => "10111000",89 => "11011110",90 => "00010001",91 => "01111111",92 => "10001011",93 => "11111101",94 => "00100000",95 => "00001010",96 => "01101100",97 => "11011110",98 => "00010001",99 => "11111001",100 => "00001110",101 => "01011100",102 => "00000001",103 => "10000000",104 => "01100111",105 => "10010010",106 => "11110000",107 => "10110101",108 => "11001010",109 => "11100111",110 => "10110011",111 => "10010110",112 => "00110101",113 => "10001101",114 => "10100010",115 => "00001001",116 => "10110000",117 => "10011101",118 => "01111001",119 => "11010011",120 => "10110101",121 => "11001010",122 => "00000110",123 => "11011111",124 => "10100111",125 => "11100100",126 => "11010101",127 => "01010100",128 => "11001010",129 => "11101011",130 => "00010001",131 => "11010100",132 => "01011100",133 => "11000111",134 => "11010101",135 => "10101000",136 => "10111101",137 => "01000011",138 => "10010101",139 => "00100110",140 => "01110111",141 => "10011010",142 => "01010111",143 => "00011100",144 => "10101101",145 => "00110111",146 => "10100110",147 => "11011001",148 => "11100101",149 => "00010010",150 => "00011111",151 => "00100001",152 => "00100110",153 => "10100110",154 => "11010010",155 => "11110111",156 => "00100100",157 => "00111000",158 => "10000011",159 => "00010010",160 => "10111100",161 => "00101101",162 => "11001011",163 => "00001010",164 => "11101110",165 => "01110100",166 => "01110000",167 => "01101001",168 => "11000111",169 => "10001110",170 => "11001111",171 => "01011111",172 => "00110000",173 => "01111111",174 => "11010011",175 => "11110001",176 => "10101001",177 => "01010011",178 => "01000000",179 => "10010001",180 => "01110110",181 => "00000111",182 => "01001000",183 => "11010100",184 => "10010000",185 => "11011001",186 => "00001010",187 => "11101101",188 => "11111110",189 => "10100111",190 => "10000101",191 => "11000000",192 => "00001000",193 => "10101111",194 => "11011011",195 => "10111001",196 => "11001100",197 => "00110101",198 => "10111010",199 => "00001100",200 => "11110101",201 => "00010111",202 => "01010111",203 => "10000110",204 => "11100010",205 => "00011110",206 => "11110100",207 => "01001101",208 => "01001010",209 => "11011010",210 => "00111010",211 => "01101011",212 => "00010001",213 => "01011010",214 => "11010101",215 => "11100101",216 => "01110110",217 => "11011111",218 => "10111110",219 => "01010001",220 => "11000100",221 => "11110110",222 => "11110101",223 => "01000100",224 => "10011011",225 => "10111001",226 => "10000111",227 => "11110101",228 => "01001110",229 => "11110010",230 => "01010000",231 => "11111000",232 => "00100011",233 => "00101010",234 => "01101011",235 => "11110110",236 => "00001110",237 => "11000111",238 => "10010100",239 => "01111110",240 => "00110110",241 => "11001111",242 => "11011100",243 => "01000000",244 => "00101001",245 => "11111010",246 => "11101110",247 => "01000110",248 => "11001110",249 => "10000001",250 => "11010110",251 => "00001010",252 => "01100000",253 => "00010111",254 => "00111111",255 => "00001111",256 => "10101101",257 => "01110111",258 => "00011010",259 => "01111011",260 => "10111101",261 => "11000100",262 => "01101111",263 => "01010110",264 => "01111000",265 => "11001101",266 => "11011101",267 => "10011010",268 => "10111111",269 => "10100100",270 => "10100101",271 => "01000111",272 => "10010111",273 => "00101000",274 => "01000111",275 => "00011000",276 => "11110110",277 => "01110110",278 => "01010110",279 => "11011010",280 => "00100100",281 => "10001011",282 => "11001000",283 => "01100111",284 => "10011001",285 => "11111000",286 => "10100000",287 => "01110101",288 => "01011100",289 => "01001100",290 => "01101001",291 => "00110001",292 => "10001011",293 => "01100100",294 => "00001001",295 => "10101111",296 => "00000011",297 => "11100101",298 => "10110110",299 => "10101011",300 => "00111011",301 => "11010111",302 => "11011100",303 => "01000011",304 => "01110011",305 => "01111100",306 => "10111100",307 => "00001001",308 => "01111110",309 => "00100010",310 => "11101101",311 => "10110110",312 => "10010100",313 => "10100011",314 => "10010001",315 => "00001111",316 => "00010011",317 => "11000101",318 => "11101000",319 => "00101000",320 => "10000101",321 => "00100100",322 => "01010110",323 => "01011010",324 => "10110011",325 => "11111000",326 => "10110011",327 => "10100000",328 => "01000000",329 => "11001010",330 => "11001110",331 => "01100111",332 => "11111110",333 => "01101111",334 => "11001101",335 => "00010101",336 => "00100101",337 => "01001000",338 => "11011101",339 => "11001101",340 => "10101000",341 => "10001001",342 => "11010111",343 => "10100111",344 => "01101000",345 => "01110010",346 => "11001000",347 => "11101110",348 => "00100100",349 => "11000110",350 => "01101111",351 => "00111101",352 => "10010001",353 => "00110100",354 => "00111001",355 => "01100011",356 => "11111001",357 => "10000101",358 => "01011110",359 => "10011100",360 => "10000001",361 => "10001010",362 => "00110111",363 => "01110001",364 => "11100100",365 => "10100111",366 => "11001101",367 => "10001000",368 => "01100010",369 => "01101000",370 => "00111110",371 => "01000110",372 => "10110000",373 => "11001010",374 => "10001110",375 => "00011111",376 => "00110111",377 => "01000000",378 => "10111000",379 => "00100000",380 => "10110011",381 => "00111100",382 => "00111011",383 => "00000101",384 => "01011000",385 => "11010011",386 => "01101110",387 => "10100011",388 => "10101101",389 => "00101111",390 => "01110101",391 => "01100000",392 => "11001110",393 => "00001010",394 => "01010100",395 => "01111011",396 => "00111001",397 => "11010111",398 => "01001100",399 => "00010101",400 => "00010001",401 => "01011000",402 => "00110000",403 => "00011000",404 => "11111101",405 => "10011000",406 => "10011000",407 => "10100101",408 => "10011100",409 => "01111110",410 => "11010110",411 => "10101000",412 => "01100000",413 => "01010001",414 => "01100010",415 => "00011010",416 => "01001000",417 => "10010111",418 => "00111011",419 => "01101000",420 => "11011100",421 => "00110111",422 => "10000101",423 => "01100000",424 => "00110010",425 => "00000000",426 => "01000101",427 => "01001110",428 => "01011011",429 => "11111100",430 => "11100001",431 => "01100111",432 => "00100110",433 => "01101000",434 => "10010011",435 => "01101110",436 => "01100111",437 => "01101000",438 => "01101100",439 => "00100100",440 => "11001110",441 => "11110010",442 => "11111101",443 => "10101101",444 => "01110001",445 => "10000101",446 => "01010101",447 => "11100001",448 => "10101100",449 => "10111100",450 => "10001111",451 => "01101011",452 => "10101111",453 => "01000001",454 => "10010000",455 => "10000001",456 => "11111101",457 => "10110100",458 => "11000011",459 => "01110001",460 => "01010101",461 => "11101101",462 => "00010111",463 => "00111001",464 => "00100000",465 => "11111101",466 => "11110100",467 => "10000011",468 => "00101011",469 => "10010011",470 => "00000000",471 => "01011001",472 => "10111001",473 => "00001101",474 => "11011100",475 => "11011011",476 => "00010111",477 => "00110101",478 => "11110011",479 => "01100011",480 => "00010110",481 => "00011101",482 => "01111101",483 => "10010101",484 => "10011111",485 => "10011100",486 => "01101111",487 => "00001110",488 => "11101011",489 => "10000100",490 => "11101101",491 => "01011000",492 => "00010011",493 => "11011010",494 => "00100000",495 => "00101001",496 => "10100111",497 => "11010111",498 => "00011101",499 => "01100010",500 => "01011100",501 => "00101101",502 => "00001010",503 => "01001110",504 => "11001110",505 => "00001011",506 => "11110000",507 => "00000111",508 => "11110111",509 => "10001010",510 => "10100111",511 => "00100101",512 => "11100110",513 => "00000100",514 => "00011010",515 => "01100001",516 => "01110101",517 => "11110100",518 => "11001000",519 => "11011001",520 => "01000100",521 => "10111011",522 => "01000010",523 => "01010101",524 => "10011101",525 => "00011010",526 => "11111001",527 => "11001110",528 => "01110000",529 => "00010100",530 => "00010111",531 => "10111101",532 => "11101000",533 => "10101000",534 => "10101010",535 => "11101111",536 => "11011100",537 => "11101011",538 => "10110100",539 => "01110011",540 => "11101111",541 => "10111110",542 => "11111100",543 => "01110110",544 => "11000001",545 => "01111000",546 => "11010101",547 => "00110010",548 => "01100001",549 => "10100110",550 => "00011010",551 => "01100010",552 => "00100000",553 => "10111010",554 => "00111100",555 => "10111111",556 => "11010111",557 => "01111000",558 => "11101100",559 => "00100101",560 => "11100110",561 => "01010100",562 => "10101010",563 => "01100010",564 => "11000110",565 => "01000100",566 => "10110110",567 => "00111011",568 => "10110001",569 => "01100000",570 => "00101111",571 => "01010000",572 => "11010000",573 => "00100001",574 => "00001100",575 => "00110111",576 => "11011111",577 => "10100111",578 => "01010101",579 => "10100111",580 => "01101111",581 => "00001010",582 => "00001000",583 => "01001001",584 => "11111011",585 => "10001010",586 => "01100101",587 => "11010000",588 => "10000010",589 => "01101010",590 => "00111010",591 => "01100111",592 => "01100110",593 => "01100011",594 => "11111110",595 => "11101001",596 => "01110111",597 => "00011110",598 => "01111110",599 => "11010000",600 => "11001111",601 => "10001101",602 => "10100110",603 => "11111111",604 => "11000011",605 => "11011000",606 => "01110001",607 => "00110101",608 => "00111001",609 => "00101100",610 => "10110000",611 => "01011101",612 => "00000011",613 => "01110010",614 => "01000000",615 => "00110100",616 => "01010101",617 => "10101010",618 => "10110010",619 => "01101111",620 => "10111010",621 => "00110000",622 => "11111111",623 => "01011100",624 => "00011100",625 => "01011101",626 => "00101010",627 => "11100001",628 => "10100111",629 => "10011100",630 => "10011000",631 => "00100010",632 => "11110110",633 => "00111101",634 => "10110000",635 => "01101000",636 => "01001111",637 => "01001000",638 => "11101101",639 => "10110011",640 => "10110011",641 => "11101110",642 => "11100110",643 => "11100110",644 => "00101010",645 => "10011010",646 => "01011011",647 => "10010000",648 => "11000101",649 => "10010001",650 => "11100011",651 => "00100111",652 => "00011000",653 => "00101111",654 => "00100001",655 => "10111100",656 => "10000110",657 => "01110111",658 => "10110011",659 => "00111001",660 => "10010110",661 => "10000000",662 => "00001011",663 => "11001100",664 => "11110001",665 => "10011010",666 => "01000110",667 => "11001010",668 => "10111010",669 => "10011100",670 => "00000000",671 => "01100101",672 => "01011111",673 => "11010111",674 => "10001100",675 => "10000001",676 => "10100110",677 => "10000101",678 => "00111110",679 => "11111011",680 => "01110110",681 => "00110010",682 => "11011000",683 => "10100001",684 => "00101110",685 => "10111111",686 => "11101101",687 => "00111110",688 => "11111011",689 => "00100010",690 => "11011000",691 => "10010000",692 => "10100000",693 => "11100000",694 => "10000011",695 => "10001101",696 => "11110110",697 => "11101001",698 => "11101010",699 => "00111110",700 => "11000101",701 => "01100100",702 => "01100001",703 => "01110001",704 => "10010111",705 => "11111110",706 => "11101011",707 => "11000101",708 => "01100000",709 => "11011100",710 => "10000110",711 => "11101110",712 => "00010001",713 => "10000001",714 => "10100110",715 => "10001011",716 => "01000010",717 => "00010110",718 => "10110100",719 => "01110101",720 => "11110110",721 => "00111000",722 => "01010000",723 => "11000110",724 => "01010000",725 => "10000001",726 => "00111000",727 => "11000110",728 => "01001001",729 => "11101000",730 => "01011010",731 => "10001000",732 => "01111011",733 => "01111110",734 => "10101101",735 => "11110110",736 => "10101100",737 => "11001000",738 => "01100100",739 => "11010010",740 => "01111010",741 => "11010000",742 => "10010100",743 => "01100001",744 => "00000000",745 => "10101111",746 => "00000111",747 => "11010100",748 => "01010000",749 => "10110111",750 => "01101010",751 => "00100111",752 => "01110101",753 => "01011000",754 => "01010101",755 => "01001001",756 => "11011101",757 => "10011100",758 => "10101000",759 => "10111000",760 => "01000011",761 => "11011001",762 => "00101000",763 => "00000111",764 => "10101111",765 => "00110100",766 => "10110100",767 => "00001000",768 => "01010000",769 => "11101101",770 => "01101110",771 => "10101011",772 => "00001000",773 => "11011010",774 => "11010101",775 => "11110101",776 => "00000011",777 => "10001011",778 => "01011010",779 => "01100000",780 => "10111111",781 => "00100111",782 => "10100001",783 => "01110110",784 => "00001101",785 => "11011111",786 => "00111101",787 => "00110111",788 => "10001101",789 => "00010010",790 => "00100001",791 => "00100010",792 => "00110011",793 => "10101000",794 => "11001101",795 => "00000010",796 => "11010100",797 => "10011111",798 => "10001001",799 => "11101101",800 => "11011010",801 => "10101001",802 => "10011001",803 => "10001000",804 => "11000011",805 => "01001010",806 => "01011100",807 => "11111111",808 => "10010000",809 => "01010111",810 => "01000010",811 => "10101100",812 => "11111100",813 => "01111101",814 => "01001000",815 => "11011010",816 => "01010101",817 => "01100010",818 => "01011101",819 => "10001110",820 => "11111101",821 => "10000101",822 => "10011110",823 => "10010111",824 => "11000111",825 => "00010101",826 => "00111100",827 => "00011001",828 => "00111101",829 => "00010100",830 => "00111100",831 => "11011110",832 => "01111111",833 => "10111100",834 => "00100110",835 => "01111110",836 => "01111000",837 => "01011111",838 => "01000011",839 => "01101011",840 => "01011101",841 => "01001110",842 => "11100011",843 => "00101110",844 => "10011111",845 => "10111010",846 => "10001110",847 => "01010011",848 => "10000000",849 => "00111100",850 => "00000100",851 => "10100110",852 => "11001101",853 => "01001010",854 => "00101111",855 => "10101110",856 => "11111010",857 => "01100000",858 => "11010010",859 => "01001110",860 => "11001000",861 => "01010011",862 => "10000000",863 => "10001011",864 => "01110010",865 => "11000011",866 => "00111010",867 => "00110011",868 => "01110010",869 => "10010000",870 => "01101001",871 => "00100001",872 => "11001101",873 => "00100011",874 => "10010011",875 => "10010000",876 => "10100001",877 => "00001110",878 => "10100111",879 => "10101110",880 => "10110110",881 => "01111001",882 => "10001001",883 => "00001001",884 => "10000000",885 => "10100101",886 => "10000010",887 => "11111011",888 => "11011001",889 => "10110101",890 => "11100000",891 => "00011101",892 => "00111001",893 => "11011101",894 => "11010101",895 => "00010011",896 => "01000111",897 => "11111101",898 => "10000011",899 => "11011101",900 => "00010001",901 => "11110011",902 => "00111101",903 => "01101011",904 => "11101001",905 => "10101100",906 => "00111000",907 => "10011011",908 => "00000100",909 => "10110100",910 => "10101001",911 => "10010000",912 => "00000101",913 => "11111101",914 => "00101000",915 => "01110110",916 => "10010000",917 => "11110110",918 => "00111011",919 => "11110000",920 => "11101010",921 => "11000101",922 => "10100111",923 => "01110100",924 => "01101011",925 => "11111100",926 => "11100000",927 => "11011101",928 => "00001110",929 => "00011000",930 => "00001001",931 => "01001100",932 => "01111100",933 => "11000101",934 => "01001100",935 => "00110111",936 => "00101000",937 => "01001001",938 => "01000011",939 => "00001101",940 => "10011001",941 => "00101111",942 => "11111001",943 => "00011000",944 => "10101111",945 => "01111001",946 => "10111110",947 => "00010110",948 => "11011101",949 => "11010000",950 => "01000000",951 => "00000001",952 => "01100100",953 => "11001001",954 => "10010000",955 => "01111111",956 => "11001011",957 => "00010110",958 => "01111111",959 => "11001001",960 => "11011011",961 => "01100110",962 => "11000110",963 => "00011011",964 => "01011000",965 => "10110110",966 => "00001101",967 => "11100100",968 => "10111110",969 => "01001011",970 => "10100011",971 => "10110101",972 => "11111111",973 => "01001011",974 => "00111100",975 => "00101001",976 => "00001110",977 => "11100110",978 => "00101100",979 => "00000010",980 => "10001101",981 => "00111011",982 => "00101001",983 => "10010111",984 => "11101110",985 => "11010111",986 => "10111110",987 => "11101110",988 => "00111100",989 => "01011001",990 => "11000011",991 => "10010100",992 => "10100110",993 => "10001000",994 => "00110100",995 => "00110100",996 => "01101100",997 => "10000101",998 => "00100110",999 => "01101100",1000 => "11010011",1001 => "01001000",1002 => "00010111",1003 => "00101101",1004 => "10111111",1005 => "10100111",1006 => "11111011",1007 => "00111100",1008 => "01011101",1009 => "10101100",1010 => "00001110",1011 => "01000010",1012 => "11111100",1013 => "10000001",1014 => "00100011",1015 => "01101010",1016 => "10001001",1017 => "11001011",1018 => "10001111",1019 => "01110111",1020 => "11000011",1021 => "10011111",1022 => "01000110",1023 => "01101110",1024 => "11110101",1025 => "00000101",1026 => "10111000",1027 => "10011100",1028 => "01101101",1029 => "00110100",1030 => "11110000",1031 => "11100000",1032 => "10010111",1033 => "10011111",1034 => "00110010",1035 => "01100001",1036 => "01011001",1037 => "11101110",1038 => "01010011",1039 => "00110011",1040 => "00100100",1041 => "10000010",1042 => "01011101",1043 => "00011010",1044 => "11000110",1045 => "11100111",1046 => "10010000",1047 => "00101101",1048 => "01010001",1049 => "00000001",1050 => "01000001",1051 => "10101011",1052 => "10101010",1053 => "01001000",1054 => "01101000",1055 => "00101111",1056 => "00110101",1057 => "00010111",1058 => "00100101",1059 => "00101001",1060 => "11000001",1061 => "01010101",1062 => "10110111",1063 => "10000010",1064 => "10010101",1065 => "01101100",1066 => "10111000",1067 => "00000011",1068 => "00011100",1069 => "00101000",1070 => "01101010",1071 => "10001110",1072 => "11001110",1073 => "01110111",1074 => "10110001",1075 => "11100110",1076 => "10100010",1077 => "10111010",1078 => "11111111",1079 => "10001001",1080 => "00110100",1081 => "10000011",1082 => "11100001",1083 => "10101110",1084 => "00000101",1085 => "10000011",1086 => "00101101",1087 => "10110110",1088 => "10011111",1089 => "10010010",1090 => "00011101",1091 => "11101111",1092 => "00100001",1093 => "00011000",1094 => "00010100",1095 => "11111111",1096 => "10001101",1097 => "00010010",1098 => "10101000",1099 => "11011000",1100 => "10111011",1101 => "11110101",1102 => "01000110",1103 => "00111100",1104 => "11101101",1105 => "11101111",1106 => "00010001",1107 => "10011101",1108 => "00110101",1109 => "00001111",1110 => "01101001",1111 => "10001010",1112 => "01010000",1113 => "00011100",1114 => "01101011",1115 => "01011001",1116 => "10100100",1117 => "11011010",1118 => "00101110",1119 => "00010110",1120 => "00001100",1121 => "01101011",1122 => "01010001",1123 => "10110000",1124 => "00001110",1125 => "00100100",1126 => "00100001",1127 => "10010110",1128 => "10010100",1129 => "11011110",1130 => "00111000",1131 => "10100000",1132 => "01110011",1133 => "10001100",1134 => "10000000",1135 => "11000011",1136 => "01001101",1137 => "11100000",1138 => "00110110",1139 => "01110111",1140 => "10100100",1141 => "11100110",1142 => "01101010",1143 => "00011101",1144 => "11110111",1145 => "11000100",1146 => "00011101",1147 => "00110111",1148 => "10101100",1149 => "11011110",1150 => "00000001",1151 => "11100011",1152 => "11110101",1153 => "11010000",1154 => "00110011",1155 => "10000111",1156 => "01010101",1157 => "10011011",1158 => "11101110",1159 => "10011010",1160 => "01000000",1161 => "01111010",1162 => "11011110",1163 => "11010001",1164 => "01100101",1165 => "01011110",1166 => "10100010",1167 => "00110100",1168 => "10110001",1169 => "11011111",1170 => "00111101",1171 => "01011010",1172 => "01000010",1173 => "11011001",1174 => "01101110",1175 => "11110100",1176 => "00111111",1177 => "10101000",1178 => "10100000",1179 => "01010111",1180 => "01010010",1181 => "00010111",1182 => "00111111",1183 => "11001001",1184 => "01110010",1185 => "10000011",1186 => "11111010",1187 => "11101110",1188 => "01111011",1189 => "01101011",1190 => "00101000",1191 => "10011000",1192 => "11011111",1193 => "00011000",1194 => "01110000",1195 => "01111100",1196 => "00111000",1197 => "01110011",1198 => "11010010",1199 => "11000101",1200 => "00100011",1201 => "11101000",1202 => "10000111",1203 => "11110010",1204 => "11010010",1205 => "00001111",1206 => "01000111",1207 => "10110101",1208 => "00100011",1209 => "10011110",1210 => "10010010",1211 => "00000100",1212 => "10111010",1213 => "11111010",1214 => "11110100",1215 => "11100011",1216 => "00011011",1217 => "00001110",1218 => "01110000",1219 => "10011001",1220 => "10001110",1221 => "11101110",1222 => "11001001",1223 => "01100010",1224 => "00000111",1225 => "11100100",1226 => "11110110",1227 => "11111111",1228 => "01110101",1229 => "00000100",1230 => "01110010",1231 => "01010010",1232 => "10111111",1233 => "11110010",1234 => "11100100",1235 => "00000111",1236 => "00010100",1237 => "10110001",1238 => "11100011",1239 => "00100110",1240 => "01011010",1241 => "01000001",1242 => "00100111",1243 => "10000110",1244 => "11001001",1245 => "01111111",1246 => "00001001",1247 => "11110111",1248 => "11100000",1249 => "11101101",1250 => "10000000",1251 => "10010000",1252 => "10000011",1253 => "10011101",1254 => "01010000",1255 => "11100001",1256 => "11111010",1257 => "00110000",1258 => "10110001",1259 => "01100100",1260 => "11100001",1261 => "10100001",1262 => "11001111",1263 => "10101110",1264 => "11111100",1265 => "11111000",1266 => "00100000",1267 => "00000001",1268 => "11110000",1269 => "10010010",1270 => "10011011",1271 => "01101100",1272 => "01100010",1273 => "01001011",1274 => "00000000",1275 => "00101100",1276 => "01010101",1277 => "10010000",1278 => "11011111",1279 => "10001101",1280 => "00001111",1281 => "10001000",1282 => "01011010",1283 => "10001011",1284 => "10100100",1285 => "01001010",1286 => "11010111",1287 => "00001111",1288 => "11101001",1289 => "10110001",1290 => "11100010",1291 => "11001001",1292 => "01111011",1293 => "00010010",1294 => "11001011",1295 => "11011011",1296 => "10010010",1297 => "10011001",1298 => "01101111",1299 => "01000010",1300 => "11000011",1301 => "01000111",1302 => "01100011",1303 => "11111111",1304 => "00101101",1305 => "01110010",1306 => "00100100",1307 => "00111101",1308 => "11110110",1309 => "11001111",1310 => "10110000",1311 => "00000011",1312 => "01000110",1313 => "11100000",1314 => "01001111",1315 => "01110001",1316 => "01100110",1317 => "01100011",1318 => "11000001",1319 => "10110011",1320 => "11101011",1321 => "10111001",1322 => "11001011",1323 => "11001000",1324 => "01000110",1325 => "00011100",1326 => "01100100",1327 => "01001011",1328 => "00011001",1329 => "10000011",1330 => "10110000",1331 => "00111000",1332 => "00001011",1333 => "11011001",1334 => "10100001",1335 => "00101011",1336 => "01001010",1337 => "01100001",1338 => "11010110",1339 => "00110011",1340 => "10000011",1341 => "10111100",1342 => "11010111",1343 => "00010111",1344 => "01010111",1345 => "10010111",1346 => "10011011",1347 => "11010101",1348 => "10100010",1349 => "10000010",1350 => "00100010",1351 => "10110001",1352 => "01011101",1353 => "01001100",1354 => "11011001",1355 => "10101110",1356 => "00111001",1357 => "11010111",1358 => "11010111",1359 => "10010110",1360 => "00000011",1361 => "01011111",1362 => "01100001",1363 => "11101110",1364 => "01000101",1365 => "00101110",1366 => "10100110",1367 => "00011010",1368 => "10100010",1369 => "11110001",1370 => "10111100",1371 => "10000101",1372 => "01111001",1373 => "11101110",1374 => "10000101",1375 => "00101011",1376 => "11111001",1377 => "11010110",1378 => "11001100",1379 => "11110010",1380 => "11000111",1381 => "11010010",1382 => "00011000",1383 => "01110011",1384 => "11001100",1385 => "11001101",1386 => "11111001",1387 => "10100100",1388 => "10011010",1389 => "01011111",1390 => "10011100",1391 => "01111110",1392 => "01100001",1393 => "11111000",1394 => "11011010",1395 => "00000101",1396 => "11011101",1397 => "00100010",1398 => "10010010",1399 => "00100110",1400 => "10011001",1401 => "01010101",1402 => "00111010",1403 => "11110111",1404 => "10010001",1405 => "00011100",1406 => "01101011",1407 => "01000010",1408 => "01110011",1409 => "11001101",1410 => "11101010",1411 => "11010010",1412 => "10100000",1413 => "00100110",1414 => "01010101",1415 => "00001110",1416 => "11000000",1417 => "10011110",1418 => "00111111",1419 => "10100101",1420 => "10101011",1421 => "01000111",1422 => "00010100",1423 => "10011111",1424 => "01111100",1425 => "10000100",1426 => "01011101",1427 => "00011110",1428 => "10110110",1429 => "01011100",1430 => "01000111",1431 => "01001110",1432 => "00011000",1433 => "00101101",1434 => "10101101",1435 => "11011000",1436 => "01100111",1437 => "10111001",1438 => "11000111",1439 => "10100101",1440 => "11111101",1441 => "10010111",1442 => "11110110",1443 => "11110110",1444 => "00000100",1445 => "10111110",1446 => "00110101",1447 => "00001111",1448 => "11111101",1449 => "00101111",1450 => "00110100",1451 => "10101110",1452 => "00011100",1453 => "10010011",1454 => "00000110",1455 => "10100100",1456 => "11100011",1457 => "11111000",1458 => "00010000",1459 => "11111110",1460 => "11000111",1461 => "01101000",1462 => "11000111",1463 => "00001100",1464 => "00111000",1465 => "01000011",1466 => "10101101",1467 => "00111110",1468 => "01010001",1469 => "10011011",1470 => "01010110",1471 => "11110111",1472 => "10101011",1473 => "01110010",1474 => "11101111",1475 => "01110000",1476 => "00001100",1477 => "01010010",1478 => "11000010",1479 => "00010001",1480 => "01110110",1481 => "01101010",1482 => "11011000",1483 => "00110010",1484 => "10010001",1485 => "11110100",1486 => "11000100",1487 => "00001000",1488 => "01100001",1489 => "01011000",1490 => "10000110",1491 => "10001001",1492 => "01110111",1493 => "00010000",1494 => "10010110",1495 => "10111000",1496 => "01000010",1497 => "01001101",1498 => "10100000",1499 => "00110100",1500 => "00110110",1501 => "10000001",1502 => "01100001",1503 => "00110111",1504 => "00100000",1505 => "10001110",1506 => "11000001",1507 => "10000100",1508 => "01111111",1509 => "11001110",1510 => "11000000",1511 => "01101110",1512 => "11010110",1513 => "00111101",1514 => "01011001",1515 => "00011101",1516 => "01110010",1517 => "01101110",1518 => "10110101",1519 => "11101111",1520 => "10110101",1521 => "11001010",1522 => "01011110",1523 => "00011000",1524 => "10101100",1525 => "01000001",1526 => "01000000",1527 => "00110001",1528 => "01000111",1529 => "11011101",1530 => "00000110",1531 => "11000010",1532 => "10001011",1533 => "00010000",1534 => "00011001",1535 => "01110001",1536 => "11010011",1537 => "10101111",1538 => "10011111",1539 => "11011101",1540 => "01010000",1541 => "01011000",1542 => "11110100",1543 => "01011110",1544 => "10101111",1545 => "00100101",1546 => "00000000",1547 => "11100011",1548 => "00001110",1549 => "11110000",1550 => "11001111",1551 => "10100100",1552 => "01001000",1553 => "11001111",1554 => "11111010",1555 => "01000100",1556 => "00101111",1557 => "11101011",1558 => "11100011",1559 => "10011011",1560 => "01111101",1561 => "11100110",1562 => "10011001",1563 => "01110110",1564 => "11000110",1565 => "01110101",1566 => "01010000",1567 => "01010010",1568 => "00100101",1569 => "11101000",1570 => "10110101",1571 => "10110010",1572 => "10111010",1573 => "00010111",1574 => "11011010",1575 => "10100111",1576 => "11011100",1577 => "10000001",1578 => "00000011",1579 => "01110010",1580 => "11111101",1581 => "00101001",1582 => "10111010",1583 => "01111110",1584 => "11011010",1585 => "01010110",1586 => "11001000",1587 => "01000010",1588 => "10000011",1589 => "11000010",1590 => "10110101",1591 => "01110111",1592 => "10001110",1593 => "00110100",1594 => "10100001",1595 => "11111111",1596 => "11011111",1597 => "00001100",1598 => "10001011",1599 => "00111100",1600 => "01010011",1601 => "01001000",1602 => "01000100",1603 => "01001111",1604 => "11000100",1605 => "01000000",1606 => "01010001",1607 => "10011011",1608 => "01101101",1609 => "00000011",1610 => "01101111",1611 => "11101111",1612 => "11000010",1613 => "11101000",1614 => "11100100",1615 => "01000100",1616 => "11100000",1617 => "11110000",1618 => "00101001",1619 => "01010001",1620 => "10001011",1621 => "00101000",1622 => "10111111",1623 => "01101110",1624 => "00111110",1625 => "00000001",1626 => "01000110",1627 => "10000001",1628 => "01111011",1629 => "01011110",1630 => "00000111",1631 => "00101010",1632 => "10000110",1633 => "01110100",1634 => "11011101",1635 => "11000001",1636 => "01010101",1637 => "00111010",1638 => "00110011",1639 => "11101100",1640 => "01100110",1641 => "00100010",1642 => "01001100",1643 => "10011011",1644 => "11111010",1645 => "10001110",1646 => "10100110",1647 => "01000011",1648 => "11010100",1649 => "11001111",1650 => "01000000",1651 => "11010000",1652 => "01001111",1653 => "10101111",1654 => "11000000",1655 => "10001101",1656 => "11000101",1657 => "00010111",1658 => "01100101",1659 => "00011101",1660 => "00001110",1661 => "11111010",1662 => "10100111",1663 => "01110111",1664 => "10010110",1665 => "10000101",1666 => "01000011",1667 => "10111110",1668 => "00000101",1669 => "11101010",1670 => "01000101",1671 => "10001000",1672 => "11011100",1673 => "01001000",1674 => "10110010",1675 => "01010111",1676 => "10111100",1677 => "10001010",1678 => "10001011",1679 => "10001100",1680 => "10101111",1681 => "00001000",1682 => "11110110",1683 => "11010000",1684 => "00110111",1685 => "11001010",1686 => "11000100",1687 => "11101000",1688 => "00101000",1689 => "11010100",1690 => "11001001",1691 => "10100111",1692 => "11001110",1693 => "00001101",1694 => "11001001",1695 => "01111110",1696 => "01010011",1697 => "01101111",1698 => "00011000",1699 => "00101111",1700 => "11100011",1701 => "10111101",1702 => "01101101",1703 => "11010110",1704 => "01101010",1705 => "01110010",1706 => "11101101",1707 => "10110101",1708 => "01110010",1709 => "01111011",1710 => "11101110",1711 => "01000111",1712 => "10010110",1713 => "00001011",1714 => "11000100",1715 => "11111100",1716 => "11111100",1717 => "10101101",1718 => "11000110",1719 => "00001101",1720 => "11110011",1721 => "00111110",1722 => "10111101",1723 => "01000111",1724 => "11101101",1725 => "10000100",1726 => "01010000",1727 => "00101011",1728 => "01010011",1729 => "00101000",1730 => "00110111",1731 => "00000010",1732 => "10011100",1733 => "11100010",1734 => "10101010",1735 => "00111100",1736 => "10110000",1737 => "10001100",1738 => "01101000",1739 => "10100110",1740 => "11101000",1741 => "11101100",1742 => "01010110",1743 => "01001110",1744 => "01001010",1745 => "11111010",1746 => "11110011",1747 => "01101100",1748 => "01110010",1749 => "00000010",1750 => "00011110",1751 => "11110101",1752 => "11101100",1753 => "01111011",1754 => "01011001",1755 => "01110000",1756 => "01001100",1757 => "00100101",1758 => "11010011",1759 => "10001100",1760 => "01000110",1761 => "11100111",1762 => "01001110",1763 => "10100100",1764 => "01111111",1765 => "00010011",1766 => "00000001",1767 => "10100111",1768 => "11001010",1769 => "11001001",1770 => "11000000",1771 => "01010110",1772 => "01010000",1773 => "11100100",1774 => "10000111",1775 => "11000001",1776 => "01001001",1777 => "10001100",1778 => "01010110",1779 => "00011000",1780 => "00111100",1781 => "00101001",1782 => "11110111",1783 => "01100011",1784 => "10111111",1785 => "11111000",1786 => "00011101",1787 => "11000111",1788 => "00100111",1789 => "00110111",1790 => "01110000",1791 => "10100111",1792 => "10101110",1793 => "11001111",1794 => "01101100",1795 => "00100100",1796 => "00000110",1797 => "00000100",1798 => "10100111",1799 => "11001101",1800 => "10010100",1801 => "10010100",1802 => "11000111",1803 => "10100010",1804 => "01111101",1805 => "01011010",1806 => "00001011",1807 => "11110011",1808 => "10111101",1809 => "11011001",1810 => "11000011",1811 => "10100010",1812 => "01101100",1813 => "11010001",1814 => "11000100",1815 => "11110001",1816 => "10101111",1817 => "11100100",1818 => "10101101",1819 => "01011110",1820 => "11110011",1821 => "11001111",1822 => "01001111",1823 => "01100010",1824 => "01100011",1825 => "10011001",1826 => "10111010",1827 => "00111110",1828 => "00001010",1829 => "00100101",1830 => "01000001",1831 => "11110111",1832 => "01010000",1833 => "00011100",1834 => "11011101",1835 => "00110100",1836 => "01100010",1837 => "10001100",1838 => "10100011",1839 => "00100010",1840 => "10000101",1841 => "11100011",1842 => "00100001",1843 => "00100111",1844 => "10110100",1845 => "00111100",1846 => "10111110",1847 => "11101010",1848 => "01101011",1849 => "11000000",1850 => "00101011",1851 => "00000000",1852 => "10011101",1853 => "10000110",1854 => "10010011",1855 => "10110001",1856 => "11111100",1857 => "10010011",1858 => "11000110",1859 => "10101011",1860 => "11011000",1861 => "10100100",1862 => "11000001",1863 => "10111010",1864 => "01000111",1865 => "11111111",1866 => "01011110",1867 => "10011101",1868 => "10011100",1869 => "10010100",1870 => "11010001",1871 => "01110011",1872 => "10110110",1873 => "10100001",1874 => "11100110",1875 => "11001110",1876 => "10110010",1877 => "11001010",1878 => "10101000",1879 => "10011101",1880 => "11010101",1881 => "10100001",1882 => "10111001",1883 => "01011101",1884 => "11000011",1885 => "01100010",1886 => "11011000",1887 => "01100010",1888 => "01101011",1889 => "11010000",1890 => "10111010",1891 => "11111010",1892 => "01100000",1893 => "11100101",1894 => "11011010",1895 => "10110011",1896 => "00001101",1897 => "01001001",1898 => "10001111",1899 => "01001111",1900 => "11010010",1901 => "10101001",1902 => "11010010",1903 => "10000111",1904 => "11010100",1905 => "11010110",1906 => "01000000",1907 => "11000000",1908 => "01011010",1909 => "01101011",1910 => "11001001",1911 => "00101010",1912 => "01100001",1913 => "11101111",1914 => "00001001",1915 => "01110000",1916 => "01000111",1917 => "01010100",1918 => "10000111",1919 => "10011010",1920 => "10011100",1921 => "11111110",1922 => "01011101",1923 => "11011100",1924 => "10101110",1925 => "00000010",1926 => "10000100",1927 => "10000010",1928 => "01101000",1929 => "01010111",1930 => "10001110",1931 => "01011010",1932 => "10101110",1933 => "01011001",1934 => "00101011",1935 => "10010011",1936 => "10100000",1937 => "11011000",1938 => "01111000",1939 => "10010000",1940 => "11100101",1941 => "11100110",1942 => "10100101",1943 => "11110011",1944 => "01110110",1945 => "10101010",1946 => "11000111",1947 => "11000100",1948 => "10110101",1949 => "11000110",1950 => "01001010",1951 => "00100000",1952 => "11011110",1953 => "00110001",1954 => "01001110",1955 => "00001010",1956 => "10111100",1957 => "10010100",1958 => "01100111",1959 => "11100111",1960 => "00011000",1961 => "00001110",1962 => "00011111",1963 => "00000110",1964 => "01111011",1965 => "00111111",1966 => "11001000",1967 => "10101111",1968 => "00000111",1969 => "01111100",1970 => "00000110",1971 => "00010010",1972 => "10111110",1973 => "11001001",1974 => "01001101",1975 => "10110001",1976 => "00011101",1977 => "11001011",1978 => "00000000",1979 => "10011001",1980 => "11000110",1981 => "01010101",1982 => "00011100",1983 => "10101011",1984 => "01101010",1985 => "01011100",1986 => "11001110",1987 => "00000101",1988 => "01010011",1989 => "01100100",1990 => "00100001",1991 => "10000110",1992 => "11000000",1993 => "01001010",1994 => "00110011",1995 => "11110010",1996 => "10010011",1997 => "11100100",1998 => "10110011",1999 => "00100011",2000 => "10101011",2001 => "00111010",2002 => "01001000",2003 => "11110011",2004 => "10011100",2005 => "10111111",2006 => "00010000",2007 => "00001101",2008 => "01100010",2009 => "00111000",2010 => "01001111",2011 => "01100110",2012 => "11010101",2013 => "11100011",2014 => "00011001",2015 => "10001011",2016 => "01101110",2017 => "11101111",2018 => "11010010",2019 => "11001010",2020 => "01001101",2021 => "00010101",2022 => "11101000",2023 => "11101110",2024 => "01001010",2025 => "11000100",2026 => "11110001",2027 => "01111101",2028 => "10111110",2029 => "11100110",2030 => "00000111",2031 => "11010011",2032 => "00011111",2033 => "10111100",2034 => "10010111",2035 => "10010010",2036 => "01000111",2037 => "11001010",2038 => "11111000",2039 => "01000100",2040 => "01010010",2041 => "10000111",2042 => "11010100",2043 => "00011010",2044 => "01001111",2045 => "00011110",2046 => "10110100",2047 => "01111000",2048 => "10101111",2049 => "00110011",2050 => "00000001",2051 => "10111110",2052 => "00001100",2053 => "11000000",2054 => "01111000",2055 => "00010111",2056 => "01110011",2057 => "01110010",2058 => "00111110",2059 => "01001101",2060 => "10000110",2061 => "11100000",2062 => "01001000",2063 => "10111000",2064 => "00110100",2065 => "00000111",2066 => "00100111",2067 => "00000011",2068 => "11111111",2069 => "01010000",2070 => "10000111",2071 => "11100110",2072 => "01011011",2073 => "11100001",2074 => "10000110",2075 => "11001101",2076 => "00011001",2077 => "11011011",2078 => "01100011",2079 => "01000100",2080 => "11100100",2081 => "11110100",2082 => "00101000",2083 => "10000100",2084 => "01011101",2085 => "11010010",2086 => "10111100",2087 => "11010000",2088 => "01110011",2089 => "10010101",2090 => "10010110",2091 => "11111110",2092 => "00001001",2093 => "10100111",2094 => "01001100",2095 => "00010000",2096 => "11000111",2097 => "11101110",2098 => "11001001",2099 => "10111001",2100 => "10000111",2101 => "00000110",2102 => "01011111",2103 => "01011111",2104 => "00110010",2105 => "01010111",2106 => "01011011",2107 => "10011001",2108 => "11111000",2109 => "01111000",2110 => "10110001",2111 => "01011110",2112 => "10000101",2113 => "01100010",2114 => "11011011",2115 => "00110000",2116 => "00101100",2117 => "11001000",2118 => "11111000",2119 => "00011000",2120 => "10111010",2121 => "10100111",2122 => "11101100",2123 => "00010111",2124 => "00011001",2125 => "00100000",2126 => "10100011",2127 => "10111011",2128 => "11111011",2129 => "00011110",2130 => "00101110",2131 => "10000110",2132 => "01010011",2133 => "01110100",2134 => "10110110",2135 => "11100101",2136 => "00111101",2137 => "00011100",2138 => "00111010",2139 => "01111010",2140 => "00100010",2141 => "11000100",2142 => "01010110",2143 => "10111010",2144 => "10110010",2145 => "00010101",2146 => "00000111",2147 => "00101111",2148 => "01000001",2149 => "11000110",2150 => "10001110",2151 => "00010001",2152 => "10111001",2153 => "10001101",2154 => "10011100",2155 => "00010111",2156 => "10111111",2157 => "10001100",2158 => "00111011",2159 => "11000010",2160 => "11110001",2161 => "10010001",2162 => "11000000",2163 => "00100010",2164 => "01011000",2165 => "11000111",2166 => "10001010",2167 => "01100101",2168 => "00010001",2169 => "01001001",2170 => "11101011",2171 => "10011110",2172 => "00001000",2173 => "01101100",2174 => "11011011",2175 => "01111111",2176 => "11011110",2177 => "00010001",2178 => "10011100",2179 => "00010111",2180 => "00111101",2181 => "01111011",2182 => "10000100",2183 => "01100100",2184 => "10001010",2185 => "10001010",2186 => "11101110",2187 => "01000001",2188 => "00000001",2189 => "10011011",2190 => "10000100",2191 => "10101001",2192 => "10001100",2193 => "01101010",2194 => "11111111",2195 => "01001110",2196 => "00100100",2197 => "10010101",2198 => "01111100",2199 => "11111011",2200 => "01001011",2201 => "01100001",2202 => "10100110",2203 => "01100110",2204 => "01000001",2205 => "01101010",2206 => "10101001",2207 => "10110001",2208 => "11000101",2209 => "00001111",2210 => "11001100",2211 => "11011110",2212 => "10011100",2213 => "10110110",2214 => "01000110",2215 => "10100110",2216 => "00111010",2217 => "10110110",2218 => "01011101",2219 => "00001111",2220 => "11101010",2221 => "10111101",2222 => "00010011",2223 => "01000111",2224 => "01110010",2225 => "01010011",2226 => "10011000",2227 => "10101011",2228 => "11000001",2229 => "11010110",2230 => "00101101",2231 => "11010111",2232 => "01000111",2233 => "10101010",2234 => "01011001",2235 => "11100000",2236 => "10110101",2237 => "01101001",2238 => "01111100",2239 => "10001001",2240 => "11110101",2241 => "01001101",2242 => "00110101",2243 => "01100000",2244 => "10000100",2245 => "10011101",2246 => "10001001",2247 => "11100011",2248 => "10011100",2249 => "11011101",2250 => "00011011",2251 => "01011111",2252 => "00101100",2253 => "00001100",2254 => "10011000",2255 => "00111111",2256 => "00111001",2257 => "11101010",2258 => "11111010",2259 => "11111001",2260 => "01000000",2261 => "11101011",2262 => "01110000",2263 => "00111010",2264 => "10101110",2265 => "01001110",2266 => "10111011",2267 => "00010011",2268 => "10100011",2269 => "01101011",2270 => "00001110",2271 => "01101100",2272 => "11000011",2273 => "00011000",2274 => "11100110",2275 => "11111100",2276 => "01110001",2277 => "00110001",2278 => "01110001",2279 => "11010011",2280 => "01100001",2281 => "11110101",2282 => "00000100",2283 => "00111111",2284 => "00100010",2285 => "00000100",2286 => "01111010",2287 => "00001111",2288 => "01111100",2289 => "10011110",2290 => "01010011",2291 => "00101100",2292 => "00011010",2293 => "01001000",2294 => "11010010",2295 => "01111010",2296 => "00100100",2297 => "10101001",2298 => "00000101",2299 => "10101000",2300 => "10100001",2301 => "00111001",2302 => "11111010",2303 => "01111011",2304 => "10101110",2305 => "11001100",2306 => "01110000",2307 => "11000000",2308 => "11111110",2309 => "01010101",2310 => "00101100",2311 => "00110101",2312 => "10111000",2313 => "11100001",2314 => "01110010",2315 => "01001101",2316 => "01100000",2317 => "10110100",2318 => "10100010",2319 => "11010101",2320 => "11001000",2321 => "00101011",2322 => "00000111",2323 => "01101001",2324 => "01011101",2325 => "11101101",2326 => "00100001",2327 => "10100110",2328 => "00111100",2329 => "01111101",2330 => "11010000",2331 => "01110111",2332 => "11111010",2333 => "10101000",2334 => "10001011",2335 => "11110001",2336 => "00101101",2337 => "11000100",2338 => "11110010",2339 => "00010000",2340 => "01000110",2341 => "11010011",2342 => "00011000",2343 => "00101100",2344 => "00101011",2345 => "00100010",2346 => "00001000",2347 => "11000110",2348 => "11101001",2349 => "10101010",2350 => "11101011",2351 => "00111110",2352 => "10100000",2353 => "10010000",2354 => "00110011",2355 => "11001001",2356 => "11011110",2357 => "10010110",2358 => "00101010",2359 => "11100001",2360 => "00001001",2361 => "01100110",2362 => "01011110",2363 => "11000111",2364 => "01111010",2365 => "00000100",2366 => "11011101",2367 => "00100010",2368 => "01001110",2369 => "10101000",2370 => "00100100",2371 => "01110111",2372 => "10101101",2373 => "01010110",2374 => "00111101",2375 => "10011011",2376 => "11011111",2377 => "00010000",2378 => "01011111",2379 => "00001110",2380 => "00011011",2381 => "01000001",2382 => "01101110",2383 => "10101000",2384 => "00110110",2385 => "10101101",2386 => "10011100",2387 => "00001011",2388 => "01101111",2389 => "11111101",2390 => "10000111",2391 => "10000000",2392 => "11100011",2393 => "01000100",2394 => "01101001",2395 => "10011001",2396 => "01010110",2397 => "01111001",2398 => "11000010",2399 => "00110010",2400 => "10010010",2401 => "11000011",2402 => "00100011",2403 => "11111100",2404 => "00110101",2405 => "00001110",2406 => "01000100",2407 => "00100110",2408 => "00000011",2409 => "11011101",2410 => "10001000",2411 => "00001101",2412 => "10100001",2413 => "10110101",2414 => "10101111",2415 => "01110111",2416 => "01001001",2417 => "10010100",2418 => "11100001",2419 => "01100111",2420 => "01100001",2421 => "11001111",2422 => "00010100",2423 => "11001111",2424 => "10110001",2425 => "11100000",2426 => "10101011",2427 => "01010001",2428 => "11010110",2429 => "10101010",2430 => "11101101",2431 => "01011101",2432 => "10111100",2433 => "11110010",2434 => "10111000",2435 => "11100011",2436 => "00110011",2437 => "11010001",2438 => "01010000",2439 => "00001011",2440 => "01001100",2441 => "01111010",2442 => "00101100",2443 => "10000010",2444 => "10010011",2445 => "10000000",2446 => "10111010",2447 => "00111011",2448 => "10001010",2449 => "10011111",2450 => "11101101",2451 => "00010011",2452 => "00001001",2453 => "11100110",2454 => "00010011",2455 => "10011000",2456 => "10101001",2457 => "01101110",2458 => "01011001",2459 => "00010010",2460 => "10101110",2461 => "10011010",2462 => "10110100",2463 => "10100110",2464 => "01111001",2465 => "00000101",2466 => "01001010",2467 => "10110000",2468 => "01000011",2469 => "00100010",2470 => "11110011",2471 => "00110011",2472 => "10110110",2473 => "11010010",2474 => "10100110",2475 => "11011010",2476 => "11110111",2477 => "10101010",2478 => "10101111",2479 => "00111011",2480 => "11001010",2481 => "00100100",2482 => "01101001",2483 => "10101011",2484 => "11001001",2485 => "11100111",2486 => "00111100",2487 => "11001011",2488 => "00110010",2489 => "11101111",2490 => "00110101",2491 => "00110101",2492 => "00000111",2493 => "11100100",2494 => "11011110",2495 => "00100101",2496 => "11011111",2497 => "10010010",2498 => "01001001",2499 => "11110110",2500 => "01001111",2501 => "00101000",2502 => "10110000",2503 => "00111000",2504 => "01111010",2505 => "01110110",2506 => "00000100",2507 => "11100001",2508 => "11010011",2509 => "00101100",2510 => "11101101",2511 => "10111001",2512 => "11101100",2513 => "01111011",2514 => "01001110",2515 => "00100111",2516 => "01111001",2517 => "01100111",2518 => "11010011",2519 => "10100011",2520 => "00010000",2521 => "00011110",2522 => "00110111",2523 => "00011100",2524 => "01111010",2525 => "00101110",2526 => "00011110",2527 => "00011001",2528 => "11011110",2529 => "11011110",2530 => "11000001",2531 => "01001111",2532 => "10010110",2533 => "10001001",2534 => "11111000",2535 => "00100100",2536 => "10001011",2537 => "11101111",2538 => "00010000",2539 => "00101101",2540 => "11001110",2541 => "00101110",2542 => "11101101",2543 => "11001000",2544 => "01111000",2545 => "11110101",2546 => "10110011",2547 => "11011000",2548 => "00100110",2549 => "11001100",2550 => "00010010",2551 => "11010111",2552 => "11101101",2553 => "10101101",2554 => "11111100",2555 => "01001101",2556 => "10111100",2557 => "00001001",2558 => "10100110",2559 => "01001110",2560 => "00100100",2561 => "01111111",2562 => "11011011",2563 => "10011100",2564 => "10100001",2565 => "00110100",2566 => "11110001",2567 => "11100110",2568 => "11011010",2569 => "10100001",2570 => "01001011",2571 => "11010111",2572 => "11100101",2573 => "01000100",2574 => "01010010",2575 => "11110010",2576 => "00000011",2577 => "00110110",2578 => "00110100",2579 => "11000000",2580 => "10110011",2581 => "00111100",2582 => "11000000",2583 => "11010010",2584 => "11101001",2585 => "00110111",2586 => "10110010",2587 => "01001011",2588 => "00000100",2589 => "10010111",2590 => "01010100",2591 => "01110100",2592 => "11001001",2593 => "10110101",2594 => "11101001",2595 => "00100111",2596 => "00110011",2597 => "01100101",2598 => "00010110",2599 => "10011001",2600 => "00110110",2601 => "01100001",2602 => "01000101",2603 => "00110010",2604 => "11000101",2605 => "01100010",2606 => "11101010",2607 => "01010000",2608 => "10000111",2609 => "01100001",2610 => "11000000",2611 => "10111001",2612 => "01100011",2613 => "11111000",2614 => "01001010",2615 => "10110011",2616 => "00000010",2617 => "01011111",2618 => "10010110",2619 => "00111100",2620 => "00110111",2621 => "01010111",2622 => "10010000",2623 => "11011100",2624 => "10000110",2625 => "10010011",2626 => "00011000",2627 => "10101001",2628 => "10100011",2629 => "11010101",2630 => "11000110",2631 => "01011100",2632 => "11100100",2633 => "00001101",2634 => "10110010",2635 => "01111000",2636 => "10011100",2637 => "00110011",2638 => "10010101",2639 => "00100000",2640 => "01100110",2641 => "00110101",2642 => "11000000",2643 => "00001000",2644 => "00101110",2645 => "01010110",2646 => "10101110",2647 => "10011001",2648 => "00011011",2649 => "00111111",2650 => "00000110",2651 => "00011001",2652 => "01000011",2653 => "01110101",2654 => "00001001",2655 => "11000011",2656 => "11000101",2657 => "00101010",2658 => "10111011",2659 => "01100010",2660 => "00011010",2661 => "11001110",2662 => "01001000",2663 => "01101100",2664 => "11011100",2665 => "01111101",2666 => "11100101",2667 => "00011010",2668 => "11000110",2669 => "00110010",2670 => "01010101",2671 => "00011011",2672 => "01111111",2673 => "01101101",2674 => "10011101",2675 => "00100010",2676 => "11111010",2677 => "10011111",2678 => "01010010",2679 => "01100001",2680 => "00110111",2681 => "11101011",2682 => "11010011",2683 => "00001001",2684 => "11001110",2685 => "11010110",2686 => "01110001",2687 => "00110100",2688 => "10101010",2689 => "10111101",2690 => "11101001",2691 => "10110111",2692 => "10110101",2693 => "10100110",2694 => "10110001",2695 => "00101101",2696 => "01101111",2697 => "11010111",2698 => "00000001",2699 => "10100101",2700 => "01010101",2701 => "10101010",2702 => "11110011",2703 => "11001001",2704 => "01101010",2705 => "10100100",2706 => "01010011",2707 => "01001111",2708 => "10011111",2709 => "00010101",2710 => "01101100",2711 => "10011101",2712 => "00101000",2713 => "11100010",2714 => "00100001",2715 => "01000100",2716 => "10101011",2717 => "10010010",2718 => "01101101",2719 => "11111011",2720 => "11010011",2721 => "00101011",2722 => "10001001",2723 => "01011111",2724 => "00110011",2725 => "10110100",2726 => "11101100",2727 => "00100111",2728 => "10101110",2729 => "10011011",2730 => "01000000",2731 => "01101010",2732 => "01110110",2733 => "11010011",2734 => "11110101",2735 => "10100101",2736 => "00000000",2737 => "10101101",2738 => "10010000",2739 => "10110010",2740 => "11001111",2741 => "11000010",2742 => "00000101",2743 => "11010011",2744 => "00010011",2745 => "11011100",2746 => "11011111",2747 => "00110010",2748 => "00000001",2749 => "01110100",2750 => "01000111",2751 => "10101011",2752 => "01001011",2753 => "11000111",2754 => "10010111",2755 => "01011110",2756 => "01011010",2757 => "11001000",2758 => "00010001",2759 => "00110001",2760 => "01010010",2761 => "00111001",2762 => "11101101",2763 => "11110011",2764 => "00101011",2765 => "01011101",2766 => "10111000",2767 => "00010100",2768 => "11010100",2769 => "00010001",2770 => "10110110",2771 => "11011011",2772 => "01100100",2773 => "01101100",2774 => "00011101",2775 => "11100101",2776 => "11110110",2777 => "00001001",2778 => "01100011",2779 => "01111111",2780 => "00011001",2781 => "00000001",2782 => "01110011",2783 => "11010101",2784 => "00010110",2785 => "11001010",2786 => "00000110",2787 => "01110010",2788 => "10111010",2789 => "00110000",2790 => "11010111",2791 => "10101100",2792 => "00000010",2793 => "01110100",2794 => "11011001",2795 => "11111101",2796 => "00101101",2797 => "11111000",2798 => "00011011",2799 => "11100001",2800 => "11001100",2801 => "10110000",2802 => "00100110",2803 => "11110001",2804 => "10100100",2805 => "11101101",2806 => "01010011",2807 => "01111100",2808 => "00010000",2809 => "11100010",2810 => "10101100",2811 => "11011111",2812 => "10100110",2813 => "00000000",2814 => "00000011",2815 => "11011011",2816 => "00011101",2817 => "00101110",2818 => "11101001",2819 => "01111111",2820 => "10110011",2821 => "11000101",2822 => "10001010",2823 => "01110000",2824 => "11111011",2825 => "11011010",2826 => "11101001",2827 => "11100101",2828 => "01001011",2829 => "01011111",2830 => "11111011",2831 => "11010000",2832 => "11010011",2833 => "10101101",2834 => "10101001",2835 => "11001011",2836 => "01011101",2837 => "01101111",2838 => "10100001",2839 => "10111001",2840 => "00000010",2841 => "00000010",2842 => "11011111",2843 => "11000101",2844 => "01010111",2845 => "01110001",2846 => "10111110",2847 => "10111001",2848 => "01101011",2849 => "10100001",2850 => "01011101",2851 => "00000100",2852 => "10111010",2853 => "01101011",2854 => "11100110",2855 => "01000100",2856 => "00111010",2857 => "01000011",2858 => "01111110",2859 => "11001101",2860 => "01100011",2861 => "01001100",2862 => "00101100",2863 => "00101001",2864 => "01001111",2865 => "10011110",2866 => "10110110",2867 => "00111101",2868 => "00010000",2869 => "11000111",2870 => "11010100",2871 => "00011001",2872 => "11001010",2873 => "11000101",2874 => "00101111",2875 => "01000000",2876 => "00100101",2877 => "01001101",2878 => "01111000",2879 => "10111000",2880 => "11010101",2881 => "01100011",2882 => "00011111",2883 => "10011100",2884 => "01001111",2885 => "11111001",2886 => "11001110",2887 => "01110101",2888 => "11111110",2889 => "00101000",2890 => "01100000",2891 => "10001010",2892 => "01001101",2893 => "00101101",2894 => "00001001",2895 => "11001011",2896 => "11111011",2897 => "11110010",2898 => "01101011",2899 => "00000111",2900 => "01110100",2901 => "10000101",2902 => "10111101",2903 => "11110111",2904 => "00010001",2905 => "11001001",2906 => "10000101",2907 => "00101111",2908 => "10100100",2909 => "01111100",2910 => "10111101",2911 => "00010010",2912 => "11001001",2913 => "01011010",2914 => "11010010",2915 => "11011000",2916 => "10000111",2917 => "00011001",2918 => "10011110",2919 => "10000010",2920 => "11100101",2921 => "10011000",2922 => "01011101",2923 => "01000000",2924 => "10001111",2925 => "00001000",2926 => "11111100",2927 => "10010010",2928 => "01101010",2929 => "01110111",2930 => "00110111",2931 => "11011100",2932 => "10011011",2933 => "10010001",2934 => "11010101",2935 => "10010100",2936 => "00010011",2937 => "11010100",2938 => "11000101",2939 => "11101000",2940 => "10100110",2941 => "01001000",2942 => "11101110",2943 => "10101101",2944 => "11001111",2945 => "00111000",2946 => "10010011",2947 => "10101101",2948 => "10011010",2949 => "10100000",2950 => "10000001",2951 => "10001110",2952 => "01010110",2953 => "00001001",2954 => "10100110",2955 => "00110111",2956 => "00111000",2957 => "10000101",2958 => "11011000",2959 => "00101010",2960 => "00101010",2961 => "11100011",2962 => "00110111",2963 => "11001110",2964 => "00101100",2965 => "11000111",2966 => "00110010",2967 => "10011011",2968 => "11100001",2969 => "01001111",2970 => "11010011",2971 => "00011100",2972 => "10001111",2973 => "10010100",2974 => "00111001",2975 => "10001111",2976 => "00101011",2977 => "11011001",2978 => "11001010",2979 => "11110000",2980 => "01011000",2981 => "11001011",2982 => "11100000",2983 => "11001001",2984 => "01110110",2985 => "00110010",2986 => "11111110",2987 => "10000110",2988 => "01101011",2989 => "01011110",2990 => "00000011",2991 => "01111010",2992 => "10100101",2993 => "00110111",2994 => "01100010",2995 => "00011111",2996 => "10111001",2997 => "01001000",2998 => "11011011",2999 => "10001010",3000 => "10000000",3001 => "10011011",3002 => "01010100",3003 => "11001101",3004 => "11101000",3005 => "00001100",3006 => "10011101",3007 => "11000110",3008 => "00001011",3009 => "10001111",3010 => "10100110",3011 => "10100000",3012 => "01001111",3013 => "10100001",3014 => "11101100",3015 => "11110101",3016 => "00010011",3017 => "01111011",3018 => "00000100",3019 => "11111011",3020 => "10000110",3021 => "10010111",3022 => "01100010",3023 => "10100100",3024 => "11100001",3025 => "11001110",3026 => "11100111",3027 => "10110111",3028 => "10000110",3029 => "00110010",3030 => "00011010",3031 => "11110001",3032 => "01101001",3033 => "11110001",3034 => "00000101",3035 => "11111100",3036 => "11111010",3037 => "10000111",3038 => "11011100",3039 => "10101101",3040 => "11100000",3041 => "00110101",3042 => "00101111",3043 => "11001110",3044 => "10110010",3045 => "11010010",3046 => "00011110",3047 => "00100110",3048 => "10111111",3049 => "10101111",3050 => "11000111",3051 => "10101111",3052 => "10011011",3053 => "01000100",3054 => "10011011",3055 => "10001110",3056 => "00110001",3057 => "00010000",3058 => "10110100",3059 => "01011001",3060 => "10110010",3061 => "00001110",3062 => "10011001",3063 => "00100000",3064 => "01100010",3065 => "00110011",3066 => "11101011",3067 => "00101101",3068 => "00010000",3069 => "10110110",3070 => "00100011",3071 => "11011010",3072 => "11001110",3073 => "01110000",3074 => "01110010",3075 => "01010001",3076 => "10111010",3077 => "00100010",3078 => "10011101",3079 => "11100100",3080 => "11101110",3081 => "00011100",3082 => "11010001",3083 => "11100000",3084 => "00110101",3085 => "00011011",3086 => "11001010",3087 => "10101010",3088 => "01101011",3089 => "00001100",3090 => "10011111",3091 => "00010111",3092 => "11101000",3093 => "11010010",3094 => "01010111",3095 => "00111111",3096 => "00111111",3097 => "10011000",3098 => "00011010",3099 => "10010001",3100 => "01100011",3101 => "00101000",3102 => "10101000",3103 => "00011010",3104 => "11100110",3105 => "11010001",3106 => "01000111",3107 => "11001100",3108 => "01001101",3109 => "10111100",3110 => "00010101",3111 => "00100011",3112 => "10110100",3113 => "01110100",3114 => "01001001",3115 => "01111011",3116 => "11011111",3117 => "11101111",3118 => "10100010",3119 => "01011011",3120 => "10110110",3121 => "01011000",3122 => "01001011",3123 => "10001110",3124 => "11000110",3125 => "10101001",3126 => "11011111",3127 => "00101011",3128 => "10110011",3129 => "01100100",3130 => "01101001",3131 => "11000101",3132 => "11100000",3133 => "00111001",3134 => "00110010",3135 => "00101111",3136 => "00011111",3137 => "00101010",3138 => "01101010",3139 => "01010100",3140 => "11000011",3141 => "11001110",3142 => "01000111",3143 => "01001010",3144 => "11111111",3145 => "10001111",3146 => "01010110",3147 => "01010111",3148 => "10101110",3149 => "00111000",3150 => "00010000",3151 => "00010100",3152 => "00000000",3153 => "01110000",3154 => "10101100",3155 => "00010000",3156 => "10111100",3157 => "00100110",3158 => "11010100",3159 => "11111111",3160 => "01111100",3161 => "10101010",3162 => "10111110",3163 => "00110101",3164 => "10001110",3165 => "01110110",3166 => "01000111",3167 => "10011000",3168 => "11000010",3169 => "00000100",3170 => "00011100",3171 => "00001011",3172 => "01100000",3173 => "11110110",3174 => "11111001",3175 => "11011010",3176 => "00111000",3177 => "00101101",3178 => "10010110",3179 => "00000011",3180 => "01100011",3181 => "11001011",3182 => "10111110",3183 => "11100001",3184 => "01110011",3185 => "00110110",3186 => "01010101",3187 => "11100110",3188 => "01010000",3189 => "10101110",3190 => "01101001",3191 => "10011110",3192 => "10101111",3193 => "11110110",3194 => "00000000",3195 => "00001010",3196 => "01001110",3197 => "00000000",3198 => "11011111",3199 => "10110000",3200 => "01111001",3201 => "10111100",3202 => "10011010",3203 => "00011110",3204 => "01100011",3205 => "00001100",3206 => "10000101",3207 => "11010100",3208 => "10101011",3209 => "11100110",3210 => "00101101",3211 => "10011000",3212 => "00111100",3213 => "01000101",3214 => "11111011",3215 => "10111010",3216 => "10100011",3217 => "10101001",3218 => "00111001",3219 => "01100001",3220 => "11101001",3221 => "11100000",3222 => "01110011",3223 => "10000011",3224 => "11101101",3225 => "01000101",3226 => "11011110",3227 => "00111110",3228 => "11010011",3229 => "11010011",3230 => "01000000",3231 => "11010001",3232 => "00110101",3233 => "01010101",3234 => "11100101",3235 => "01110001",3236 => "00001101",3237 => "00011011",3238 => "10100111",3239 => "01111001",3240 => "01001101",3241 => "01000100",3242 => "01010110",3243 => "00100110",3244 => "01010010",3245 => "01100011",3246 => "01100110",3247 => "10011001",3248 => "01101010",3249 => "11110000",3250 => "11110000",3251 => "00001000",3252 => "01111101",3253 => "10010110",3254 => "10111011",3255 => "11011110",3256 => "01110101",3257 => "11101110",3258 => "01000110",3259 => "01000000",3260 => "01000101",3261 => "11010101",3262 => "00011001",3263 => "11111011",3264 => "00000101",3265 => "00111010",3266 => "01100000",3267 => "11101001",3268 => "10010101",3269 => "01011010",3270 => "00101111",3271 => "11000010",3272 => "01001100",3273 => "11000011",3274 => "11101101",3275 => "01010100",3276 => "11100000",3277 => "01100111",3278 => "11000000",3279 => "01000101",3280 => "00101000",3281 => "10011100",3282 => "11010011",3283 => "01110100",3284 => "10101011",3285 => "10100001",3286 => "00000111",3287 => "01011011",3288 => "01000011",3289 => "11010001",3290 => "11100011",3291 => "10010100",3292 => "01101000",3293 => "10101110",3294 => "10001101",3295 => "01110001",3296 => "00100001",3297 => "10001001",3298 => "10110110",3299 => "10000111",3300 => "11110011",3301 => "01011000",3302 => "01010000",3303 => "10100001",3304 => "01100000",3305 => "11110001",3306 => "01010101",3307 => "01000001",3308 => "00110011",3309 => "00001101",3310 => "01000001",3311 => "11000010",3312 => "00101101",3313 => "11111111",3314 => "10001010",3315 => "10010101",3316 => "11101000",3317 => "00111000",3318 => "01011000",3319 => "01001110",3320 => "01001100",3321 => "01111001",3322 => "01011000",3323 => "11001010",3324 => "00101010",3325 => "10101100",3326 => "11111010",3327 => "11100100",3328 => "11111110",3329 => "10111100",3330 => "00011001",3331 => "10111101",3332 => "00000001",3333 => "01000110",3334 => "01100111",3335 => "01010000",3336 => "00100011",3337 => "10011011",3338 => "00111111",3339 => "11111000",3340 => "00010101",3341 => "10111110",3342 => "01100111",3343 => "00100111",3344 => "11001111",3345 => "10011001",3346 => "00111101",3347 => "01110110",3348 => "11110000",3349 => "11100001",3350 => "10100110",3351 => "10000001",3352 => "01101000",3353 => "10101101",3354 => "00001110",3355 => "00000001",3356 => "10001101",3357 => "10011100",3358 => "01101110",3359 => "00111100",3360 => "01101000",3361 => "10001101",3362 => "00010101",3363 => "01011010",3364 => "10100000",3365 => "01001001",3366 => "01111110",3367 => "00111010",3368 => "10001011",3369 => "01000011",3370 => "11011111",3371 => "10111001",3372 => "10101110",3373 => "01011100",3374 => "10100101",3375 => "00001101",3376 => "00011010",3377 => "10111111",3378 => "00000100",3379 => "11010110",3380 => "10110001",3381 => "00011001",3382 => "01101001",3383 => "10100101",3384 => "01011001",3385 => "00111000",3386 => "10100011",3387 => "01101100",3388 => "10101100",3389 => "00111110",3390 => "10011110",3391 => "01011001",3392 => "11000000",3393 => "11111000",3394 => "10111100",3395 => "01001000",3396 => "10110110",3397 => "00011001",3398 => "10001110",3399 => "11110110",3400 => "10001110",3401 => "01110110",3402 => "01011000",3403 => "10000111",3404 => "01100110",3405 => "01111000",3406 => "00101111",3407 => "10011100",3408 => "01101110",3409 => "01111110",3410 => "01011101",3411 => "00111011",3412 => "10101010",3413 => "10000010",3414 => "00111011",3415 => "00010110",3416 => "11010000",3417 => "00101101",3418 => "00001111",3419 => "01111100",3420 => "00110011",3421 => "00100010",3422 => "10000111",3423 => "10101100",3424 => "01111101",3425 => "11100010",3426 => "10011111",3427 => "01001010",3428 => "01010000",3429 => "01010110",3430 => "10010000",3431 => "11001001",3432 => "01011001",3433 => "01000010",3434 => "10011100",3435 => "00111010",3436 => "10111111",3437 => "10000010",3438 => "10011101",3439 => "11001100",3440 => "10111000",3441 => "10000100",3442 => "00101000",3443 => "01110100",3444 => "01010111",3445 => "00000001",3446 => "01001110",3447 => "10000001",3448 => "11101011",3449 => "00101100",3450 => "10000110",3451 => "11011000",3452 => "01100100",3453 => "00101000",3454 => "10001110",3455 => "10001111",3456 => "00100101",3457 => "10000011",3458 => "10101010",3459 => "10001001",3460 => "10011000",3461 => "00001100",3462 => "10001011",3463 => "10001101",3464 => "10011111",3465 => "10110100",3466 => "10111000",3467 => "10101101",3468 => "01011100",3469 => "11100100",3470 => "10000010",3471 => "11001100",3472 => "01001101",3473 => "11010100",3474 => "10010010",3475 => "01110100",3476 => "00010011",3477 => "00011010",3478 => "11110101",3479 => "11100001",3480 => "00111101",3481 => "01001100",3482 => "10011011",3483 => "01100000",3484 => "10110010",3485 => "01101110",3486 => "10110000",3487 => "10110000",3488 => "11000001",3489 => "00010101",3490 => "00001101",3491 => "00100110",3492 => "10001110",3493 => "00011111",3494 => "11101100",3495 => "01001101",3496 => "10100100",3497 => "01111111",3498 => "10000010",3499 => "11001110",3500 => "11000001",3501 => "00110101",3502 => "10100111",3503 => "11110101",3504 => "00010000",3505 => "00010101",3506 => "01111010",3507 => "11110100",3508 => "10100010",3509 => "10000110",3510 => "01001000",3511 => "01001001",3512 => "11001111",3513 => "00111111",3514 => "01010000",3515 => "11110011",3516 => "01001000",3517 => "00001110",3518 => "00101110",3519 => "01101000",3520 => "10110001",3521 => "10011110",3522 => "01100001",3523 => "01101111",3524 => "00111001",3525 => "00101001",3526 => "01011100",3527 => "10111111",3528 => "00001101",3529 => "01111011",3530 => "01010001",3531 => "01011111",3532 => "10000111",3533 => "00100100",3534 => "01111110",3535 => "10111011",3536 => "00100010",3537 => "01110111",3538 => "00110111",3539 => "11010010",3540 => "10111010",3541 => "00110100",3542 => "00000011",3543 => "01101100",3544 => "11101111",3545 => "01011110",3546 => "01011001",3547 => "01001101",3548 => "11110000",3549 => "11101110",3550 => "00110011",3551 => "10100100",3552 => "11100011",3553 => "10000010",3554 => "01101101",3555 => "01010000",3556 => "10100010",3557 => "10101010",3558 => "01111011",3559 => "01110111",3560 => "00000110",3561 => "11111100",3562 => "00010100",3563 => "11111000",3564 => "11001010",3565 => "11101010",3566 => "11000000",3567 => "00111111",3568 => "01001110",3569 => "10100011",3570 => "10110001",3571 => "10011111",3572 => "00001110",3573 => "11001001",3574 => "01101010",3575 => "01001010",3576 => "01000101",3577 => "01000001",3578 => "00011001",3579 => "10011100",3580 => "10010111",3581 => "11100001",3582 => "00001001",3583 => "01101000",3584 => "10101010",3585 => "00011110",3586 => "01111001",3587 => "01010001",3588 => "11010000",3589 => "10011011",3590 => "11110100",3591 => "00010010",3592 => "01111001",3593 => "01010111",3594 => "11101111",3595 => "00000011",3596 => "10010000",3597 => "01110100",3598 => "11000010",3599 => "10110001",3600 => "01010000",3601 => "01001100",3602 => "11101101",3603 => "10001000",3604 => "10010100",3605 => "11000010",3606 => "11100101",3607 => "11001011",3608 => "01110011",3609 => "01110000",3610 => "00101010",3611 => "01001110",3612 => "01100111",3613 => "01010001",3614 => "11111111",3615 => "01111100",3616 => "01111111",3617 => "00111111",3618 => "11010111",3619 => "00101111",3620 => "10011011",3621 => "01101111",3622 => "00001000",3623 => "00111000",3624 => "01000011",3625 => "11010111",3626 => "00000110",3627 => "11011101",3628 => "00100010",3629 => "11011000",3630 => "01100001",3631 => "10111000",3632 => "01010011",3633 => "00100101",3634 => "01100010",3635 => "11100110",3636 => "00100010",3637 => "01110111",3638 => "01111110",3639 => "10100000",3640 => "01010011",3641 => "00000011",3642 => "10001100",3643 => "10010011",3644 => "11111011",3645 => "10110111",3646 => "00011100",3647 => "11100101",3648 => "11010001",3649 => "11000010",3650 => "10000000",3651 => "00111011",3652 => "00101110",3653 => "00101110",3654 => "10010101",3655 => "01010111",3656 => "10101010",3657 => "11110011",3658 => "01101001",3659 => "00101011",3660 => "00010010",3661 => "01010001",3662 => "00011111",3663 => "10010011",3664 => "00111111",3665 => "11101100",3666 => "10010011",3667 => "01101000",3668 => "11000011",3669 => "00010000",3670 => "11110111",3671 => "00110110",3672 => "10011101",3673 => "10001110",3674 => "01001000",3675 => "01110110",3676 => "11100100",3677 => "00110000",3678 => "01111111",3679 => "01101100",3680 => "10100001",3681 => "10011010",3682 => "01001101",3683 => "10001011",3684 => "01011000",3685 => "00010010",3686 => "00100101",3687 => "11100001",3688 => "00100110",3689 => "10101100",3690 => "01011001",3691 => "10101110",3692 => "00011101",3693 => "10001110",3694 => "01111000",3695 => "00011011",3696 => "01110111",3697 => "11110101",3698 => "00001010",3699 => "10111001",3700 => "01011001",3701 => "11110101",3702 => "01101010",3703 => "11010011",3704 => "01100010",3705 => "11001100",3706 => "11010000",3707 => "00101101",3708 => "11011011",3709 => "10100010",3710 => "00001100",3711 => "01100101",3712 => "01000110",3713 => "01110000",3714 => "10100000",3715 => "11010110",3716 => "10101111",3717 => "11001000",3718 => "10110011",3719 => "10111010",3720 => "01010100",3721 => "11010110",3722 => "11000100",3723 => "00010101",3724 => "00111111",3725 => "01010010",3726 => "00101111",3727 => "10110100",3728 => "10011111",3729 => "10111010",3730 => "01100011",3731 => "01011101",3732 => "01001100",3733 => "11101100",3734 => "01011000",3735 => "01111001",3736 => "11001100",3737 => "00010011",3738 => "10001110",3739 => "11101000",3740 => "10110000",3741 => "01110101",3742 => "10011010",3743 => "11010011",3744 => "00100111",3745 => "10011101",3746 => "10000100",3747 => "11100001",3748 => "01111100",3749 => "01110110",3750 => "00010101",3751 => "10011101",3752 => "10110010",3753 => "10010101",3754 => "01110101",3755 => "10000101",3756 => "10111110",3757 => "00010010",3758 => "01001010",3759 => "10011111",3760 => "01011110",3761 => "11001000",3762 => "11111100",3763 => "00101110",3764 => "00101011",3765 => "10101001",3766 => "01000101",3767 => "11010011",3768 => "11101000",3769 => "01000000",3770 => "00010000",3771 => "01110110",3772 => "01111011",3773 => "10010011",3774 => "00000110",3775 => "00001100",3776 => "11010101",3777 => "01111100",3778 => "01011000",3779 => "01000101",3780 => "01000001",3781 => "01000101",3782 => "10100100",3783 => "10100101",3784 => "00110010",3785 => "01110111",3786 => "11110001",3787 => "10110010",3788 => "10011011",3789 => "10111000",3790 => "11010100",3791 => "00111100",3792 => "10010011",3793 => "01010101",3794 => "00101001",3795 => "11000110",3796 => "10011111",3797 => "01011101",3798 => "11011000",3799 => "11100001",3800 => "10010101",3801 => "00000011",3802 => "00011010",3803 => "10010111",3804 => "01101000",3805 => "01000110",3806 => "10101101",3807 => "01111100",3808 => "11011001",3809 => "01101000",3810 => "10110001",3811 => "11111100",3812 => "00010011",3813 => "11001000",3814 => "10111101",3815 => "11000001",3816 => "10110110",3817 => "00011000",3818 => "01001001",3819 => "10100101",3820 => "00100011",3821 => "00011011",3822 => "00111110",3823 => "11101110",3824 => "00011001",3825 => "10001011",3826 => "00101011",3827 => "01000001",3828 => "01101111",3829 => "00110111",3830 => "11110001",3831 => "10001110",3832 => "10010100",3833 => "01000101",3834 => "01000100",3835 => "10110111",3836 => "01011101",3837 => "10111010",3838 => "11000010",3839 => "01111101",3840 => "11000001",3841 => "01111100",3842 => "10100011",3843 => "01110000",3844 => "01001001",3845 => "11011100",3846 => "11000111",3847 => "11010011",3848 => "00101011",3849 => "10110001",3850 => "01101001",3851 => "10111010",3852 => "01101010",3853 => "01100101",3854 => "11100101",3855 => "10111001",3856 => "11001110",3857 => "11100001",3858 => "10000010",3859 => "11100000",3860 => "10000111",3861 => "10011101",3862 => "01000000",3863 => "01000111",3864 => "01111011",3865 => "11011110",3866 => "00111101",3867 => "11110100",3868 => "00111010",3869 => "00011011",3870 => "11110000",3871 => "01010111",3872 => "00001100",3873 => "10110110",3874 => "11011100",3875 => "11111001",3876 => "10101011",3877 => "11000000",3878 => "11101101",3879 => "10110111",3880 => "01101010",3881 => "01100010",3882 => "01001000",3883 => "01101000",3884 => "10110111",3885 => "01010010",3886 => "00100001",3887 => "10111011",3888 => "00010110",3889 => "01110100",3890 => "01101101",3891 => "11101101",3892 => "00001011",3893 => "00000111",3894 => "10111000",3895 => "10010110",3896 => "10101010",3897 => "11000101",3898 => "10110101",3899 => "00110000",3900 => "00110010",3901 => "01000001",3902 => "01111100",3903 => "10001011",3904 => "10100011",3905 => "01110000",3906 => "01000011",3907 => "01101100",3908 => "01000101",3909 => "10000101",3910 => "00000010",3911 => "00101110",3912 => "00101001",3913 => "00001111",3914 => "11110001",3915 => "01001110",3916 => "01001110",3917 => "11001101",3918 => "10000011",3919 => "11010000",3920 => "10101000",3921 => "01010110",3922 => "00001110",3923 => "10111000",3924 => "10100110",3925 => "00000110",3926 => "00001101",3927 => "11011111",3928 => "11001100",3929 => "11101000",3930 => "01111110",3931 => "10001001",3932 => "01101100",3933 => "10000011",3934 => "10001011",3935 => "00101000",3936 => "01000001",3937 => "11011001",3938 => "01001011",3939 => "10101110",3940 => "10000111",3941 => "10001100",3942 => "10110000",3943 => "00010001",3944 => "00111101",3945 => "00110000",3946 => "01111000",3947 => "11110011",3948 => "10101111",3949 => "11011001",3950 => "01100110",3951 => "10110000",3952 => "00111100",3953 => "00010101",3954 => "11101000",3955 => "01001010",3956 => "01010111",3957 => "01001101",3958 => "00110010",3959 => "11101101",3960 => "01001001",3961 => "10011100",3962 => "01101111",3963 => "00110001",3964 => "01110001",3965 => "10011000",3966 => "00100110",3967 => "10000001",3968 => "01001100",3969 => "11101100",3970 => "11101101",3971 => "11001010",3972 => "00001101",3973 => "00110110",3974 => "11110100",3975 => "01001000",3976 => "01101111",3977 => "00010101",3978 => "00010010",3979 => "00001010",3980 => "01101011",3981 => "01101011",3982 => "11110000",3983 => "10110110",3984 => "11001011",3985 => "11011001",3986 => "11110000",3987 => "11110101",3988 => "10110011",3989 => "10000110",3990 => "01011011",3991 => "01010101",3992 => "01000100",3993 => "01110010",3994 => "01011001",3995 => "10110001",3996 => "10000010",3997 => "00101000",3998 => "11111011",3999 => "10000011",4000 => "11011011",4001 => "10111001",4002 => "00101110",4003 => "00010100",4004 => "00100001",4005 => "10110001",4006 => "00110010",4007 => "11000111",4008 => "11111001",4009 => "00100010",4010 => "00110100",4011 => "10011000",4012 => "11010101",4013 => "10011010",4014 => "11001011",4015 => "11000100",4016 => "01100101",4017 => "11111110",4018 => "00101101",4019 => "00000001",4020 => "11000110",4021 => "00000100",4022 => "11100011",4023 => "10101100",4024 => "00010010",4025 => "01101100",4026 => "01110101",4027 => "11001011",4028 => "01011001",4029 => "01110001",4030 => "11010000",4031 => "01100011",4032 => "01001001",4033 => "00111000",4034 => "10011101",4035 => "10010010",4036 => "01011111",4037 => "00101110",4038 => "10000111",4039 => "01011111",4040 => "11011010",4041 => "00100111",4042 => "00000101",4043 => "11100111",4044 => "11111011",4045 => "10010001",4046 => "10100101",4047 => "10100101",4048 => "00110011",4049 => "01100010",4050 => "00110110",4051 => "00110000",4052 => "01100000",4053 => "01000111",4054 => "01100010",4055 => "11001001",4056 => "10011101",4057 => "11100110",4058 => "00110011",4059 => "11110101",4060 => "11000101",4061 => "01101111",4062 => "01110101",4063 => "01000111",4064 => "01100011",4065 => "11110000",4066 => "11001011",4067 => "10000111",4068 => "11100101",4069 => "11010011",4070 => "00110010",4071 => "11111001",4072 => "10001001",4073 => "10101001",4074 => "11000001",4075 => "11011110",4076 => "10111010",4077 => "01000000",4078 => "00110100",4079 => "10101010",4080 => "00011110",4081 => "10111110",4082 => "00011101",4083 => "10101001",4084 => "00010011",4085 => "00000001",4086 => "10111101",4087 => "10101101",4088 => "11110010",4089 => "00100001",4090 => "11001000",4091 => "01011100",4092 => "01000111",4093 => "10010010",4094 => "00110010",4095 => "10110111",4096 => "01010010",4097 => "00011000",4098 => "00010010",4099 => "10110000",4100 => "10100111",4101 => "10110111",4102 => "11001001",4103 => "10010001",4104 => "10001011",4105 => "10101001",4106 => "00110100",4107 => "11100110",4108 => "11000010",4109 => "10001000",4110 => "00010000",4111 => "01100000",4112 => "11100100",4113 => "11001010",4114 => "01011011",4115 => "11111001",4116 => "01101101",4117 => "00110001",4118 => "00101110",4119 => "10001001",4120 => "11111010",4121 => "00011001",4122 => "11000101",4123 => "10110010",4124 => "01000000",4125 => "11110001",4126 => "00011100",4127 => "10100100",4128 => "11010011",4129 => "01010010",4130 => "00001110",4131 => "01000010",4132 => "01011111",4133 => "00111001",4134 => "01111001",4135 => "11110100",4136 => "01010011",4137 => "00100011",4138 => "01111011",4139 => "00011111",4140 => "10111110",4141 => "11011001",4142 => "00100101",4143 => "00101100",4144 => "01011011",4145 => "10110010",4146 => "00110101",4147 => "10110010",4148 => "01001100",4149 => "01011101",4150 => "11100000",4151 => "00110000",4152 => "10011000",4153 => "00010010",4154 => "10001101",4155 => "01111111",4156 => "00011001",4157 => "01111001",4158 => "10110000",4159 => "11000010",4160 => "00001001",4161 => "10011110",4162 => "00011011",4163 => "00100100",4164 => "10001111",4165 => "00111101",4166 => "10011001",4167 => "10001111",4168 => "10011100",4169 => "11111011",4170 => "01010111",4171 => "11101110",4172 => "00001101",4173 => "01000100",4174 => "01100110",4175 => "10100011",4176 => "10011100",4177 => "11110000",4178 => "01000010",4179 => "00101111",4180 => "00110011",4181 => "10100010",4182 => "01001001",4183 => "01101010",4184 => "11110001",4185 => "11101000",4186 => "10111110",4187 => "00110111",4188 => "11001010",4189 => "11010100",4190 => "01110001",4191 => "11011111",4192 => "11001010",4193 => "10110111",4194 => "11010000",4195 => "01110111",4196 => "10011011",4197 => "01111011",4198 => "01101010",4199 => "10000110",4200 => "11100111",4201 => "00011100",4202 => "00010000",4203 => "10011011",4204 => "10001010",4205 => "00011000",4206 => "10110111",4207 => "11111011",4208 => "00010010",4209 => "01101101",4210 => "01001001",4211 => "11111011",4212 => "00001101",4213 => "00100100",4214 => "11111011",4215 => "10101101",4216 => "11110011",4217 => "00101101",4218 => "01100011",4219 => "11100100",4220 => "11100010",4221 => "01110110",4222 => "10101000",4223 => "01000000",4224 => "01110110",4225 => "10111011",4226 => "10111001",4227 => "11101100",4228 => "11100011",4229 => "10000100",4230 => "01101010",4231 => "11100111",4232 => "00101111",4233 => "00100010",4234 => "10010010",4235 => "10011100",4236 => "00000100",4237 => "10001000",4238 => "10100100",4239 => "01011110",4240 => "11011000",4241 => "11111101",4242 => "11001011",4243 => "10000100",4244 => "11000001",4245 => "00101000",4246 => "00001111",4247 => "01101000",4248 => "10101001",4249 => "00100000",4250 => "01100100",4251 => "10001101",4252 => "01111111",4253 => "00010110",4254 => "01010110",4255 => "11011100",4256 => "00110011",4257 => "11111111",4258 => "00001110",4259 => "00101110",4260 => "10111001",4261 => "11010111",4262 => "10111000",4263 => "01011010",4264 => "01111111",4265 => "11100101",4266 => "00000101",4267 => "00101110",4268 => "11010111",4269 => "00110110",4270 => "01111011",4271 => "10001100",4272 => "01110100",4273 => "10101101",4274 => "01110001",4275 => "11001111",4276 => "00011101",4277 => "01100110",4278 => "01010000",4279 => "11101010",4280 => "11101101",4281 => "11111010",4282 => "11110001",4283 => "00100100",4284 => "10100011",4285 => "10010011",4286 => "01111001",4287 => "11000101",4288 => "10110101",4289 => "00010101",4290 => "01001010",4291 => "11110110",4292 => "01001011",4293 => "11100011",4294 => "10110010",4295 => "11100000",4296 => "11100100",4297 => "01000101",4298 => "10101010",4299 => "10000010",4300 => "01111001",4301 => "10111101",4302 => "11110001",4303 => "10101111",4304 => "11111101",4305 => "10011111",4306 => "00000010",4307 => "01011110",4308 => "10111100",4309 => "11100011",4310 => "10111010",4311 => "01111011",4312 => "10101101",4313 => "00000011",4314 => "11110001",4315 => "11110001",4316 => "11111011",4317 => "10010111",4318 => "00011100",4319 => "01100000",4320 => "11111101",4321 => "01101011",4322 => "00001001",4323 => "11001001",4324 => "10111110",4325 => "10000010",4326 => "11001001",4327 => "10110001",4328 => "01011010",4329 => "10111100",4330 => "10000110",4331 => "10100001",4332 => "10011010",4333 => "00001000",4334 => "01101011",4335 => "10011000",4336 => "01110011",4337 => "00010111",4338 => "00111000",4339 => "00110111",4340 => "01110000",4341 => "01001111",4342 => "11111110",4343 => "01011100",4344 => "01010100",4345 => "01011100",4346 => "11010000",4347 => "00110111",4348 => "11010001",4349 => "00010101",4350 => "10001111",4351 => "11101110",4352 => "11000011",4353 => "00110110",4354 => "11010111",4355 => "00000010",4356 => "00100001",4357 => "10101010",4358 => "11011001",4359 => "11010010",4360 => "11011001",4361 => "11010011",4362 => "00101001",4363 => "01001110",4364 => "01110001",4365 => "00001100",4366 => "11010001",4367 => "11001100",4368 => "01010000",4369 => "01100101",4370 => "10111101",4371 => "01111010",4372 => "11111101",4373 => "01100101",4374 => "10010011",4375 => "10010001",4376 => "10010110",4377 => "11001110",4378 => "10010001",4379 => "00010100",4380 => "01001010",4381 => "01011000",4382 => "10101101",4383 => "10000111",4384 => "01100111",4385 => "01101100",4386 => "10101101",4387 => "10110111",4388 => "01010011",4389 => "00110111",4390 => "01000010",4391 => "11011100",4392 => "11000111",4393 => "01110011",4394 => "10101111",4395 => "01000111",4396 => "10100001",4397 => "10011011",4398 => "11110001",4399 => "01001010",4400 => "10011101",4401 => "00110110",4402 => "00010001",4403 => "11000110",4404 => "10110101",4405 => "00000001",4406 => "11100011",4407 => "01011001",4408 => "11001110",4409 => "10001011",4410 => "10100011",4411 => "00010101",4412 => "00010010",4413 => "10000001",4414 => "00101100",4415 => "00101000",4416 => "00011000",4417 => "10011110",4418 => "10010110",4419 => "00111111",4420 => "00000111",4421 => "11110001",4422 => "00001001",4423 => "10010010",4424 => "10011110",4425 => "11101110",4426 => "10001001",4427 => "10011101",4428 => "01010110",4429 => "11010110",4430 => "01110000",4431 => "11001110",4432 => "11001000",4433 => "00010101",4434 => "00011010",4435 => "11110011",4436 => "00111001",4437 => "00011101",4438 => "00110111",4439 => "01011110",4440 => "01000100",4441 => "01101111",4442 => "00010100",4443 => "00110001",4444 => "01111001",4445 => "10100110",4446 => "01001001",4447 => "00001110",4448 => "01010010",4449 => "11111101",4450 => "11010010",4451 => "11100110",4452 => "11100101",4453 => "00110010",4454 => "10000001",4455 => "11001110",4456 => "10010011",4457 => "00001001",4458 => "00011110",4459 => "10111000",4460 => "00011011",4461 => "11011110",4462 => "10000010",4463 => "11011101",4464 => "10000100",4465 => "01100111",4466 => "01110010",4467 => "10110011",4468 => "00100100",4469 => "10000110",4470 => "00100011",4471 => "01010101",4472 => "10110010",4473 => "01101101",4474 => "11001010",4475 => "10001011",4476 => "01100111",4477 => "11110101",4478 => "01010011",4479 => "10011101",4480 => "01101100",4481 => "01001111",4482 => "01001000",4483 => "01111011",4484 => "01110011",4485 => "00011110",4486 => "00000110",4487 => "00001110",4488 => "10000101",4489 => "00110111",4490 => "01001101",4491 => "11000111",4492 => "11011001",4493 => "00111101",4494 => "10111101",4495 => "00100111",4496 => "00101000",4497 => "01111100",4498 => "01001110",4499 => "11101011",4500 => "00101010",4501 => "00111101",4502 => "10110110",4503 => "11010110",4504 => "11100001",4505 => "11011001",4506 => "11011010",4507 => "01110001",4508 => "01000111",4509 => "00100111",4510 => "11000110",4511 => "11101001",4512 => "11111011",4513 => "00001001",4514 => "00111010",4515 => "10100101",4516 => "00100001",4517 => "10111100",4518 => "01110001",4519 => "00101101",4520 => "10101011",4521 => "01100111",4522 => "11101001",4523 => "01000010",4524 => "10000111",4525 => "01001000",4526 => "00011000",4527 => "10011010",4528 => "11100010",4529 => "01010011",4530 => "11111011",4531 => "11010101",4532 => "10111001",4533 => "00101110",4534 => "01100011",4535 => "10000110",4536 => "10101100",4537 => "11111110",4538 => "00100101",4539 => "10111101",4540 => "11010011",4541 => "11010010",4542 => "11110001",4543 => "00100000",4544 => "11110101",4545 => "01011011",4546 => "11111101",4547 => "00010100",4548 => "01010111",4549 => "11101110",4550 => "00101011",4551 => "01100111",4552 => "10111100",4553 => "11000010",4554 => "00111111",4555 => "01011100",4556 => "00011011",4557 => "10000010",4558 => "00000001",4559 => "11111111",4560 => "01001010",4561 => "11110100",4562 => "01110000",4563 => "11100000",4564 => "00000001",4565 => "00010011",4566 => "10110100",4567 => "01110100",4568 => "00011110",4569 => "00010010",4570 => "01100011",4571 => "11001011",4572 => "10111011",4573 => "11101001",4574 => "10001100",4575 => "11101010",4576 => "10001011",4577 => "01010101",4578 => "00010111",4579 => "10110110",4580 => "01101001",4581 => "11011000",4582 => "00100111",4583 => "00011110",4584 => "00011011",4585 => "10111000",4586 => "10110100",4587 => "01101101",4588 => "01011101",4589 => "00101011",4590 => "01000011",4591 => "00100101",4592 => "10100111",4593 => "10111001",4594 => "10011101",4595 => "00111010",4596 => "11110000",4597 => "00001111",4598 => "11000100",4599 => "10001101",4600 => "01001010",4601 => "00101011",4602 => "11001011",4603 => "10110101",4604 => "11001111",4605 => "11111101",4606 => "00000000",4607 => "01011110",4608 => "10011110",4609 => "01110100",4610 => "11011100",4611 => "00111101",4612 => "11110101",4613 => "00100011",4614 => "00101001",4615 => "00101100",4616 => "01110010",4617 => "00001000",4618 => "11111101",4619 => "01000010",4620 => "00101100",4621 => "01101111",4622 => "11011110",4623 => "10100011",4624 => "10001011",4625 => "10111111",4626 => "00111000",4627 => "11111011",4628 => "10100111",4629 => "01101000",4630 => "00010011",4631 => "11011101",4632 => "00100001",4633 => "01010001",4634 => "01011110",4635 => "00010100",4636 => "01110100",4637 => "10010000",4638 => "11010011",4639 => "00100101",4640 => "01010011",4641 => "00100011",4642 => "00010000",4643 => "01100001",4644 => "01101011",4645 => "01011001",4646 => "10111101",4647 => "11111000",4648 => "11111010",4649 => "00111101",4650 => "01111110",4651 => "11110111",4652 => "01011101",4653 => "11010011",4654 => "01010101",4655 => "10110010",4656 => "00010100",4657 => "01000100",4658 => "10000000",4659 => "01001110",4660 => "10001100",4661 => "00100111",4662 => "11000110",4663 => "01010101",4664 => "01101001",4665 => "10000000",4666 => "00111111",4667 => "10110100",4668 => "00001011",4669 => "10101000",4670 => "00011100",4671 => "10011101",4672 => "10111000",4673 => "11010110",4674 => "00110001",4675 => "10111101",4676 => "00100011",4677 => "00100100",4678 => "01001010",4679 => "10111100",4680 => "00100111",4681 => "00100100",4682 => "10000000",4683 => "01100101",4684 => "01011000",4685 => "11001101",4686 => "10001000",4687 => "10011011",4688 => "01010001",4689 => "00110110",4690 => "11100101",4691 => "11001011",4692 => "10010000",4693 => "01000110",4694 => "00111100",4695 => "10110000",4696 => "11111010",4697 => "10010100",4698 => "11011110",4699 => "00010100",4700 => "10111010",4701 => "00001010",4702 => "01010111",4703 => "00000100",4704 => "10011011",4705 => "11001000",4706 => "00100111",4707 => "00001100",4708 => "11110000",4709 => "10101110",4710 => "11101101",4711 => "01111000",4712 => "00111010",4713 => "01001100",4714 => "01010100",4715 => "11110101",4716 => "01111110",4717 => "01110111",4718 => "10011011",4719 => "01110010",4720 => "10010000",4721 => "01010111",4722 => "10110001",4723 => "11111101",4724 => "11000101",4725 => "10011110",4726 => "00010000",4727 => "00111011",4728 => "11101101",4729 => "00101010",4730 => "10101000",4731 => "10010110",4732 => "11000111",4733 => "00010101",4734 => "11100000",4735 => "01010000",4736 => "11000110",4737 => "01000001",4738 => "11011001",4739 => "00000011",4740 => "10101100",4741 => "01111011",4742 => "00011111",4743 => "10010101",4744 => "00110101",4745 => "11110110",4746 => "11000011",4747 => "11101100",4748 => "01010001",4749 => "10011101",4750 => "00110000",4751 => "00011001",4752 => "01010100",4753 => "00000000",4754 => "11110001",4755 => "10110000",4756 => "00101001",4757 => "10010110",4758 => "00100001",4759 => "00110010",4760 => "10101000",4761 => "00101000",4762 => "10011011",4763 => "00111100",4764 => "01011100",4765 => "10001011",4766 => "01011111",4767 => "00010111",4768 => "01110000",4769 => "11101110",4770 => "01001011",4771 => "10111011",4772 => "11101011",4773 => "00010010",4774 => "11110101",4775 => "11110101",4776 => "01100010",4777 => "00011100",4778 => "00011001",4779 => "01001101",4780 => "01001011",4781 => "00100101",4782 => "10101111",4783 => "01101101",4784 => "01111000",4785 => "00010001",4786 => "11000010",4787 => "11001111",4788 => "10111111",4789 => "10001110",4790 => "01110011",4791 => "11101001",4792 => "01101010",4793 => "10101111",4794 => "00100111",4795 => "01110111",4796 => "11100001",4797 => "01111011",4798 => "00111010",4799 => "00001001",4800 => "11011001",4801 => "01000001",4802 => "11110100",4803 => "00000111",4804 => "10110101",4805 => "10010001",4806 => "01100011",4807 => "11100000",4808 => "01010010",4809 => "11100010",4810 => "10100111",4811 => "01101000",4812 => "01101010",4813 => "01011101",4814 => "00101100",4815 => "01111111",4816 => "11000001",4817 => "00010001",4818 => "01100110",4819 => "11001000",4820 => "01010011",4821 => "01100100",4822 => "11110111",4823 => "00001111",4824 => "00100011",4825 => "10110111",4826 => "00110000",4827 => "10011111",4828 => "01110101",4829 => "00010111",4830 => "11000001",4831 => "01100100",4832 => "01011010",4833 => "11101010",4834 => "11110011",4835 => "10110001",4836 => "00101100",4837 => "10100000",4838 => "00001000",4839 => "00000001",4840 => "10011111",4841 => "10010110",4842 => "01101101",4843 => "11000010",4844 => "11001000",4845 => "11100010",4846 => "00110100",4847 => "01100001",4848 => "10100100",4849 => "10001110",4850 => "00011011",4851 => "10011011",4852 => "01100000",4853 => "00011001",4854 => "00011111",4855 => "10111110",4856 => "10110011",4857 => "00001101",4858 => "10111000",4859 => "00011111",4860 => "01101100",4861 => "00100111",4862 => "10110011",4863 => "10000100",4864 => "11111000",4865 => "01011011",4866 => "01101110",4867 => "00111010",4868 => "01000101",4869 => "01010110",4870 => "11000011",4871 => "10100101",4872 => "01100000",4873 => "01010000",4874 => "01011100",4875 => "10101010",4876 => "10011001",4877 => "01100001",4878 => "10000001",4879 => "01100010",4880 => "01101101",4881 => "11011111",4882 => "00110111",4883 => "11110111",4884 => "10100101",4885 => "11100000",4886 => "00100100",4887 => "11011101",4888 => "00011100",4889 => "11011100",4890 => "00001011",4891 => "00000101",4892 => "01101101",4893 => "10011111",4894 => "11010110",4895 => "11110110",4896 => "01001111",4897 => "11110110",4898 => "10101100",4899 => "01010100",4900 => "01111111",4901 => "11101101",4902 => "11000011",4903 => "11101110",4904 => "11010001",4905 => "00010101",4906 => "10011011",4907 => "11000100",4908 => "00001010",4909 => "10100000",4910 => "11100000",4911 => "01100001",4912 => "11011010",4913 => "11100111",4914 => "01010010",4915 => "10001010",4916 => "00101111",4917 => "01010100",4918 => "10111001",4919 => "10111000",4920 => "01010010",4921 => "10111011",4922 => "00001111",4923 => "10000111",4924 => "00010101",4925 => "00110100",4926 => "01011111",4927 => "01110000",4928 => "01001010",4929 => "01101000",4930 => "11100000",4931 => "11111110",4932 => "10000111",4933 => "00000110",4934 => "00011100",4935 => "00000111",4936 => "01111111",4937 => "01011001",4938 => "11001011",4939 => "01100100",4940 => "01010111",4941 => "11100111",4942 => "11011010",4943 => "00000011",4944 => "01000011",4945 => "01010011",4946 => "10111100",4947 => "11110110",4948 => "01010100",4949 => "10010010",4950 => "10111001",4951 => "01100001",4952 => "10011000",4953 => "01001001",4954 => "00000001",4955 => "11100111",4956 => "01000101",4957 => "11000101",4958 => "01011001",4959 => "01101000",4960 => "01000101",4961 => "11110101",4962 => "10110010",4963 => "11000000",4964 => "00011100",4965 => "01010000",4966 => "10010101",4967 => "01110100",4968 => "11100110",4969 => "11010000",4970 => "10011100",4971 => "01101111",4972 => "01101100",4973 => "11100100",4974 => "10111111",4975 => "10110011",4976 => "01000011",4977 => "11111100",4978 => "11111111",4979 => "01101001",4980 => "01101100",4981 => "10010000",4982 => "01110100",4983 => "10010101",4984 => "00110011",4985 => "11110011",4986 => "00110010",4987 => "10110110",4988 => "00001001",4989 => "01010011",4990 => "10111111",4991 => "00001101",4992 => "00000110",4993 => "01110110",4994 => "01010001",4995 => "01110011",4996 => "01100101",4997 => "10110000",4998 => "11110100",4999 => "00000111",5000 => "10011010",5001 => "00111110",5002 => "11011010",5003 => "11010010",5004 => "00000110",5005 => "00000001",5006 => "11100000",5007 => "10010100",5008 => "01101011",5009 => "10011010",5010 => "11111010",5011 => "10101111",5012 => "11100110",5013 => "01101001",5014 => "11010101",5015 => "10001111",5016 => "01100101",5017 => "11011101",5018 => "01101111",5019 => "00110010",5020 => "10000110",5021 => "01001100",5022 => "10011011",5023 => "11010110",5024 => "10001111",5025 => "01111111",5026 => "00010001",5027 => "10000000",5028 => "11000010",5029 => "10111001",5030 => "11110001",5031 => "00000101",5032 => "00110100",5033 => "11011011",5034 => "01000100",5035 => "11010001",5036 => "01101111",5037 => "11101111",5038 => "01100010",5039 => "01101001",5040 => "01001110",5041 => "11010001",5042 => "10110000",5043 => "00111011",5044 => "10011111",5045 => "10011010",5046 => "11100101",5047 => "10100100",5048 => "01010100",5049 => "00011010",5050 => "10100110",5051 => "00000100",5052 => "10101101",5053 => "11111000",5054 => "00011011",5055 => "00011101",5056 => "00000000",5057 => "01111000",5058 => "00101000",5059 => "11110001",5060 => "00111000",5061 => "01110011",5062 => "10001100",5063 => "10011010",5064 => "00010100",5065 => "01001110",5066 => "10010010",5067 => "00101010",5068 => "01100010",5069 => "11110001",5070 => "01000010",5071 => "00100000",5072 => "10100011",5073 => "00110100",5074 => "11101100",5075 => "10000010",5076 => "10100111",5077 => "01111011",5078 => "10110000",5079 => "00100101",5080 => "00110110",5081 => "00000011",5082 => "00101100",5083 => "01100110",5084 => "00011011",5085 => "11110010",5086 => "01111111",5087 => "01011000",5088 => "01100110",5089 => "01001000",5090 => "00101110",5091 => "01101111",5092 => "01110101",5093 => "01101011",5094 => "00010010",5095 => "01000000",5096 => "01101110",5097 => "10000100",5098 => "01011101",5099 => "01101100",5100 => "00010100",5101 => "10001110",5102 => "10101010",5103 => "10100010",5104 => "11011110",5105 => "00111001",5106 => "01000001",5107 => "10110001",5108 => "00111010",5109 => "01001000",5110 => "01111011",5111 => "10011111",5112 => "01100100",5113 => "10011011",5114 => "01101100",5115 => "10101110",5116 => "10001011",5117 => "11000011",5118 => "00101001",5119 => "00111010",5120 => "11001001",5121 => "10111110",5122 => "00100000",5123 => "11001000",5124 => "10000100",5125 => "00110001",5126 => "11100011",5127 => "01111111",5128 => "11101000",5129 => "01000110",5130 => "00000110",5131 => "01111100",5132 => "10101111",5133 => "11110110",5134 => "01100100",5135 => "01101010",5136 => "11101001",5137 => "11000011",5138 => "10000000",5139 => "10110110",5140 => "10101111",5141 => "11110010",5142 => "00010100",5143 => "01110011",5144 => "01001111",5145 => "01011010",5146 => "01101000",5147 => "11001010",5148 => "01100000",5149 => "10001000",5150 => "11110001",5151 => "10110000",5152 => "00100101",5153 => "10010000",5154 => "10101010",5155 => "10101010",5156 => "01010110",5157 => "01100011",5158 => "00110001",5159 => "01110111",5160 => "01100011",5161 => "10001011",5162 => "01110001",5163 => "11100101",5164 => "11100110",5165 => "00000101",5166 => "11110001",5167 => "00111100",5168 => "01000011",5169 => "11001011",5170 => "11110000",5171 => "01101000",5172 => "01100010",5173 => "01111110",5174 => "11101110",5175 => "01100001",5176 => "11000000",5177 => "10001101",5178 => "11110000",5179 => "11100101",5180 => "11011100",5181 => "10011011",5182 => "11101101",5183 => "10111010",5184 => "11100101",5185 => "11010011",5186 => "01001101",5187 => "00011010",5188 => "01111000",5189 => "00001011",5190 => "10110010",5191 => "01101011",5192 => "01000000",5193 => "01110101",5194 => "11000011",5195 => "11111111",5196 => "10011011",5197 => "00111000",5198 => "10011111",5199 => "11010101",5200 => "10000011",5201 => "10011011",5202 => "00011000",5203 => "11001111",5204 => "10000011",5205 => "11100011",5206 => "01011000",5207 => "00101010",5208 => "01011001",5209 => "00100001",5210 => "00001011",5211 => "10111100",5212 => "11100001",5213 => "00101010",5214 => "01111001",5215 => "00111100",5216 => "01010110",5217 => "10101000",5218 => "10010010",5219 => "00100001",5220 => "01110010",5221 => "00010001",5222 => "11001101",5223 => "11110100",5224 => "01101101",5225 => "00110101",5226 => "01111011",5227 => "10001101",5228 => "01101100",5229 => "01011010",5230 => "00101001",5231 => "00010000",5232 => "01110010",5233 => "11101110",5234 => "11001111",5235 => "01001010",5236 => "01010010",5237 => "00001001",5238 => "11001110",5239 => "01001110",5240 => "11111101",5241 => "10111000",5242 => "10000101",5243 => "01110111",5244 => "10000111",5245 => "11000111",5246 => "11001100",5247 => "00100000",5248 => "11001000",5249 => "11100111",5250 => "10000000",5251 => "01000001",5252 => "00101001",5253 => "11111011",5254 => "10001011",5255 => "11010001",5256 => "01111010",5257 => "11100011",5258 => "01101000",5259 => "01000110",5260 => "11101011",5261 => "00011001",5262 => "00001010",5263 => "10101110",5264 => "10001001",5265 => "00001010",5266 => "11011001",5267 => "10011101",5268 => "00101011",5269 => "11111011",5270 => "00101110",5271 => "11100010",5272 => "11101000",5273 => "10101111",5274 => "11110001",5275 => "00000000",5276 => "01110001",5277 => "00000000",5278 => "01111010",5279 => "00001000",5280 => "00000011",5281 => "00111100",5282 => "10110011",5283 => "11100100",5284 => "11110110",5285 => "11101000",5286 => "10001101",5287 => "01000011",5288 => "00100111",5289 => "01000010",5290 => "00011111",5291 => "01110000",5292 => "11000101",5293 => "11011100",5294 => "00111011",5295 => "10011100",5296 => "01010010",5297 => "00111000",5298 => "11000111",5299 => "01000100",5300 => "11111111",5301 => "11101001",5302 => "11110111",5303 => "10100101",5304 => "11101101",5305 => "10011101",5306 => "01101100",5307 => "11110011",5308 => "01000110",5309 => "01111110",5310 => "01000101",5311 => "01110001",5312 => "11100110",5313 => "00111111",5314 => "01011001",5315 => "00011111",5316 => "01010001",5317 => "01010100",5318 => "10101001",5319 => "10001100",5320 => "10110001",5321 => "00100111",5322 => "10001011",5323 => "00000100",5324 => "00001011",5325 => "10010010",5326 => "11100011",5327 => "00010011",5328 => "00010100",5329 => "10111111",5330 => "11000001",5331 => "01010001",5332 => "11101111",5333 => "00011001",5334 => "01010111",5335 => "10011100",5336 => "10101111",5337 => "01100111",5338 => "00011010",5339 => "01111100",5340 => "00101110",5341 => "00101000",5342 => "01110111",5343 => "11111000",5344 => "11111101",5345 => "00001101",5346 => "11001010",5347 => "11111111",5348 => "00110000",5349 => "10010011",5350 => "01101000",5351 => "11001110",5352 => "00100011",5353 => "10101000",5354 => "10111011",5355 => "00000111",5356 => "11010011",5357 => "00000001",5358 => "01010110",5359 => "01111010",5360 => "00110011",5361 => "00011000",5362 => "11011100",5363 => "10001001",5364 => "11001111",5365 => "01011011",5366 => "01101000",5367 => "01110110",5368 => "00001010",5369 => "00010000",5370 => "10101011",5371 => "10110110",5372 => "11110011",5373 => "01100100",5374 => "11001100",5375 => "10001100",5376 => "00001011",5377 => "11111110",5378 => "10010011",5379 => "11100100",5380 => "01011010",5381 => "00011001",5382 => "10010111",5383 => "01101010",5384 => "10110001",5385 => "11000101",5386 => "01010110",5387 => "01000100",5388 => "11000100",5389 => "11110011",5390 => "10010100",5391 => "11010011",5392 => "11111100",5393 => "01111011",5394 => "11010010",5395 => "00000100",5396 => "00100011",5397 => "00010010",5398 => "00101111",5399 => "11100101",5400 => "10100000",5401 => "10111110",5402 => "01110011",5403 => "01111011",5404 => "10001110",5405 => "10101111",5406 => "11000001",5407 => "00100100",5408 => "01101100",5409 => "00010000",5410 => "10000100",5411 => "01001100",5412 => "11010010",5413 => "00010001",5414 => "11100011",5415 => "11010101",5416 => "11001110",5417 => "01111010",5418 => "01001111",5419 => "11011010",5420 => "11100110",5421 => "00111000",5422 => "10001101",5423 => "01110110",5424 => "01000001",5425 => "01000110",5426 => "11000010",5427 => "10011011",5428 => "10001010",5429 => "01110001",5430 => "00011110",5431 => "00000101",5432 => "10001111",5433 => "00100010",5434 => "10101011",5435 => "00100001",5436 => "00000101",5437 => "00000100",5438 => "10101101",5439 => "10000000",5440 => "11101111",5441 => "01000001",5442 => "11101000",5443 => "01000101",5444 => "01001000",5445 => "01100011",5446 => "11101010",5447 => "01111100",5448 => "01101100",5449 => "10000011",5450 => "01100110",5451 => "10001100",5452 => "11101000",5453 => "00000011",5454 => "00000100",5455 => "00010011",5456 => "01101001",5457 => "11101110",5458 => "11000010",5459 => "11111000",5460 => "10010011",5461 => "01101110",5462 => "00111110",5463 => "10000001",5464 => "00111000",5465 => "11100111",5466 => "01011010",5467 => "10011100",5468 => "01010111",5469 => "11100110",5470 => "01011000",5471 => "11011101",5472 => "01000010",5473 => "00101100",5474 => "11001111",5475 => "10101011",5476 => "11000110",5477 => "01100110",5478 => "00011011",5479 => "10011000",5480 => "10111111",5481 => "10000111",5482 => "00001011",5483 => "10000001",5484 => "00111000",5485 => "11011000",5486 => "10011001",5487 => "11001110",5488 => "01100000",5489 => "00000000",5490 => "01011010",5491 => "00010001",5492 => "10100101",5493 => "10000001",5494 => "01110111",5495 => "11011100",5496 => "10011110",5497 => "10001101",5498 => "11101000",5499 => "00100100",5500 => "11010110",5501 => "10010001",5502 => "01111010",5503 => "00011111",5504 => "10101100",5505 => "01000101",5506 => "01001001",5507 => "01110111",5508 => "10010001",5509 => "00110011",5510 => "00101101",5511 => "11111010",5512 => "01111110",5513 => "10110100",5514 => "11000000",5515 => "01011101",5516 => "01111010",others => (others =>'0'));


component project_reti_logiche is 
    port (
            i_clk         : in  std_logic;
            i_start       : in  std_logic;
            i_rst         : in  std_logic;
            i_data       : in  std_logic_vector(7 downto 0); --1 byte
            o_address     : out std_logic_vector(15 downto 0); --16 bit addr: max size is 255*255 + 3 more for max x and y and thresh.
            o_done            : out std_logic;
            o_en         : out std_logic;
            o_we       : out std_logic;
            o_data            : out std_logic_vector (7 downto 0)
          );
end component project_reti_logiche;


begin 
	UUT: project_reti_logiche
	port map (
		  i_clk      	=> tb_clk,	
          i_start       => tb_start,
          i_rst      	=> tb_rst,
          i_data    	=> mem_o_data,
          o_address  	=> mem_address, 
          o_done      	=> tb_done,
          o_en   	=> enable_wire,
		  o_we 	=> mem_we,
          o_data    => mem_i_data
);

p_CLK_GEN : process is
  begin
    wait for c_CLOCK_PERIOD/2;
    tb_clk <= not tb_clk;
  end process p_CLK_GEN; 
  
  
MEM : process(tb_clk)
   begin
    if tb_clk'event and tb_clk = '1' then
     if enable_wire = '1' then
      if mem_we = '1' then
       RAM(conv_integer(mem_address))              <= mem_i_data;
       mem_o_data                      <= mem_i_data;
      else
       mem_o_data <= RAM(conv_integer(mem_address));
      end if;
     end if;
    end if;
   end process;
 
  
  
test : process is
begin 
wait for 100 ns;
wait for c_CLOCK_PERIOD;
tb_rst <= '1';
wait for c_CLOCK_PERIOD;
tb_rst <= '0';
wait for c_CLOCK_PERIOD;
tb_start <= '1';
wait for c_CLOCK_PERIOD; 
tb_start <= '0';
wait until tb_done = '1';
wait until tb_done = '0';
wait until rising_edge(tb_clk); 

assert RAM(1) = "00010101" report "FAIL high bits" severity failure;
assert RAM(0) = "10001100" report "FAIL low bits" severity failure;


assert false report "Simulation Ended!, test passed" severity failure;
end process test;

end projecttb; 
